# ________________________________________________________________________________________________
# 
# 
#             Synchronous One-Port Register File Compiler
# 
#                 UMC 0.11um LL AE Logic Process
# 
# ________________________________________________________________________________________________
# 
#               
#         Copyright (C) 2024 Faraday Technology Corporation. All Rights Reserved.       
#                
#         This source code is an unpublished work belongs to Faraday Technology Corporation       
#         It is considered a trade secret and is not to be divulged or       
#         used by parties who have not received written authorization from       
#         Faraday Technology Corporation       
#                
#         Faraday's home page can be found at: http://www.faraday-tech.com/       
#                
# ________________________________________________________________________________________________
# 
#        IP Name            :  FSR0K_B_SY                
#        IP Version         :  1.4.0                     
#        IP Release Status  :  Active                    
#        Word               :  32                        
#        Bit                :  8                         
#        Byte               :  16                        
#        Mux                :  2                         
#        Output Loading     :  0.01                      
#        Clock Input Slew   :  0.016                     
#        Data Input Slew    :  0.016                     
#        Ring Type          :  Ringless Model            
#        Ring Width         :  0                         
#        Bus Format         :  0                         
#        Memaker Path       :  /home/mem/Desktop/memlib  
#        GUI Version        :  m20230904                 
#        Date               :  2024/11/05 22:37:10       
# ________________________________________________________________________________________________
# 

VERSION 5.5 ;
NAMESCASESENSITIVE ON ;
MACRO SYKB110_32X8X16CM2
CLASS BLOCK ;
FOREIGN SYKB110_32X8X16CM2 0.000 0.000 ;
ORIGIN 0.000 0.000 ;
SIZE 554.411 BY 66.831 ;
SYMMETRY x y r90 ;
SITE core ;
PIN GND
  DIRECTION INOUT ;
  USE GROUND ;
 PORT
  LAYER ME4 ;
  RECT 299.078 1.781 299.418 66.831 ;
 END
 PORT
  LAYER ME4 ;
  RECT 295.074 1.781 295.414 66.831 ;
 END
 PORT
  LAYER ME4 ;
  RECT 297.076 1.781 297.416 66.831 ;
 END
 PORT
  LAYER ME4 ;
  RECT 297.887 0.000 298.607 44.094 ;
 END
 PORT
  LAYER ME4 ;
  RECT 303.082 1.781 303.422 66.831 ;
 END
 PORT
  LAYER ME4 ;
  RECT 301.080 1.781 301.420 66.831 ;
 END
 PORT
  LAYER ME4 ;
  RECT 301.891 0.000 302.611 44.094 ;
 END
 PORT
  LAYER ME4 ;
  RECT 307.086 1.781 307.426 66.831 ;
 END
 PORT
  LAYER ME4 ;
  RECT 305.084 1.781 305.424 66.831 ;
 END
 PORT
  LAYER ME4 ;
  RECT 305.895 0.000 306.615 44.094 ;
 END
 PORT
  LAYER ME4 ;
  RECT 311.090 1.781 311.430 66.831 ;
 END
 PORT
  LAYER ME4 ;
  RECT 309.088 1.781 309.428 66.831 ;
 END
 PORT
  LAYER ME4 ;
  RECT 309.899 0.000 310.619 44.094 ;
 END
 PORT
  LAYER ME4 ;
  RECT 315.094 1.781 315.434 66.831 ;
 END
 PORT
  LAYER ME4 ;
  RECT 313.092 1.781 313.432 66.831 ;
 END
 PORT
  LAYER ME4 ;
  RECT 313.903 0.000 314.623 44.094 ;
 END
 PORT
  LAYER ME4 ;
  RECT 319.098 1.781 319.438 66.831 ;
 END
 PORT
  LAYER ME4 ;
  RECT 317.096 1.781 317.436 66.831 ;
 END
 PORT
  LAYER ME4 ;
  RECT 317.907 0.000 318.627 44.094 ;
 END
 PORT
  LAYER ME4 ;
  RECT 323.102 1.781 323.442 66.831 ;
 END
 PORT
  LAYER ME4 ;
  RECT 321.100 1.781 321.440 66.831 ;
 END
 PORT
  LAYER ME4 ;
  RECT 321.911 0.000 322.631 44.094 ;
 END
 PORT
  LAYER ME4 ;
  RECT 327.106 1.781 327.446 66.831 ;
 END
 PORT
  LAYER ME4 ;
  RECT 325.104 1.781 325.444 66.831 ;
 END
 PORT
  LAYER ME4 ;
  RECT 325.915 0.000 326.635 44.094 ;
 END
 PORT
  LAYER ME4 ;
  RECT 331.110 1.781 331.450 66.831 ;
 END
 PORT
  LAYER ME4 ;
  RECT 329.108 1.781 329.448 66.831 ;
 END
 PORT
  LAYER ME4 ;
  RECT 329.919 0.000 330.639 44.094 ;
 END
 PORT
  LAYER ME4 ;
  RECT 335.114 1.781 335.454 66.831 ;
 END
 PORT
  LAYER ME4 ;
  RECT 333.112 1.781 333.452 66.831 ;
 END
 PORT
  LAYER ME4 ;
  RECT 333.923 0.000 334.643 44.094 ;
 END
 PORT
  LAYER ME4 ;
  RECT 339.118 1.781 339.458 66.831 ;
 END
 PORT
  LAYER ME4 ;
  RECT 337.116 1.781 337.456 66.831 ;
 END
 PORT
  LAYER ME4 ;
  RECT 337.927 0.000 338.647 44.094 ;
 END
 PORT
  LAYER ME4 ;
  RECT 343.122 1.781 343.462 66.831 ;
 END
 PORT
  LAYER ME4 ;
  RECT 341.120 1.781 341.460 66.831 ;
 END
 PORT
  LAYER ME4 ;
  RECT 341.931 0.000 342.651 44.094 ;
 END
 PORT
  LAYER ME4 ;
  RECT 347.126 1.781 347.466 66.831 ;
 END
 PORT
  LAYER ME4 ;
  RECT 345.124 1.781 345.464 66.831 ;
 END
 PORT
  LAYER ME4 ;
  RECT 345.935 0.000 346.655 44.094 ;
 END
 PORT
  LAYER ME4 ;
  RECT 351.130 1.781 351.470 66.831 ;
 END
 PORT
  LAYER ME4 ;
  RECT 349.128 1.781 349.468 66.831 ;
 END
 PORT
  LAYER ME4 ;
  RECT 349.939 0.000 350.659 44.094 ;
 END
 PORT
  LAYER ME4 ;
  RECT 355.134 1.781 355.474 66.831 ;
 END
 PORT
  LAYER ME4 ;
  RECT 353.132 1.781 353.472 66.831 ;
 END
 PORT
  LAYER ME4 ;
  RECT 353.943 0.000 354.663 44.094 ;
 END
 PORT
  LAYER ME4 ;
  RECT 359.138 1.781 359.478 66.831 ;
 END
 PORT
  LAYER ME4 ;
  RECT 357.136 1.781 357.476 66.831 ;
 END
 PORT
  LAYER ME4 ;
  RECT 357.947 0.000 358.667 44.094 ;
 END
 PORT
  LAYER ME4 ;
  RECT 363.142 1.781 363.482 66.831 ;
 END
 PORT
  LAYER ME4 ;
  RECT 361.140 1.781 361.480 66.831 ;
 END
 PORT
  LAYER ME4 ;
  RECT 361.951 0.000 362.671 44.094 ;
 END
 PORT
  LAYER ME4 ;
  RECT 367.146 1.781 367.486 66.831 ;
 END
 PORT
  LAYER ME4 ;
  RECT 365.144 1.781 365.484 66.831 ;
 END
 PORT
  LAYER ME4 ;
  RECT 365.955 0.000 366.675 44.094 ;
 END
 PORT
  LAYER ME4 ;
  RECT 371.150 1.781 371.490 66.831 ;
 END
 PORT
  LAYER ME4 ;
  RECT 369.148 1.781 369.488 66.831 ;
 END
 PORT
  LAYER ME4 ;
  RECT 369.959 0.000 370.679 44.094 ;
 END
 PORT
  LAYER ME4 ;
  RECT 375.154 1.781 375.494 66.831 ;
 END
 PORT
  LAYER ME4 ;
  RECT 373.152 1.781 373.492 66.831 ;
 END
 PORT
  LAYER ME4 ;
  RECT 373.963 0.000 374.683 44.094 ;
 END
 PORT
  LAYER ME4 ;
  RECT 379.158 1.781 379.498 66.831 ;
 END
 PORT
  LAYER ME4 ;
  RECT 377.156 1.781 377.496 66.831 ;
 END
 PORT
  LAYER ME4 ;
  RECT 377.967 0.000 378.687 44.094 ;
 END
 PORT
  LAYER ME4 ;
  RECT 383.162 1.781 383.502 66.831 ;
 END
 PORT
  LAYER ME4 ;
  RECT 381.160 1.781 381.500 66.831 ;
 END
 PORT
  LAYER ME4 ;
  RECT 381.971 0.000 382.691 44.094 ;
 END
 PORT
  LAYER ME4 ;
  RECT 387.166 1.781 387.506 66.831 ;
 END
 PORT
  LAYER ME4 ;
  RECT 385.164 1.781 385.504 66.831 ;
 END
 PORT
  LAYER ME4 ;
  RECT 385.975 0.000 386.695 44.094 ;
 END
 PORT
  LAYER ME4 ;
  RECT 391.170 1.781 391.510 66.831 ;
 END
 PORT
  LAYER ME4 ;
  RECT 389.168 1.781 389.508 66.831 ;
 END
 PORT
  LAYER ME4 ;
  RECT 389.979 0.000 390.699 44.094 ;
 END
 PORT
  LAYER ME4 ;
  RECT 395.174 1.781 395.514 66.831 ;
 END
 PORT
  LAYER ME4 ;
  RECT 393.172 1.781 393.512 66.831 ;
 END
 PORT
  LAYER ME4 ;
  RECT 393.983 0.000 394.703 44.094 ;
 END
 PORT
  LAYER ME4 ;
  RECT 399.178 1.781 399.518 66.831 ;
 END
 PORT
  LAYER ME4 ;
  RECT 397.176 1.781 397.516 66.831 ;
 END
 PORT
  LAYER ME4 ;
  RECT 397.987 0.000 398.707 44.094 ;
 END
 PORT
  LAYER ME4 ;
  RECT 403.182 1.781 403.522 66.831 ;
 END
 PORT
  LAYER ME4 ;
  RECT 401.180 1.781 401.520 66.831 ;
 END
 PORT
  LAYER ME4 ;
  RECT 401.991 0.000 402.711 44.094 ;
 END
 PORT
  LAYER ME4 ;
  RECT 407.186 1.781 407.526 66.831 ;
 END
 PORT
  LAYER ME4 ;
  RECT 405.184 1.781 405.524 66.831 ;
 END
 PORT
  LAYER ME4 ;
  RECT 405.995 0.000 406.715 44.094 ;
 END
 PORT
  LAYER ME4 ;
  RECT 411.190 1.781 411.530 66.831 ;
 END
 PORT
  LAYER ME4 ;
  RECT 409.188 1.781 409.528 66.831 ;
 END
 PORT
  LAYER ME4 ;
  RECT 409.999 0.000 410.719 44.094 ;
 END
 PORT
  LAYER ME4 ;
  RECT 415.194 1.781 415.534 66.831 ;
 END
 PORT
  LAYER ME4 ;
  RECT 413.192 1.781 413.532 66.831 ;
 END
 PORT
  LAYER ME4 ;
  RECT 414.003 0.000 414.723 44.094 ;
 END
 PORT
  LAYER ME4 ;
  RECT 419.198 1.781 419.538 66.831 ;
 END
 PORT
  LAYER ME4 ;
  RECT 417.196 1.781 417.536 66.831 ;
 END
 PORT
  LAYER ME4 ;
  RECT 418.007 0.000 418.727 44.094 ;
 END
 PORT
  LAYER ME4 ;
  RECT 423.202 1.781 423.542 66.831 ;
 END
 PORT
  LAYER ME4 ;
  RECT 421.200 1.781 421.540 66.831 ;
 END
 PORT
  LAYER ME4 ;
  RECT 422.011 0.000 422.731 44.094 ;
 END
 PORT
  LAYER ME4 ;
  RECT 427.206 1.781 427.546 66.831 ;
 END
 PORT
  LAYER ME4 ;
  RECT 425.204 1.781 425.544 66.831 ;
 END
 PORT
  LAYER ME4 ;
  RECT 426.015 0.000 426.735 44.094 ;
 END
 PORT
  LAYER ME4 ;
  RECT 431.210 1.781 431.550 66.831 ;
 END
 PORT
  LAYER ME4 ;
  RECT 429.208 1.781 429.548 66.831 ;
 END
 PORT
  LAYER ME4 ;
  RECT 430.019 0.000 430.739 44.094 ;
 END
 PORT
  LAYER ME4 ;
  RECT 435.214 1.781 435.554 66.831 ;
 END
 PORT
  LAYER ME4 ;
  RECT 433.212 1.781 433.552 66.831 ;
 END
 PORT
  LAYER ME4 ;
  RECT 434.023 0.000 434.743 44.094 ;
 END
 PORT
  LAYER ME4 ;
  RECT 439.218 1.781 439.558 66.831 ;
 END
 PORT
  LAYER ME4 ;
  RECT 437.216 1.781 437.556 66.831 ;
 END
 PORT
  LAYER ME4 ;
  RECT 438.027 0.000 438.747 44.094 ;
 END
 PORT
  LAYER ME4 ;
  RECT 443.222 1.781 443.562 66.831 ;
 END
 PORT
  LAYER ME4 ;
  RECT 441.220 1.781 441.560 66.831 ;
 END
 PORT
  LAYER ME4 ;
  RECT 442.031 0.000 442.751 44.094 ;
 END
 PORT
  LAYER ME4 ;
  RECT 447.226 1.781 447.566 66.831 ;
 END
 PORT
  LAYER ME4 ;
  RECT 445.224 1.781 445.564 66.831 ;
 END
 PORT
  LAYER ME4 ;
  RECT 446.035 0.000 446.755 44.094 ;
 END
 PORT
  LAYER ME4 ;
  RECT 451.230 1.781 451.570 66.831 ;
 END
 PORT
  LAYER ME4 ;
  RECT 449.228 1.781 449.568 66.831 ;
 END
 PORT
  LAYER ME4 ;
  RECT 450.039 0.000 450.759 44.094 ;
 END
 PORT
  LAYER ME4 ;
  RECT 455.234 1.781 455.574 66.831 ;
 END
 PORT
  LAYER ME4 ;
  RECT 453.232 1.781 453.572 66.831 ;
 END
 PORT
  LAYER ME4 ;
  RECT 454.043 0.000 454.763 44.094 ;
 END
 PORT
  LAYER ME4 ;
  RECT 459.238 1.781 459.578 66.831 ;
 END
 PORT
  LAYER ME4 ;
  RECT 457.236 1.781 457.576 66.831 ;
 END
 PORT
  LAYER ME4 ;
  RECT 458.047 0.000 458.767 44.094 ;
 END
 PORT
  LAYER ME4 ;
  RECT 463.242 1.781 463.582 66.831 ;
 END
 PORT
  LAYER ME4 ;
  RECT 461.240 1.781 461.580 66.831 ;
 END
 PORT
  LAYER ME4 ;
  RECT 462.051 0.000 462.771 44.094 ;
 END
 PORT
  LAYER ME4 ;
  RECT 467.246 1.781 467.586 66.831 ;
 END
 PORT
  LAYER ME4 ;
  RECT 465.244 1.781 465.584 66.831 ;
 END
 PORT
  LAYER ME4 ;
  RECT 466.055 0.000 466.775 44.094 ;
 END
 PORT
  LAYER ME4 ;
  RECT 471.250 1.781 471.590 66.831 ;
 END
 PORT
  LAYER ME4 ;
  RECT 469.248 1.781 469.588 66.831 ;
 END
 PORT
  LAYER ME4 ;
  RECT 470.059 0.000 470.779 44.094 ;
 END
 PORT
  LAYER ME4 ;
  RECT 475.254 1.781 475.594 66.831 ;
 END
 PORT
  LAYER ME4 ;
  RECT 473.252 1.781 473.592 66.831 ;
 END
 PORT
  LAYER ME4 ;
  RECT 474.063 0.000 474.783 44.094 ;
 END
 PORT
  LAYER ME4 ;
  RECT 479.258 1.781 479.598 66.831 ;
 END
 PORT
  LAYER ME4 ;
  RECT 477.256 1.781 477.596 66.831 ;
 END
 PORT
  LAYER ME4 ;
  RECT 478.067 0.000 478.787 44.094 ;
 END
 PORT
  LAYER ME4 ;
  RECT 483.262 1.781 483.602 66.831 ;
 END
 PORT
  LAYER ME4 ;
  RECT 481.260 1.781 481.600 66.831 ;
 END
 PORT
  LAYER ME4 ;
  RECT 482.071 0.000 482.791 44.094 ;
 END
 PORT
  LAYER ME4 ;
  RECT 487.266 1.781 487.606 66.831 ;
 END
 PORT
  LAYER ME4 ;
  RECT 485.264 1.781 485.604 66.831 ;
 END
 PORT
  LAYER ME4 ;
  RECT 486.075 0.000 486.795 44.094 ;
 END
 PORT
  LAYER ME4 ;
  RECT 491.270 1.781 491.610 66.831 ;
 END
 PORT
  LAYER ME4 ;
  RECT 489.268 1.781 489.608 66.831 ;
 END
 PORT
  LAYER ME4 ;
  RECT 490.079 0.000 490.799 44.094 ;
 END
 PORT
  LAYER ME4 ;
  RECT 495.274 1.781 495.614 66.831 ;
 END
 PORT
  LAYER ME4 ;
  RECT 493.272 1.781 493.612 66.831 ;
 END
 PORT
  LAYER ME4 ;
  RECT 494.083 0.000 494.803 44.094 ;
 END
 PORT
  LAYER ME4 ;
  RECT 499.278 1.781 499.618 66.831 ;
 END
 PORT
  LAYER ME4 ;
  RECT 497.276 1.781 497.616 66.831 ;
 END
 PORT
  LAYER ME4 ;
  RECT 498.087 0.000 498.807 44.094 ;
 END
 PORT
  LAYER ME4 ;
  RECT 503.282 1.781 503.622 66.831 ;
 END
 PORT
  LAYER ME4 ;
  RECT 501.280 1.781 501.620 66.831 ;
 END
 PORT
  LAYER ME4 ;
  RECT 502.091 0.000 502.811 44.094 ;
 END
 PORT
  LAYER ME4 ;
  RECT 507.286 1.781 507.626 66.831 ;
 END
 PORT
  LAYER ME4 ;
  RECT 505.284 1.781 505.624 66.831 ;
 END
 PORT
  LAYER ME4 ;
  RECT 506.095 0.000 506.815 44.094 ;
 END
 PORT
  LAYER ME4 ;
  RECT 511.290 1.781 511.630 66.831 ;
 END
 PORT
  LAYER ME4 ;
  RECT 509.288 1.781 509.628 66.831 ;
 END
 PORT
  LAYER ME4 ;
  RECT 510.099 0.000 510.819 44.094 ;
 END
 PORT
  LAYER ME4 ;
  RECT 515.294 1.781 515.634 66.831 ;
 END
 PORT
  LAYER ME4 ;
  RECT 513.292 1.781 513.632 66.831 ;
 END
 PORT
  LAYER ME4 ;
  RECT 514.103 0.000 514.823 44.094 ;
 END
 PORT
  LAYER ME4 ;
  RECT 519.298 1.781 519.638 66.831 ;
 END
 PORT
  LAYER ME4 ;
  RECT 517.296 1.781 517.636 66.831 ;
 END
 PORT
  LAYER ME4 ;
  RECT 518.107 0.000 518.827 44.094 ;
 END
 PORT
  LAYER ME4 ;
  RECT 523.302 1.781 523.642 66.831 ;
 END
 PORT
  LAYER ME4 ;
  RECT 521.300 1.781 521.640 66.831 ;
 END
 PORT
  LAYER ME4 ;
  RECT 522.111 0.000 522.831 44.094 ;
 END
 PORT
  LAYER ME4 ;
  RECT 527.306 1.781 527.646 66.831 ;
 END
 PORT
  LAYER ME4 ;
  RECT 525.304 1.781 525.644 66.831 ;
 END
 PORT
  LAYER ME4 ;
  RECT 526.115 0.000 526.835 44.094 ;
 END
 PORT
  LAYER ME4 ;
  RECT 531.310 1.781 531.650 66.831 ;
 END
 PORT
  LAYER ME4 ;
  RECT 529.308 1.781 529.648 66.831 ;
 END
 PORT
  LAYER ME4 ;
  RECT 530.119 0.000 530.839 44.094 ;
 END
 PORT
  LAYER ME4 ;
  RECT 535.314 1.781 535.654 66.831 ;
 END
 PORT
  LAYER ME4 ;
  RECT 533.312 1.781 533.652 66.831 ;
 END
 PORT
  LAYER ME4 ;
  RECT 534.123 0.000 534.843 44.094 ;
 END
 PORT
  LAYER ME4 ;
  RECT 539.318 1.781 539.658 66.831 ;
 END
 PORT
  LAYER ME4 ;
  RECT 537.316 1.781 537.656 66.831 ;
 END
 PORT
  LAYER ME4 ;
  RECT 538.127 0.000 538.847 44.094 ;
 END
 PORT
  LAYER ME4 ;
  RECT 543.322 1.781 543.662 66.831 ;
 END
 PORT
  LAYER ME4 ;
  RECT 541.320 1.781 541.660 66.831 ;
 END
 PORT
  LAYER ME4 ;
  RECT 542.131 0.000 542.851 44.094 ;
 END
 PORT
  LAYER ME4 ;
  RECT 547.326 1.781 547.666 66.831 ;
 END
 PORT
  LAYER ME4 ;
  RECT 545.324 1.781 545.664 66.831 ;
 END
 PORT
  LAYER ME4 ;
  RECT 546.135 0.000 546.855 44.094 ;
 END
 PORT
  LAYER ME4 ;
  RECT 551.330 1.781 551.670 66.831 ;
 END
 PORT
  LAYER ME4 ;
  RECT 549.328 1.781 549.668 66.831 ;
 END
 PORT
  LAYER ME4 ;
  RECT 550.139 0.000 550.859 44.094 ;
 END
 PORT
  LAYER ME4 ;
  RECT 552.331 0.000 552.671 66.831 ;
 END
 PORT
  LAYER ME4 ;
  RECT 276.217 0.000 276.937 66.831 ;
 END
 PORT
  LAYER ME4 ;
  RECT 282.211 0.000 282.931 66.831 ;
 END
 PORT
  LAYER ME4 ;
  RECT 287.682 0.000 288.402 66.831 ;
 END
 PORT
  LAYER ME4 ;
  RECT 289.397 0.000 290.117 66.831 ;
 END
 PORT
  LAYER ME4 ;
  RECT 292.393 0.000 292.993 66.831 ;
 END
 PORT
  LAYER ME4 ;
  RECT 294.073 1.781 294.413 66.831 ;
 END
 PORT
  LAYER ME4 ;
  RECT 268.658 0.000 269.378 66.831 ;
 END
 PORT
  LAYER ME4 ;
  RECT 266.618 1.781 267.338 66.072 ;
 END
 PORT
  LAYER ME4 ;
  RECT 1.740 0.000 2.080 66.831 ;
 END
 PORT
  LAYER ME4 ;
  RECT 6.745 1.781 7.085 66.831 ;
 END
 PORT
  LAYER ME4 ;
  RECT 2.741 1.781 3.081 66.831 ;
 END
 PORT
  LAYER ME4 ;
  RECT 4.743 1.781 5.083 66.831 ;
 END
 PORT
  LAYER ME4 ;
  RECT 5.554 0.000 6.274 44.094 ;
 END
 PORT
  LAYER ME4 ;
  RECT 10.749 1.781 11.089 66.831 ;
 END
 PORT
  LAYER ME4 ;
  RECT 8.747 1.781 9.087 66.831 ;
 END
 PORT
  LAYER ME4 ;
  RECT 9.558 0.000 10.278 44.094 ;
 END
 PORT
  LAYER ME4 ;
  RECT 14.753 1.781 15.093 66.831 ;
 END
 PORT
  LAYER ME4 ;
  RECT 12.751 1.781 13.091 66.831 ;
 END
 PORT
  LAYER ME4 ;
  RECT 13.562 0.000 14.282 44.094 ;
 END
 PORT
  LAYER ME4 ;
  RECT 18.757 1.781 19.097 66.831 ;
 END
 PORT
  LAYER ME4 ;
  RECT 16.755 1.781 17.095 66.831 ;
 END
 PORT
  LAYER ME4 ;
  RECT 17.566 0.000 18.286 44.094 ;
 END
 PORT
  LAYER ME4 ;
  RECT 22.761 1.781 23.101 66.831 ;
 END
 PORT
  LAYER ME4 ;
  RECT 20.759 1.781 21.099 66.831 ;
 END
 PORT
  LAYER ME4 ;
  RECT 21.570 0.000 22.290 44.094 ;
 END
 PORT
  LAYER ME4 ;
  RECT 26.765 1.781 27.105 66.831 ;
 END
 PORT
  LAYER ME4 ;
  RECT 24.763 1.781 25.103 66.831 ;
 END
 PORT
  LAYER ME4 ;
  RECT 25.574 0.000 26.294 44.094 ;
 END
 PORT
  LAYER ME4 ;
  RECT 30.769 1.781 31.109 66.831 ;
 END
 PORT
  LAYER ME4 ;
  RECT 28.767 1.781 29.107 66.831 ;
 END
 PORT
  LAYER ME4 ;
  RECT 29.578 0.000 30.298 44.094 ;
 END
 PORT
  LAYER ME4 ;
  RECT 34.773 1.781 35.113 66.831 ;
 END
 PORT
  LAYER ME4 ;
  RECT 32.771 1.781 33.111 66.831 ;
 END
 PORT
  LAYER ME4 ;
  RECT 33.582 0.000 34.302 44.094 ;
 END
 PORT
  LAYER ME4 ;
  RECT 38.777 1.781 39.117 66.831 ;
 END
 PORT
  LAYER ME4 ;
  RECT 36.775 1.781 37.115 66.831 ;
 END
 PORT
  LAYER ME4 ;
  RECT 37.586 0.000 38.306 44.094 ;
 END
 PORT
  LAYER ME4 ;
  RECT 42.781 1.781 43.121 66.831 ;
 END
 PORT
  LAYER ME4 ;
  RECT 40.779 1.781 41.119 66.831 ;
 END
 PORT
  LAYER ME4 ;
  RECT 41.590 0.000 42.310 44.094 ;
 END
 PORT
  LAYER ME4 ;
  RECT 46.785 1.781 47.125 66.831 ;
 END
 PORT
  LAYER ME4 ;
  RECT 44.783 1.781 45.123 66.831 ;
 END
 PORT
  LAYER ME4 ;
  RECT 45.594 0.000 46.314 44.094 ;
 END
 PORT
  LAYER ME4 ;
  RECT 50.789 1.781 51.129 66.831 ;
 END
 PORT
  LAYER ME4 ;
  RECT 48.787 1.781 49.127 66.831 ;
 END
 PORT
  LAYER ME4 ;
  RECT 49.598 0.000 50.318 44.094 ;
 END
 PORT
  LAYER ME4 ;
  RECT 54.793 1.781 55.133 66.831 ;
 END
 PORT
  LAYER ME4 ;
  RECT 52.791 1.781 53.131 66.831 ;
 END
 PORT
  LAYER ME4 ;
  RECT 53.602 0.000 54.322 44.094 ;
 END
 PORT
  LAYER ME4 ;
  RECT 58.797 1.781 59.137 66.831 ;
 END
 PORT
  LAYER ME4 ;
  RECT 56.795 1.781 57.135 66.831 ;
 END
 PORT
  LAYER ME4 ;
  RECT 57.606 0.000 58.326 44.094 ;
 END
 PORT
  LAYER ME4 ;
  RECT 62.801 1.781 63.141 66.831 ;
 END
 PORT
  LAYER ME4 ;
  RECT 60.799 1.781 61.139 66.831 ;
 END
 PORT
  LAYER ME4 ;
  RECT 61.610 0.000 62.330 44.094 ;
 END
 PORT
  LAYER ME4 ;
  RECT 66.805 1.781 67.145 66.831 ;
 END
 PORT
  LAYER ME4 ;
  RECT 64.803 1.781 65.143 66.831 ;
 END
 PORT
  LAYER ME4 ;
  RECT 65.614 0.000 66.334 44.094 ;
 END
 PORT
  LAYER ME4 ;
  RECT 70.809 1.781 71.149 66.831 ;
 END
 PORT
  LAYER ME4 ;
  RECT 68.807 1.781 69.147 66.831 ;
 END
 PORT
  LAYER ME4 ;
  RECT 69.618 0.000 70.338 44.094 ;
 END
 PORT
  LAYER ME4 ;
  RECT 74.813 1.781 75.153 66.831 ;
 END
 PORT
  LAYER ME4 ;
  RECT 72.811 1.781 73.151 66.831 ;
 END
 PORT
  LAYER ME4 ;
  RECT 73.622 0.000 74.342 44.094 ;
 END
 PORT
  LAYER ME4 ;
  RECT 78.817 1.781 79.157 66.831 ;
 END
 PORT
  LAYER ME4 ;
  RECT 76.815 1.781 77.155 66.831 ;
 END
 PORT
  LAYER ME4 ;
  RECT 77.626 0.000 78.346 44.094 ;
 END
 PORT
  LAYER ME4 ;
  RECT 82.821 1.781 83.161 66.831 ;
 END
 PORT
  LAYER ME4 ;
  RECT 80.819 1.781 81.159 66.831 ;
 END
 PORT
  LAYER ME4 ;
  RECT 81.630 0.000 82.350 44.094 ;
 END
 PORT
  LAYER ME4 ;
  RECT 86.825 1.781 87.165 66.831 ;
 END
 PORT
  LAYER ME4 ;
  RECT 84.823 1.781 85.163 66.831 ;
 END
 PORT
  LAYER ME4 ;
  RECT 85.634 0.000 86.354 44.094 ;
 END
 PORT
  LAYER ME4 ;
  RECT 90.829 1.781 91.169 66.831 ;
 END
 PORT
  LAYER ME4 ;
  RECT 88.827 1.781 89.167 66.831 ;
 END
 PORT
  LAYER ME4 ;
  RECT 89.638 0.000 90.358 44.094 ;
 END
 PORT
  LAYER ME4 ;
  RECT 94.833 1.781 95.173 66.831 ;
 END
 PORT
  LAYER ME4 ;
  RECT 92.831 1.781 93.171 66.831 ;
 END
 PORT
  LAYER ME4 ;
  RECT 93.642 0.000 94.362 44.094 ;
 END
 PORT
  LAYER ME4 ;
  RECT 98.837 1.781 99.177 66.831 ;
 END
 PORT
  LAYER ME4 ;
  RECT 96.835 1.781 97.175 66.831 ;
 END
 PORT
  LAYER ME4 ;
  RECT 97.646 0.000 98.366 44.094 ;
 END
 PORT
  LAYER ME4 ;
  RECT 102.841 1.781 103.181 66.831 ;
 END
 PORT
  LAYER ME4 ;
  RECT 100.839 1.781 101.179 66.831 ;
 END
 PORT
  LAYER ME4 ;
  RECT 101.650 0.000 102.370 44.094 ;
 END
 PORT
  LAYER ME4 ;
  RECT 106.845 1.781 107.185 66.831 ;
 END
 PORT
  LAYER ME4 ;
  RECT 104.843 1.781 105.183 66.831 ;
 END
 PORT
  LAYER ME4 ;
  RECT 105.654 0.000 106.374 44.094 ;
 END
 PORT
  LAYER ME4 ;
  RECT 110.849 1.781 111.189 66.831 ;
 END
 PORT
  LAYER ME4 ;
  RECT 108.847 1.781 109.187 66.831 ;
 END
 PORT
  LAYER ME4 ;
  RECT 109.658 0.000 110.378 44.094 ;
 END
 PORT
  LAYER ME4 ;
  RECT 114.853 1.781 115.193 66.831 ;
 END
 PORT
  LAYER ME4 ;
  RECT 112.851 1.781 113.191 66.831 ;
 END
 PORT
  LAYER ME4 ;
  RECT 113.662 0.000 114.382 44.094 ;
 END
 PORT
  LAYER ME4 ;
  RECT 118.857 1.781 119.197 66.831 ;
 END
 PORT
  LAYER ME4 ;
  RECT 116.855 1.781 117.195 66.831 ;
 END
 PORT
  LAYER ME4 ;
  RECT 117.666 0.000 118.386 44.094 ;
 END
 PORT
  LAYER ME4 ;
  RECT 122.861 1.781 123.201 66.831 ;
 END
 PORT
  LAYER ME4 ;
  RECT 120.859 1.781 121.199 66.831 ;
 END
 PORT
  LAYER ME4 ;
  RECT 121.670 0.000 122.390 44.094 ;
 END
 PORT
  LAYER ME4 ;
  RECT 126.865 1.781 127.205 66.831 ;
 END
 PORT
  LAYER ME4 ;
  RECT 124.863 1.781 125.203 66.831 ;
 END
 PORT
  LAYER ME4 ;
  RECT 125.674 0.000 126.394 44.094 ;
 END
 PORT
  LAYER ME4 ;
  RECT 130.869 1.781 131.209 66.831 ;
 END
 PORT
  LAYER ME4 ;
  RECT 128.867 1.781 129.207 66.831 ;
 END
 PORT
  LAYER ME4 ;
  RECT 129.678 0.000 130.398 44.094 ;
 END
 PORT
  LAYER ME4 ;
  RECT 134.873 1.781 135.213 66.831 ;
 END
 PORT
  LAYER ME4 ;
  RECT 132.871 1.781 133.211 66.831 ;
 END
 PORT
  LAYER ME4 ;
  RECT 133.682 0.000 134.402 44.094 ;
 END
 PORT
  LAYER ME4 ;
  RECT 138.877 1.781 139.217 66.831 ;
 END
 PORT
  LAYER ME4 ;
  RECT 136.875 1.781 137.215 66.831 ;
 END
 PORT
  LAYER ME4 ;
  RECT 137.686 0.000 138.406 44.094 ;
 END
 PORT
  LAYER ME4 ;
  RECT 142.881 1.781 143.221 66.831 ;
 END
 PORT
  LAYER ME4 ;
  RECT 140.879 1.781 141.219 66.831 ;
 END
 PORT
  LAYER ME4 ;
  RECT 141.690 0.000 142.410 44.094 ;
 END
 PORT
  LAYER ME4 ;
  RECT 146.885 1.781 147.225 66.831 ;
 END
 PORT
  LAYER ME4 ;
  RECT 144.883 1.781 145.223 66.831 ;
 END
 PORT
  LAYER ME4 ;
  RECT 145.694 0.000 146.414 44.094 ;
 END
 PORT
  LAYER ME4 ;
  RECT 150.889 1.781 151.229 66.831 ;
 END
 PORT
  LAYER ME4 ;
  RECT 148.887 1.781 149.227 66.831 ;
 END
 PORT
  LAYER ME4 ;
  RECT 149.698 0.000 150.418 44.094 ;
 END
 PORT
  LAYER ME4 ;
  RECT 154.893 1.781 155.233 66.831 ;
 END
 PORT
  LAYER ME4 ;
  RECT 152.891 1.781 153.231 66.831 ;
 END
 PORT
  LAYER ME4 ;
  RECT 153.702 0.000 154.422 44.094 ;
 END
 PORT
  LAYER ME4 ;
  RECT 158.897 1.781 159.237 66.831 ;
 END
 PORT
  LAYER ME4 ;
  RECT 156.895 1.781 157.235 66.831 ;
 END
 PORT
  LAYER ME4 ;
  RECT 157.706 0.000 158.426 44.094 ;
 END
 PORT
  LAYER ME4 ;
  RECT 162.901 1.781 163.241 66.831 ;
 END
 PORT
  LAYER ME4 ;
  RECT 160.899 1.781 161.239 66.831 ;
 END
 PORT
  LAYER ME4 ;
  RECT 161.710 0.000 162.430 44.094 ;
 END
 PORT
  LAYER ME4 ;
  RECT 166.905 1.781 167.245 66.831 ;
 END
 PORT
  LAYER ME4 ;
  RECT 164.903 1.781 165.243 66.831 ;
 END
 PORT
  LAYER ME4 ;
  RECT 165.714 0.000 166.434 44.094 ;
 END
 PORT
  LAYER ME4 ;
  RECT 170.909 1.781 171.249 66.831 ;
 END
 PORT
  LAYER ME4 ;
  RECT 168.907 1.781 169.247 66.831 ;
 END
 PORT
  LAYER ME4 ;
  RECT 169.718 0.000 170.438 44.094 ;
 END
 PORT
  LAYER ME4 ;
  RECT 174.913 1.781 175.253 66.831 ;
 END
 PORT
  LAYER ME4 ;
  RECT 172.911 1.781 173.251 66.831 ;
 END
 PORT
  LAYER ME4 ;
  RECT 173.722 0.000 174.442 44.094 ;
 END
 PORT
  LAYER ME4 ;
  RECT 178.917 1.781 179.257 66.831 ;
 END
 PORT
  LAYER ME4 ;
  RECT 176.915 1.781 177.255 66.831 ;
 END
 PORT
  LAYER ME4 ;
  RECT 177.726 0.000 178.446 44.094 ;
 END
 PORT
  LAYER ME4 ;
  RECT 182.921 1.781 183.261 66.831 ;
 END
 PORT
  LAYER ME4 ;
  RECT 180.919 1.781 181.259 66.831 ;
 END
 PORT
  LAYER ME4 ;
  RECT 181.730 0.000 182.450 44.094 ;
 END
 PORT
  LAYER ME4 ;
  RECT 186.925 1.781 187.265 66.831 ;
 END
 PORT
  LAYER ME4 ;
  RECT 184.923 1.781 185.263 66.831 ;
 END
 PORT
  LAYER ME4 ;
  RECT 185.734 0.000 186.454 44.094 ;
 END
 PORT
  LAYER ME4 ;
  RECT 190.929 1.781 191.269 66.831 ;
 END
 PORT
  LAYER ME4 ;
  RECT 188.927 1.781 189.267 66.831 ;
 END
 PORT
  LAYER ME4 ;
  RECT 189.738 0.000 190.458 44.094 ;
 END
 PORT
  LAYER ME4 ;
  RECT 194.933 1.781 195.273 66.831 ;
 END
 PORT
  LAYER ME4 ;
  RECT 192.931 1.781 193.271 66.831 ;
 END
 PORT
  LAYER ME4 ;
  RECT 193.742 0.000 194.462 44.094 ;
 END
 PORT
  LAYER ME4 ;
  RECT 198.937 1.781 199.277 66.831 ;
 END
 PORT
  LAYER ME4 ;
  RECT 196.935 1.781 197.275 66.831 ;
 END
 PORT
  LAYER ME4 ;
  RECT 197.746 0.000 198.466 44.094 ;
 END
 PORT
  LAYER ME4 ;
  RECT 202.941 1.781 203.281 66.831 ;
 END
 PORT
  LAYER ME4 ;
  RECT 200.939 1.781 201.279 66.831 ;
 END
 PORT
  LAYER ME4 ;
  RECT 201.750 0.000 202.470 44.094 ;
 END
 PORT
  LAYER ME4 ;
  RECT 206.945 1.781 207.285 66.831 ;
 END
 PORT
  LAYER ME4 ;
  RECT 204.943 1.781 205.283 66.831 ;
 END
 PORT
  LAYER ME4 ;
  RECT 205.754 0.000 206.474 44.094 ;
 END
 PORT
  LAYER ME4 ;
  RECT 210.949 1.781 211.289 66.831 ;
 END
 PORT
  LAYER ME4 ;
  RECT 208.947 1.781 209.287 66.831 ;
 END
 PORT
  LAYER ME4 ;
  RECT 209.758 0.000 210.478 44.094 ;
 END
 PORT
  LAYER ME4 ;
  RECT 214.953 1.781 215.293 66.831 ;
 END
 PORT
  LAYER ME4 ;
  RECT 212.951 1.781 213.291 66.831 ;
 END
 PORT
  LAYER ME4 ;
  RECT 213.762 0.000 214.482 44.094 ;
 END
 PORT
  LAYER ME4 ;
  RECT 218.957 1.781 219.297 66.831 ;
 END
 PORT
  LAYER ME4 ;
  RECT 216.955 1.781 217.295 66.831 ;
 END
 PORT
  LAYER ME4 ;
  RECT 217.766 0.000 218.486 44.094 ;
 END
 PORT
  LAYER ME4 ;
  RECT 222.961 1.781 223.301 66.831 ;
 END
 PORT
  LAYER ME4 ;
  RECT 220.959 1.781 221.299 66.831 ;
 END
 PORT
  LAYER ME4 ;
  RECT 221.770 0.000 222.490 44.094 ;
 END
 PORT
  LAYER ME4 ;
  RECT 226.965 1.781 227.305 66.831 ;
 END
 PORT
  LAYER ME4 ;
  RECT 224.963 1.781 225.303 66.831 ;
 END
 PORT
  LAYER ME4 ;
  RECT 225.774 0.000 226.494 44.094 ;
 END
 PORT
  LAYER ME4 ;
  RECT 230.969 1.781 231.309 66.831 ;
 END
 PORT
  LAYER ME4 ;
  RECT 228.967 1.781 229.307 66.831 ;
 END
 PORT
  LAYER ME4 ;
  RECT 229.778 0.000 230.498 44.094 ;
 END
 PORT
  LAYER ME4 ;
  RECT 234.973 1.781 235.313 66.831 ;
 END
 PORT
  LAYER ME4 ;
  RECT 232.971 1.781 233.311 66.831 ;
 END
 PORT
  LAYER ME4 ;
  RECT 233.782 0.000 234.502 44.094 ;
 END
 PORT
  LAYER ME4 ;
  RECT 238.977 1.781 239.317 66.831 ;
 END
 PORT
  LAYER ME4 ;
  RECT 236.975 1.781 237.315 66.831 ;
 END
 PORT
  LAYER ME4 ;
  RECT 237.786 0.000 238.506 44.094 ;
 END
 PORT
  LAYER ME4 ;
  RECT 242.981 1.781 243.321 66.831 ;
 END
 PORT
  LAYER ME4 ;
  RECT 240.979 1.781 241.319 66.831 ;
 END
 PORT
  LAYER ME4 ;
  RECT 241.790 0.000 242.510 44.094 ;
 END
 PORT
  LAYER ME4 ;
  RECT 246.985 1.781 247.325 66.831 ;
 END
 PORT
  LAYER ME4 ;
  RECT 244.983 1.781 245.323 66.831 ;
 END
 PORT
  LAYER ME4 ;
  RECT 245.794 0.000 246.514 44.094 ;
 END
 PORT
  LAYER ME4 ;
  RECT 250.989 1.781 251.329 66.831 ;
 END
 PORT
  LAYER ME4 ;
  RECT 248.987 1.781 249.327 66.831 ;
 END
 PORT
  LAYER ME4 ;
  RECT 249.798 0.000 250.518 44.094 ;
 END
 PORT
  LAYER ME4 ;
  RECT 254.993 1.781 255.333 66.831 ;
 END
 PORT
  LAYER ME4 ;
  RECT 252.991 1.781 253.331 66.831 ;
 END
 PORT
  LAYER ME4 ;
  RECT 253.802 0.000 254.522 44.094 ;
 END
 PORT
  LAYER ME4 ;
  RECT 258.997 1.781 259.337 66.831 ;
 END
 PORT
  LAYER ME4 ;
  RECT 256.995 1.781 257.335 66.831 ;
 END
 PORT
  LAYER ME4 ;
  RECT 257.806 0.000 258.526 44.094 ;
 END
 PORT
  LAYER ME4 ;
  RECT 264.498 0.000 265.218 66.831 ;
 END
 PORT
  LAYER ME4 ;
  RECT 262.458 0.000 263.178 66.831 ;
 END
 PORT
  LAYER ME4 ;
  RECT 259.998 0.000 260.338 66.831 ;
 END
END GND
PIN VCC
  DIRECTION INOUT ;
  USE POWER ;
 PORT
  LAYER ME4 ;
  RECT 298.077 45.394 298.417 66.831 ;
 END
 PORT
  LAYER ME4 ;
  RECT 295.885 0.000 296.605 46.394 ;
 END
 PORT
  LAYER ME4 ;
  RECT 302.081 45.394 302.421 66.831 ;
 END
 PORT
  LAYER ME4 ;
  RECT 299.889 0.000 300.609 46.394 ;
 END
 PORT
  LAYER ME4 ;
  RECT 306.085 45.394 306.425 66.831 ;
 END
 PORT
  LAYER ME4 ;
  RECT 303.893 0.000 304.613 46.394 ;
 END
 PORT
  LAYER ME4 ;
  RECT 310.089 45.394 310.429 66.831 ;
 END
 PORT
  LAYER ME4 ;
  RECT 307.897 0.000 308.617 46.394 ;
 END
 PORT
  LAYER ME4 ;
  RECT 314.093 45.394 314.433 66.831 ;
 END
 PORT
  LAYER ME4 ;
  RECT 311.901 0.000 312.621 46.394 ;
 END
 PORT
  LAYER ME4 ;
  RECT 318.097 45.394 318.437 66.831 ;
 END
 PORT
  LAYER ME4 ;
  RECT 315.905 0.000 316.625 46.394 ;
 END
 PORT
  LAYER ME4 ;
  RECT 322.101 45.394 322.441 66.831 ;
 END
 PORT
  LAYER ME4 ;
  RECT 319.909 0.000 320.629 46.394 ;
 END
 PORT
  LAYER ME4 ;
  RECT 326.105 45.394 326.445 66.831 ;
 END
 PORT
  LAYER ME4 ;
  RECT 323.913 0.000 324.633 46.394 ;
 END
 PORT
  LAYER ME4 ;
  RECT 330.109 45.394 330.449 66.831 ;
 END
 PORT
  LAYER ME4 ;
  RECT 327.917 0.000 328.637 46.394 ;
 END
 PORT
  LAYER ME4 ;
  RECT 334.113 45.394 334.453 66.831 ;
 END
 PORT
  LAYER ME4 ;
  RECT 331.921 0.000 332.641 46.394 ;
 END
 PORT
  LAYER ME4 ;
  RECT 338.117 45.394 338.457 66.831 ;
 END
 PORT
  LAYER ME4 ;
  RECT 335.925 0.000 336.645 46.394 ;
 END
 PORT
  LAYER ME4 ;
  RECT 342.121 45.394 342.461 66.831 ;
 END
 PORT
  LAYER ME4 ;
  RECT 339.929 0.000 340.649 46.394 ;
 END
 PORT
  LAYER ME4 ;
  RECT 346.125 45.394 346.465 66.831 ;
 END
 PORT
  LAYER ME4 ;
  RECT 343.933 0.000 344.653 46.394 ;
 END
 PORT
  LAYER ME4 ;
  RECT 350.129 45.394 350.469 66.831 ;
 END
 PORT
  LAYER ME4 ;
  RECT 347.937 0.000 348.657 46.394 ;
 END
 PORT
  LAYER ME4 ;
  RECT 354.133 45.394 354.473 66.831 ;
 END
 PORT
  LAYER ME4 ;
  RECT 351.941 0.000 352.661 46.394 ;
 END
 PORT
  LAYER ME4 ;
  RECT 358.137 45.394 358.477 66.831 ;
 END
 PORT
  LAYER ME4 ;
  RECT 355.945 0.000 356.665 46.394 ;
 END
 PORT
  LAYER ME4 ;
  RECT 362.141 45.394 362.481 66.831 ;
 END
 PORT
  LAYER ME4 ;
  RECT 359.949 0.000 360.669 46.394 ;
 END
 PORT
  LAYER ME4 ;
  RECT 366.145 45.394 366.485 66.831 ;
 END
 PORT
  LAYER ME4 ;
  RECT 363.953 0.000 364.673 46.394 ;
 END
 PORT
  LAYER ME4 ;
  RECT 370.149 45.394 370.489 66.831 ;
 END
 PORT
  LAYER ME4 ;
  RECT 367.957 0.000 368.677 46.394 ;
 END
 PORT
  LAYER ME4 ;
  RECT 374.153 45.394 374.493 66.831 ;
 END
 PORT
  LAYER ME4 ;
  RECT 371.961 0.000 372.681 46.394 ;
 END
 PORT
  LAYER ME4 ;
  RECT 378.157 45.394 378.497 66.831 ;
 END
 PORT
  LAYER ME4 ;
  RECT 375.965 0.000 376.685 46.394 ;
 END
 PORT
  LAYER ME4 ;
  RECT 382.161 45.394 382.501 66.831 ;
 END
 PORT
  LAYER ME4 ;
  RECT 379.969 0.000 380.689 46.394 ;
 END
 PORT
  LAYER ME4 ;
  RECT 386.165 45.394 386.505 66.831 ;
 END
 PORT
  LAYER ME4 ;
  RECT 383.973 0.000 384.693 46.394 ;
 END
 PORT
  LAYER ME4 ;
  RECT 390.169 45.394 390.509 66.831 ;
 END
 PORT
  LAYER ME4 ;
  RECT 387.977 0.000 388.697 46.394 ;
 END
 PORT
  LAYER ME4 ;
  RECT 394.173 45.394 394.513 66.831 ;
 END
 PORT
  LAYER ME4 ;
  RECT 391.981 0.000 392.701 46.394 ;
 END
 PORT
  LAYER ME4 ;
  RECT 398.177 45.394 398.517 66.831 ;
 END
 PORT
  LAYER ME4 ;
  RECT 395.985 0.000 396.705 46.394 ;
 END
 PORT
  LAYER ME4 ;
  RECT 402.181 45.394 402.521 66.831 ;
 END
 PORT
  LAYER ME4 ;
  RECT 399.989 0.000 400.709 46.394 ;
 END
 PORT
  LAYER ME4 ;
  RECT 406.185 45.394 406.525 66.831 ;
 END
 PORT
  LAYER ME4 ;
  RECT 403.993 0.000 404.713 46.394 ;
 END
 PORT
  LAYER ME4 ;
  RECT 410.189 45.394 410.529 66.831 ;
 END
 PORT
  LAYER ME4 ;
  RECT 407.997 0.000 408.717 46.394 ;
 END
 PORT
  LAYER ME4 ;
  RECT 414.193 45.394 414.533 66.831 ;
 END
 PORT
  LAYER ME4 ;
  RECT 412.001 0.000 412.721 46.394 ;
 END
 PORT
  LAYER ME4 ;
  RECT 418.197 45.394 418.537 66.831 ;
 END
 PORT
  LAYER ME4 ;
  RECT 416.005 0.000 416.725 46.394 ;
 END
 PORT
  LAYER ME4 ;
  RECT 422.201 45.394 422.541 66.831 ;
 END
 PORT
  LAYER ME4 ;
  RECT 420.009 0.000 420.729 46.394 ;
 END
 PORT
  LAYER ME4 ;
  RECT 426.205 45.394 426.545 66.831 ;
 END
 PORT
  LAYER ME4 ;
  RECT 424.013 0.000 424.733 46.394 ;
 END
 PORT
  LAYER ME4 ;
  RECT 430.209 45.394 430.549 66.831 ;
 END
 PORT
  LAYER ME4 ;
  RECT 428.017 0.000 428.737 46.394 ;
 END
 PORT
  LAYER ME4 ;
  RECT 434.213 45.394 434.553 66.831 ;
 END
 PORT
  LAYER ME4 ;
  RECT 432.021 0.000 432.741 46.394 ;
 END
 PORT
  LAYER ME4 ;
  RECT 438.217 45.394 438.557 66.831 ;
 END
 PORT
  LAYER ME4 ;
  RECT 436.025 0.000 436.745 46.394 ;
 END
 PORT
  LAYER ME4 ;
  RECT 442.221 45.394 442.561 66.831 ;
 END
 PORT
  LAYER ME4 ;
  RECT 440.029 0.000 440.749 46.394 ;
 END
 PORT
  LAYER ME4 ;
  RECT 446.225 45.394 446.565 66.831 ;
 END
 PORT
  LAYER ME4 ;
  RECT 444.033 0.000 444.753 46.394 ;
 END
 PORT
  LAYER ME4 ;
  RECT 450.229 45.394 450.569 66.831 ;
 END
 PORT
  LAYER ME4 ;
  RECT 448.037 0.000 448.757 46.394 ;
 END
 PORT
  LAYER ME4 ;
  RECT 454.233 45.394 454.573 66.831 ;
 END
 PORT
  LAYER ME4 ;
  RECT 452.041 0.000 452.761 46.394 ;
 END
 PORT
  LAYER ME4 ;
  RECT 458.237 45.394 458.577 66.831 ;
 END
 PORT
  LAYER ME4 ;
  RECT 456.045 0.000 456.765 46.394 ;
 END
 PORT
  LAYER ME4 ;
  RECT 462.241 45.394 462.581 66.831 ;
 END
 PORT
  LAYER ME4 ;
  RECT 460.049 0.000 460.769 46.394 ;
 END
 PORT
  LAYER ME4 ;
  RECT 466.245 45.394 466.585 66.831 ;
 END
 PORT
  LAYER ME4 ;
  RECT 464.053 0.000 464.773 46.394 ;
 END
 PORT
  LAYER ME4 ;
  RECT 470.249 45.394 470.589 66.831 ;
 END
 PORT
  LAYER ME4 ;
  RECT 468.057 0.000 468.777 46.394 ;
 END
 PORT
  LAYER ME4 ;
  RECT 474.253 45.394 474.593 66.831 ;
 END
 PORT
  LAYER ME4 ;
  RECT 472.061 0.000 472.781 46.394 ;
 END
 PORT
  LAYER ME4 ;
  RECT 478.257 45.394 478.597 66.831 ;
 END
 PORT
  LAYER ME4 ;
  RECT 476.065 0.000 476.785 46.394 ;
 END
 PORT
  LAYER ME4 ;
  RECT 482.261 45.394 482.601 66.831 ;
 END
 PORT
  LAYER ME4 ;
  RECT 480.069 0.000 480.789 46.394 ;
 END
 PORT
  LAYER ME4 ;
  RECT 486.265 45.394 486.605 66.831 ;
 END
 PORT
  LAYER ME4 ;
  RECT 484.073 0.000 484.793 46.394 ;
 END
 PORT
  LAYER ME4 ;
  RECT 490.269 45.394 490.609 66.831 ;
 END
 PORT
  LAYER ME4 ;
  RECT 488.077 0.000 488.797 46.394 ;
 END
 PORT
  LAYER ME4 ;
  RECT 494.273 45.394 494.613 66.831 ;
 END
 PORT
  LAYER ME4 ;
  RECT 492.081 0.000 492.801 46.394 ;
 END
 PORT
  LAYER ME4 ;
  RECT 498.277 45.394 498.617 66.831 ;
 END
 PORT
  LAYER ME4 ;
  RECT 496.085 0.000 496.805 46.394 ;
 END
 PORT
  LAYER ME4 ;
  RECT 502.281 45.394 502.621 66.831 ;
 END
 PORT
  LAYER ME4 ;
  RECT 500.089 0.000 500.809 46.394 ;
 END
 PORT
  LAYER ME4 ;
  RECT 506.285 45.394 506.625 66.831 ;
 END
 PORT
  LAYER ME4 ;
  RECT 504.093 0.000 504.813 46.394 ;
 END
 PORT
  LAYER ME4 ;
  RECT 510.289 45.394 510.629 66.831 ;
 END
 PORT
  LAYER ME4 ;
  RECT 508.097 0.000 508.817 46.394 ;
 END
 PORT
  LAYER ME4 ;
  RECT 514.293 45.394 514.633 66.831 ;
 END
 PORT
  LAYER ME4 ;
  RECT 512.101 0.000 512.821 46.394 ;
 END
 PORT
  LAYER ME4 ;
  RECT 518.297 45.394 518.637 66.831 ;
 END
 PORT
  LAYER ME4 ;
  RECT 516.105 0.000 516.825 46.394 ;
 END
 PORT
  LAYER ME4 ;
  RECT 522.301 45.394 522.641 66.831 ;
 END
 PORT
  LAYER ME4 ;
  RECT 520.109 0.000 520.829 46.394 ;
 END
 PORT
  LAYER ME4 ;
  RECT 526.305 45.394 526.645 66.831 ;
 END
 PORT
  LAYER ME4 ;
  RECT 524.113 0.000 524.833 46.394 ;
 END
 PORT
  LAYER ME4 ;
  RECT 530.309 45.394 530.649 66.831 ;
 END
 PORT
  LAYER ME4 ;
  RECT 528.117 0.000 528.837 46.394 ;
 END
 PORT
  LAYER ME4 ;
  RECT 534.313 45.394 534.653 66.831 ;
 END
 PORT
  LAYER ME4 ;
  RECT 532.121 0.000 532.841 46.394 ;
 END
 PORT
  LAYER ME4 ;
  RECT 538.317 45.394 538.657 66.831 ;
 END
 PORT
  LAYER ME4 ;
  RECT 536.125 0.000 536.845 46.394 ;
 END
 PORT
  LAYER ME4 ;
  RECT 542.321 45.394 542.661 66.831 ;
 END
 PORT
  LAYER ME4 ;
  RECT 540.129 0.000 540.849 46.394 ;
 END
 PORT
  LAYER ME4 ;
  RECT 546.325 45.394 546.665 66.831 ;
 END
 PORT
  LAYER ME4 ;
  RECT 544.133 0.000 544.853 46.394 ;
 END
 PORT
  LAYER ME4 ;
  RECT 550.329 45.394 550.669 66.831 ;
 END
 PORT
  LAYER ME4 ;
  RECT 548.137 0.000 548.857 46.394 ;
 END
 PORT
  LAYER ME4 ;
  RECT 553.111 0.000 553.491 66.831 ;
 END
 PORT
  LAYER ME4 ;
  RECT 278.997 0.000 279.597 66.831 ;
 END
 PORT
  LAYER ME4 ;
  RECT 283.177 0.000 283.897 66.831 ;
 END
 PORT
  LAYER ME4 ;
  RECT 285.287 0.000 286.407 66.831 ;
 END
 PORT
  LAYER ME4 ;
  RECT 291.317 0.000 292.037 66.831 ;
 END
 PORT
  LAYER ME4 ;
  RECT 293.253 1.781 293.633 66.831 ;
 END
 PORT
  LAYER ME4 ;
  RECT 274.767 0.000 275.487 66.831 ;
 END
 PORT
  LAYER ME4 ;
  RECT 272.052 0.000 273.172 66.831 ;
 END
 PORT
  LAYER ME4 ;
  RECT 269.678 0.000 270.398 66.072 ;
 END
 PORT
  LAYER ME4 ;
  RECT 267.638 1.781 268.358 66.831 ;
 END
 PORT
  LAYER ME4 ;
  RECT 0.920 0.000 1.300 66.831 ;
 END
 PORT
  LAYER ME4 ;
  RECT 5.744 45.394 6.084 66.831 ;
 END
 PORT
  LAYER ME4 ;
  RECT 3.552 0.000 4.272 46.394 ;
 END
 PORT
  LAYER ME4 ;
  RECT 9.748 45.394 10.088 66.831 ;
 END
 PORT
  LAYER ME4 ;
  RECT 7.556 0.000 8.276 46.394 ;
 END
 PORT
  LAYER ME4 ;
  RECT 13.752 45.394 14.092 66.831 ;
 END
 PORT
  LAYER ME4 ;
  RECT 11.560 0.000 12.280 46.394 ;
 END
 PORT
  LAYER ME4 ;
  RECT 17.756 45.394 18.096 66.831 ;
 END
 PORT
  LAYER ME4 ;
  RECT 15.564 0.000 16.284 46.394 ;
 END
 PORT
  LAYER ME4 ;
  RECT 21.760 45.394 22.100 66.831 ;
 END
 PORT
  LAYER ME4 ;
  RECT 19.568 0.000 20.288 46.394 ;
 END
 PORT
  LAYER ME4 ;
  RECT 25.764 45.394 26.104 66.831 ;
 END
 PORT
  LAYER ME4 ;
  RECT 23.572 0.000 24.292 46.394 ;
 END
 PORT
  LAYER ME4 ;
  RECT 29.768 45.394 30.108 66.831 ;
 END
 PORT
  LAYER ME4 ;
  RECT 27.576 0.000 28.296 46.394 ;
 END
 PORT
  LAYER ME4 ;
  RECT 33.772 45.394 34.112 66.831 ;
 END
 PORT
  LAYER ME4 ;
  RECT 31.580 0.000 32.300 46.394 ;
 END
 PORT
  LAYER ME4 ;
  RECT 37.776 45.394 38.116 66.831 ;
 END
 PORT
  LAYER ME4 ;
  RECT 35.584 0.000 36.304 46.394 ;
 END
 PORT
  LAYER ME4 ;
  RECT 41.780 45.394 42.120 66.831 ;
 END
 PORT
  LAYER ME4 ;
  RECT 39.588 0.000 40.308 46.394 ;
 END
 PORT
  LAYER ME4 ;
  RECT 45.784 45.394 46.124 66.831 ;
 END
 PORT
  LAYER ME4 ;
  RECT 43.592 0.000 44.312 46.394 ;
 END
 PORT
  LAYER ME4 ;
  RECT 49.788 45.394 50.128 66.831 ;
 END
 PORT
  LAYER ME4 ;
  RECT 47.596 0.000 48.316 46.394 ;
 END
 PORT
  LAYER ME4 ;
  RECT 53.792 45.394 54.132 66.831 ;
 END
 PORT
  LAYER ME4 ;
  RECT 51.600 0.000 52.320 46.394 ;
 END
 PORT
  LAYER ME4 ;
  RECT 57.796 45.394 58.136 66.831 ;
 END
 PORT
  LAYER ME4 ;
  RECT 55.604 0.000 56.324 46.394 ;
 END
 PORT
  LAYER ME4 ;
  RECT 61.800 45.394 62.140 66.831 ;
 END
 PORT
  LAYER ME4 ;
  RECT 59.608 0.000 60.328 46.394 ;
 END
 PORT
  LAYER ME4 ;
  RECT 65.804 45.394 66.144 66.831 ;
 END
 PORT
  LAYER ME4 ;
  RECT 63.612 0.000 64.332 46.394 ;
 END
 PORT
  LAYER ME4 ;
  RECT 69.808 45.394 70.148 66.831 ;
 END
 PORT
  LAYER ME4 ;
  RECT 67.616 0.000 68.336 46.394 ;
 END
 PORT
  LAYER ME4 ;
  RECT 73.812 45.394 74.152 66.831 ;
 END
 PORT
  LAYER ME4 ;
  RECT 71.620 0.000 72.340 46.394 ;
 END
 PORT
  LAYER ME4 ;
  RECT 77.816 45.394 78.156 66.831 ;
 END
 PORT
  LAYER ME4 ;
  RECT 75.624 0.000 76.344 46.394 ;
 END
 PORT
  LAYER ME4 ;
  RECT 81.820 45.394 82.160 66.831 ;
 END
 PORT
  LAYER ME4 ;
  RECT 79.628 0.000 80.348 46.394 ;
 END
 PORT
  LAYER ME4 ;
  RECT 85.824 45.394 86.164 66.831 ;
 END
 PORT
  LAYER ME4 ;
  RECT 83.632 0.000 84.352 46.394 ;
 END
 PORT
  LAYER ME4 ;
  RECT 89.828 45.394 90.168 66.831 ;
 END
 PORT
  LAYER ME4 ;
  RECT 87.636 0.000 88.356 46.394 ;
 END
 PORT
  LAYER ME4 ;
  RECT 93.832 45.394 94.172 66.831 ;
 END
 PORT
  LAYER ME4 ;
  RECT 91.640 0.000 92.360 46.394 ;
 END
 PORT
  LAYER ME4 ;
  RECT 97.836 45.394 98.176 66.831 ;
 END
 PORT
  LAYER ME4 ;
  RECT 95.644 0.000 96.364 46.394 ;
 END
 PORT
  LAYER ME4 ;
  RECT 101.840 45.394 102.180 66.831 ;
 END
 PORT
  LAYER ME4 ;
  RECT 99.648 0.000 100.368 46.394 ;
 END
 PORT
  LAYER ME4 ;
  RECT 105.844 45.394 106.184 66.831 ;
 END
 PORT
  LAYER ME4 ;
  RECT 103.652 0.000 104.372 46.394 ;
 END
 PORT
  LAYER ME4 ;
  RECT 109.848 45.394 110.188 66.831 ;
 END
 PORT
  LAYER ME4 ;
  RECT 107.656 0.000 108.376 46.394 ;
 END
 PORT
  LAYER ME4 ;
  RECT 113.852 45.394 114.192 66.831 ;
 END
 PORT
  LAYER ME4 ;
  RECT 111.660 0.000 112.380 46.394 ;
 END
 PORT
  LAYER ME4 ;
  RECT 117.856 45.394 118.196 66.831 ;
 END
 PORT
  LAYER ME4 ;
  RECT 115.664 0.000 116.384 46.394 ;
 END
 PORT
  LAYER ME4 ;
  RECT 121.860 45.394 122.200 66.831 ;
 END
 PORT
  LAYER ME4 ;
  RECT 119.668 0.000 120.388 46.394 ;
 END
 PORT
  LAYER ME4 ;
  RECT 125.864 45.394 126.204 66.831 ;
 END
 PORT
  LAYER ME4 ;
  RECT 123.672 0.000 124.392 46.394 ;
 END
 PORT
  LAYER ME4 ;
  RECT 129.868 45.394 130.208 66.831 ;
 END
 PORT
  LAYER ME4 ;
  RECT 127.676 0.000 128.396 46.394 ;
 END
 PORT
  LAYER ME4 ;
  RECT 133.872 45.394 134.212 66.831 ;
 END
 PORT
  LAYER ME4 ;
  RECT 131.680 0.000 132.400 46.394 ;
 END
 PORT
  LAYER ME4 ;
  RECT 137.876 45.394 138.216 66.831 ;
 END
 PORT
  LAYER ME4 ;
  RECT 135.684 0.000 136.404 46.394 ;
 END
 PORT
  LAYER ME4 ;
  RECT 141.880 45.394 142.220 66.831 ;
 END
 PORT
  LAYER ME4 ;
  RECT 139.688 0.000 140.408 46.394 ;
 END
 PORT
  LAYER ME4 ;
  RECT 145.884 45.394 146.224 66.831 ;
 END
 PORT
  LAYER ME4 ;
  RECT 143.692 0.000 144.412 46.394 ;
 END
 PORT
  LAYER ME4 ;
  RECT 149.888 45.394 150.228 66.831 ;
 END
 PORT
  LAYER ME4 ;
  RECT 147.696 0.000 148.416 46.394 ;
 END
 PORT
  LAYER ME4 ;
  RECT 153.892 45.394 154.232 66.831 ;
 END
 PORT
  LAYER ME4 ;
  RECT 151.700 0.000 152.420 46.394 ;
 END
 PORT
  LAYER ME4 ;
  RECT 157.896 45.394 158.236 66.831 ;
 END
 PORT
  LAYER ME4 ;
  RECT 155.704 0.000 156.424 46.394 ;
 END
 PORT
  LAYER ME4 ;
  RECT 161.900 45.394 162.240 66.831 ;
 END
 PORT
  LAYER ME4 ;
  RECT 159.708 0.000 160.428 46.394 ;
 END
 PORT
  LAYER ME4 ;
  RECT 165.904 45.394 166.244 66.831 ;
 END
 PORT
  LAYER ME4 ;
  RECT 163.712 0.000 164.432 46.394 ;
 END
 PORT
  LAYER ME4 ;
  RECT 169.908 45.394 170.248 66.831 ;
 END
 PORT
  LAYER ME4 ;
  RECT 167.716 0.000 168.436 46.394 ;
 END
 PORT
  LAYER ME4 ;
  RECT 173.912 45.394 174.252 66.831 ;
 END
 PORT
  LAYER ME4 ;
  RECT 171.720 0.000 172.440 46.394 ;
 END
 PORT
  LAYER ME4 ;
  RECT 177.916 45.394 178.256 66.831 ;
 END
 PORT
  LAYER ME4 ;
  RECT 175.724 0.000 176.444 46.394 ;
 END
 PORT
  LAYER ME4 ;
  RECT 181.920 45.394 182.260 66.831 ;
 END
 PORT
  LAYER ME4 ;
  RECT 179.728 0.000 180.448 46.394 ;
 END
 PORT
  LAYER ME4 ;
  RECT 185.924 45.394 186.264 66.831 ;
 END
 PORT
  LAYER ME4 ;
  RECT 183.732 0.000 184.452 46.394 ;
 END
 PORT
  LAYER ME4 ;
  RECT 189.928 45.394 190.268 66.831 ;
 END
 PORT
  LAYER ME4 ;
  RECT 187.736 0.000 188.456 46.394 ;
 END
 PORT
  LAYER ME4 ;
  RECT 193.932 45.394 194.272 66.831 ;
 END
 PORT
  LAYER ME4 ;
  RECT 191.740 0.000 192.460 46.394 ;
 END
 PORT
  LAYER ME4 ;
  RECT 197.936 45.394 198.276 66.831 ;
 END
 PORT
  LAYER ME4 ;
  RECT 195.744 0.000 196.464 46.394 ;
 END
 PORT
  LAYER ME4 ;
  RECT 201.940 45.394 202.280 66.831 ;
 END
 PORT
  LAYER ME4 ;
  RECT 199.748 0.000 200.468 46.394 ;
 END
 PORT
  LAYER ME4 ;
  RECT 205.944 45.394 206.284 66.831 ;
 END
 PORT
  LAYER ME4 ;
  RECT 203.752 0.000 204.472 46.394 ;
 END
 PORT
  LAYER ME4 ;
  RECT 209.948 45.394 210.288 66.831 ;
 END
 PORT
  LAYER ME4 ;
  RECT 207.756 0.000 208.476 46.394 ;
 END
 PORT
  LAYER ME4 ;
  RECT 213.952 45.394 214.292 66.831 ;
 END
 PORT
  LAYER ME4 ;
  RECT 211.760 0.000 212.480 46.394 ;
 END
 PORT
  LAYER ME4 ;
  RECT 217.956 45.394 218.296 66.831 ;
 END
 PORT
  LAYER ME4 ;
  RECT 215.764 0.000 216.484 46.394 ;
 END
 PORT
  LAYER ME4 ;
  RECT 221.960 45.394 222.300 66.831 ;
 END
 PORT
  LAYER ME4 ;
  RECT 219.768 0.000 220.488 46.394 ;
 END
 PORT
  LAYER ME4 ;
  RECT 225.964 45.394 226.304 66.831 ;
 END
 PORT
  LAYER ME4 ;
  RECT 223.772 0.000 224.492 46.394 ;
 END
 PORT
  LAYER ME4 ;
  RECT 229.968 45.394 230.308 66.831 ;
 END
 PORT
  LAYER ME4 ;
  RECT 227.776 0.000 228.496 46.394 ;
 END
 PORT
  LAYER ME4 ;
  RECT 233.972 45.394 234.312 66.831 ;
 END
 PORT
  LAYER ME4 ;
  RECT 231.780 0.000 232.500 46.394 ;
 END
 PORT
  LAYER ME4 ;
  RECT 237.976 45.394 238.316 66.831 ;
 END
 PORT
  LAYER ME4 ;
  RECT 235.784 0.000 236.504 46.394 ;
 END
 PORT
  LAYER ME4 ;
  RECT 241.980 45.394 242.320 66.831 ;
 END
 PORT
  LAYER ME4 ;
  RECT 239.788 0.000 240.508 46.394 ;
 END
 PORT
  LAYER ME4 ;
  RECT 245.984 45.394 246.324 66.831 ;
 END
 PORT
  LAYER ME4 ;
  RECT 243.792 0.000 244.512 46.394 ;
 END
 PORT
  LAYER ME4 ;
  RECT 249.988 45.394 250.328 66.831 ;
 END
 PORT
  LAYER ME4 ;
  RECT 247.796 0.000 248.516 46.394 ;
 END
 PORT
  LAYER ME4 ;
  RECT 253.992 45.394 254.332 66.831 ;
 END
 PORT
  LAYER ME4 ;
  RECT 251.800 0.000 252.520 46.394 ;
 END
 PORT
  LAYER ME4 ;
  RECT 257.996 45.394 258.336 66.831 ;
 END
 PORT
  LAYER ME4 ;
  RECT 255.804 0.000 256.524 46.394 ;
 END
 PORT
  LAYER ME4 ;
  RECT 265.518 0.000 266.238 66.831 ;
 END
 PORT
  LAYER ME4 ;
  RECT 263.478 0.000 264.198 66.831 ;
 END
 PORT
  LAYER ME4 ;
  RECT 261.358 0.000 262.078 66.831 ;
 END
 PORT
  LAYER ME4 ;
  RECT 260.778 0.000 261.158 66.831 ;
 END
 PORT
  LAYER ME4 ;
  RECT 296.075 47.744 296.415 66.831 ;
 END
 PORT
  LAYER ME4 ;
  RECT 300.079 47.744 300.419 66.831 ;
 END
 PORT
  LAYER ME4 ;
  RECT 304.083 47.744 304.423 66.831 ;
 END
 PORT
  LAYER ME4 ;
  RECT 308.087 47.744 308.427 66.831 ;
 END
 PORT
  LAYER ME4 ;
  RECT 312.091 47.744 312.431 66.831 ;
 END
 PORT
  LAYER ME4 ;
  RECT 316.095 47.744 316.435 66.831 ;
 END
 PORT
  LAYER ME4 ;
  RECT 320.099 47.744 320.439 66.831 ;
 END
 PORT
  LAYER ME4 ;
  RECT 324.103 47.744 324.443 66.831 ;
 END
 PORT
  LAYER ME4 ;
  RECT 328.107 47.744 328.447 66.831 ;
 END
 PORT
  LAYER ME4 ;
  RECT 332.111 47.744 332.451 66.831 ;
 END
 PORT
  LAYER ME4 ;
  RECT 336.115 47.744 336.455 66.831 ;
 END
 PORT
  LAYER ME4 ;
  RECT 340.119 47.744 340.459 66.831 ;
 END
 PORT
  LAYER ME4 ;
  RECT 344.123 47.744 344.463 66.831 ;
 END
 PORT
  LAYER ME4 ;
  RECT 348.127 47.744 348.467 66.831 ;
 END
 PORT
  LAYER ME4 ;
  RECT 352.131 47.744 352.471 66.831 ;
 END
 PORT
  LAYER ME4 ;
  RECT 356.135 47.744 356.475 66.831 ;
 END
 PORT
  LAYER ME4 ;
  RECT 360.139 47.744 360.479 66.831 ;
 END
 PORT
  LAYER ME4 ;
  RECT 364.143 47.744 364.483 66.831 ;
 END
 PORT
  LAYER ME4 ;
  RECT 368.147 47.744 368.487 66.831 ;
 END
 PORT
  LAYER ME4 ;
  RECT 372.151 47.744 372.491 66.831 ;
 END
 PORT
  LAYER ME4 ;
  RECT 376.155 47.744 376.495 66.831 ;
 END
 PORT
  LAYER ME4 ;
  RECT 380.159 47.744 380.499 66.831 ;
 END
 PORT
  LAYER ME4 ;
  RECT 384.163 47.744 384.503 66.831 ;
 END
 PORT
  LAYER ME4 ;
  RECT 388.167 47.744 388.507 66.831 ;
 END
 PORT
  LAYER ME4 ;
  RECT 392.171 47.744 392.511 66.831 ;
 END
 PORT
  LAYER ME4 ;
  RECT 396.175 47.744 396.515 66.831 ;
 END
 PORT
  LAYER ME4 ;
  RECT 400.179 47.744 400.519 66.831 ;
 END
 PORT
  LAYER ME4 ;
  RECT 404.183 47.744 404.523 66.831 ;
 END
 PORT
  LAYER ME4 ;
  RECT 408.187 47.744 408.527 66.831 ;
 END
 PORT
  LAYER ME4 ;
  RECT 412.191 47.744 412.531 66.831 ;
 END
 PORT
  LAYER ME4 ;
  RECT 416.195 47.744 416.535 66.831 ;
 END
 PORT
  LAYER ME4 ;
  RECT 420.199 47.744 420.539 66.831 ;
 END
 PORT
  LAYER ME4 ;
  RECT 424.203 47.744 424.543 66.831 ;
 END
 PORT
  LAYER ME4 ;
  RECT 428.207 47.744 428.547 66.831 ;
 END
 PORT
  LAYER ME4 ;
  RECT 432.211 47.744 432.551 66.831 ;
 END
 PORT
  LAYER ME4 ;
  RECT 436.215 47.744 436.555 66.831 ;
 END
 PORT
  LAYER ME4 ;
  RECT 440.219 47.744 440.559 66.831 ;
 END
 PORT
  LAYER ME4 ;
  RECT 444.223 47.744 444.563 66.831 ;
 END
 PORT
  LAYER ME4 ;
  RECT 448.227 47.744 448.567 66.831 ;
 END
 PORT
  LAYER ME4 ;
  RECT 452.231 47.744 452.571 66.831 ;
 END
 PORT
  LAYER ME4 ;
  RECT 456.235 47.744 456.575 66.831 ;
 END
 PORT
  LAYER ME4 ;
  RECT 460.239 47.744 460.579 66.831 ;
 END
 PORT
  LAYER ME4 ;
  RECT 464.243 47.744 464.583 66.831 ;
 END
 PORT
  LAYER ME4 ;
  RECT 468.247 47.744 468.587 66.831 ;
 END
 PORT
  LAYER ME4 ;
  RECT 472.251 47.744 472.591 66.831 ;
 END
 PORT
  LAYER ME4 ;
  RECT 476.255 47.744 476.595 66.831 ;
 END
 PORT
  LAYER ME4 ;
  RECT 480.259 47.744 480.599 66.831 ;
 END
 PORT
  LAYER ME4 ;
  RECT 484.263 47.744 484.603 66.831 ;
 END
 PORT
  LAYER ME4 ;
  RECT 488.267 47.744 488.607 66.831 ;
 END
 PORT
  LAYER ME4 ;
  RECT 492.271 47.744 492.611 66.831 ;
 END
 PORT
  LAYER ME4 ;
  RECT 496.275 47.744 496.615 66.831 ;
 END
 PORT
  LAYER ME4 ;
  RECT 500.279 47.744 500.619 66.831 ;
 END
 PORT
  LAYER ME4 ;
  RECT 504.283 47.744 504.623 66.831 ;
 END
 PORT
  LAYER ME4 ;
  RECT 508.287 47.744 508.627 66.831 ;
 END
 PORT
  LAYER ME4 ;
  RECT 512.291 47.744 512.631 66.831 ;
 END
 PORT
  LAYER ME4 ;
  RECT 516.295 47.744 516.635 66.831 ;
 END
 PORT
  LAYER ME4 ;
  RECT 520.299 47.744 520.639 66.831 ;
 END
 PORT
  LAYER ME4 ;
  RECT 524.303 47.744 524.643 66.831 ;
 END
 PORT
  LAYER ME4 ;
  RECT 528.307 47.744 528.647 66.831 ;
 END
 PORT
  LAYER ME4 ;
  RECT 532.311 47.744 532.651 66.831 ;
 END
 PORT
  LAYER ME4 ;
  RECT 536.315 47.744 536.655 66.831 ;
 END
 PORT
  LAYER ME4 ;
  RECT 540.319 47.744 540.659 66.831 ;
 END
 PORT
  LAYER ME4 ;
  RECT 544.323 47.744 544.663 66.831 ;
 END
 PORT
  LAYER ME4 ;
  RECT 548.327 47.744 548.667 66.831 ;
 END
 PORT
  LAYER ME4 ;
  RECT 3.742 47.744 4.082 66.831 ;
 END
 PORT
  LAYER ME4 ;
  RECT 7.746 47.744 8.086 66.831 ;
 END
 PORT
  LAYER ME4 ;
  RECT 11.750 47.744 12.090 66.831 ;
 END
 PORT
  LAYER ME4 ;
  RECT 15.754 47.744 16.094 66.831 ;
 END
 PORT
  LAYER ME4 ;
  RECT 19.758 47.744 20.098 66.831 ;
 END
 PORT
  LAYER ME4 ;
  RECT 23.762 47.744 24.102 66.831 ;
 END
 PORT
  LAYER ME4 ;
  RECT 27.766 47.744 28.106 66.831 ;
 END
 PORT
  LAYER ME4 ;
  RECT 31.770 47.744 32.110 66.831 ;
 END
 PORT
  LAYER ME4 ;
  RECT 35.774 47.744 36.114 66.831 ;
 END
 PORT
  LAYER ME4 ;
  RECT 39.778 47.744 40.118 66.831 ;
 END
 PORT
  LAYER ME4 ;
  RECT 43.782 47.744 44.122 66.831 ;
 END
 PORT
  LAYER ME4 ;
  RECT 47.786 47.744 48.126 66.831 ;
 END
 PORT
  LAYER ME4 ;
  RECT 51.790 47.744 52.130 66.831 ;
 END
 PORT
  LAYER ME4 ;
  RECT 55.794 47.744 56.134 66.831 ;
 END
 PORT
  LAYER ME4 ;
  RECT 59.798 47.744 60.138 66.831 ;
 END
 PORT
  LAYER ME4 ;
  RECT 63.802 47.744 64.142 66.831 ;
 END
 PORT
  LAYER ME4 ;
  RECT 67.806 47.744 68.146 66.831 ;
 END
 PORT
  LAYER ME4 ;
  RECT 71.810 47.744 72.150 66.831 ;
 END
 PORT
  LAYER ME4 ;
  RECT 75.814 47.744 76.154 66.831 ;
 END
 PORT
  LAYER ME4 ;
  RECT 79.818 47.744 80.158 66.831 ;
 END
 PORT
  LAYER ME4 ;
  RECT 83.822 47.744 84.162 66.831 ;
 END
 PORT
  LAYER ME4 ;
  RECT 87.826 47.744 88.166 66.831 ;
 END
 PORT
  LAYER ME4 ;
  RECT 91.830 47.744 92.170 66.831 ;
 END
 PORT
  LAYER ME4 ;
  RECT 95.834 47.744 96.174 66.831 ;
 END
 PORT
  LAYER ME4 ;
  RECT 99.838 47.744 100.178 66.831 ;
 END
 PORT
  LAYER ME4 ;
  RECT 103.842 47.744 104.182 66.831 ;
 END
 PORT
  LAYER ME4 ;
  RECT 107.846 47.744 108.186 66.831 ;
 END
 PORT
  LAYER ME4 ;
  RECT 111.850 47.744 112.190 66.831 ;
 END
 PORT
  LAYER ME4 ;
  RECT 115.854 47.744 116.194 66.831 ;
 END
 PORT
  LAYER ME4 ;
  RECT 119.858 47.744 120.198 66.831 ;
 END
 PORT
  LAYER ME4 ;
  RECT 123.862 47.744 124.202 66.831 ;
 END
 PORT
  LAYER ME4 ;
  RECT 127.866 47.744 128.206 66.831 ;
 END
 PORT
  LAYER ME4 ;
  RECT 131.870 47.744 132.210 66.831 ;
 END
 PORT
  LAYER ME4 ;
  RECT 135.874 47.744 136.214 66.831 ;
 END
 PORT
  LAYER ME4 ;
  RECT 139.878 47.744 140.218 66.831 ;
 END
 PORT
  LAYER ME4 ;
  RECT 143.882 47.744 144.222 66.831 ;
 END
 PORT
  LAYER ME4 ;
  RECT 147.886 47.744 148.226 66.831 ;
 END
 PORT
  LAYER ME4 ;
  RECT 151.890 47.744 152.230 66.831 ;
 END
 PORT
  LAYER ME4 ;
  RECT 155.894 47.744 156.234 66.831 ;
 END
 PORT
  LAYER ME4 ;
  RECT 159.898 47.744 160.238 66.831 ;
 END
 PORT
  LAYER ME4 ;
  RECT 163.902 47.744 164.242 66.831 ;
 END
 PORT
  LAYER ME4 ;
  RECT 167.906 47.744 168.246 66.831 ;
 END
 PORT
  LAYER ME4 ;
  RECT 171.910 47.744 172.250 66.831 ;
 END
 PORT
  LAYER ME4 ;
  RECT 175.914 47.744 176.254 66.831 ;
 END
 PORT
  LAYER ME4 ;
  RECT 179.918 47.744 180.258 66.831 ;
 END
 PORT
  LAYER ME4 ;
  RECT 183.922 47.744 184.262 66.831 ;
 END
 PORT
  LAYER ME4 ;
  RECT 187.926 47.744 188.266 66.831 ;
 END
 PORT
  LAYER ME4 ;
  RECT 191.930 47.744 192.270 66.831 ;
 END
 PORT
  LAYER ME4 ;
  RECT 195.934 47.744 196.274 66.831 ;
 END
 PORT
  LAYER ME4 ;
  RECT 199.938 47.744 200.278 66.831 ;
 END
 PORT
  LAYER ME4 ;
  RECT 203.942 47.744 204.282 66.831 ;
 END
 PORT
  LAYER ME4 ;
  RECT 207.946 47.744 208.286 66.831 ;
 END
 PORT
  LAYER ME4 ;
  RECT 211.950 47.744 212.290 66.831 ;
 END
 PORT
  LAYER ME4 ;
  RECT 215.954 47.744 216.294 66.831 ;
 END
 PORT
  LAYER ME4 ;
  RECT 219.958 47.744 220.298 66.831 ;
 END
 PORT
  LAYER ME4 ;
  RECT 223.962 47.744 224.302 66.831 ;
 END
 PORT
  LAYER ME4 ;
  RECT 227.966 47.744 228.306 66.831 ;
 END
 PORT
  LAYER ME4 ;
  RECT 231.970 47.744 232.310 66.831 ;
 END
 PORT
  LAYER ME4 ;
  RECT 235.974 47.744 236.314 66.831 ;
 END
 PORT
  LAYER ME4 ;
  RECT 239.978 47.744 240.318 66.831 ;
 END
 PORT
  LAYER ME4 ;
  RECT 243.982 47.744 244.322 66.831 ;
 END
 PORT
  LAYER ME4 ;
  RECT 247.986 47.744 248.326 66.831 ;
 END
 PORT
  LAYER ME4 ;
  RECT 251.990 47.744 252.330 66.831 ;
 END
 PORT
  LAYER ME4 ;
  RECT 255.994 47.744 256.334 66.831 ;
 END
END VCC
PIN DI63
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 257.286 0.000 257.606 0.600 ;
  LAYER ME3 ;
  RECT 257.286 0.000 257.606 0.600 ;
  LAYER ME2 ;
  RECT 257.286 0.000 257.606 0.600 ;
  LAYER ME1 ;
  RECT 257.286 0.000 257.606 0.600 ;
 END
 ANTENNAPARTIALMETALAREA                  1.058 LAYER ME2 ;
 ANTENNAGATEAREA                          0.072 LAYER ME2 ;
 ANTENNAGATEAREA                          0.072 LAYER ME3 ;
 ANTENNAGATEAREA                          0.072 LAYER ME4 ;
 ANTENNADIFFAREA                          0.160 LAYER ME2 ;
 ANTENNADIFFAREA                          0.160 LAYER ME3 ;
 ANTENNADIFFAREA                          0.160 LAYER ME4 ;
 ANTENNAMAXAREACAR                       21.782 LAYER ME2 ;
 ANTENNAMAXAREACAR                       24.449 LAYER ME3 ;
 ANTENNAMAXAREACAR                       27.116 LAYER ME4 ;
END DI63
PIN DO63
  DIRECTION OUTPUT ;
 PORT
  LAYER ME4 ;
  RECT 256.724 0.000 257.044 0.600 ;
  LAYER ME3 ;
  RECT 256.724 0.000 257.044 0.600 ;
  LAYER ME2 ;
  RECT 256.724 0.000 257.044 0.600 ;
  LAYER ME1 ;
  RECT 256.724 0.000 257.044 0.600 ;
 END
 ANTENNAPARTIALMETALAREA                  5.273 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME3 ;
 ANTENNADIFFAREA                          1.293 LAYER ME4 ;
END DO63
PIN DI62
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 253.282 0.000 253.602 0.600 ;
  LAYER ME3 ;
  RECT 253.282 0.000 253.602 0.600 ;
  LAYER ME2 ;
  RECT 253.282 0.000 253.602 0.600 ;
  LAYER ME1 ;
  RECT 253.282 0.000 253.602 0.600 ;
 END
 ANTENNAPARTIALMETALAREA                  1.058 LAYER ME2 ;
 ANTENNAGATEAREA                          0.072 LAYER ME2 ;
 ANTENNAGATEAREA                          0.072 LAYER ME3 ;
 ANTENNAGATEAREA                          0.072 LAYER ME4 ;
 ANTENNADIFFAREA                          0.160 LAYER ME2 ;
 ANTENNADIFFAREA                          0.160 LAYER ME3 ;
 ANTENNADIFFAREA                          0.160 LAYER ME4 ;
 ANTENNAMAXAREACAR                       21.782 LAYER ME2 ;
 ANTENNAMAXAREACAR                       24.449 LAYER ME3 ;
 ANTENNAMAXAREACAR                       27.116 LAYER ME4 ;
END DI62
PIN DO62
  DIRECTION OUTPUT ;
 PORT
  LAYER ME4 ;
  RECT 252.720 0.000 253.040 0.600 ;
  LAYER ME3 ;
  RECT 252.720 0.000 253.040 0.600 ;
  LAYER ME2 ;
  RECT 252.720 0.000 253.040 0.600 ;
  LAYER ME1 ;
  RECT 252.720 0.000 253.040 0.600 ;
 END
 ANTENNAPARTIALMETALAREA                  5.273 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME3 ;
 ANTENNADIFFAREA                          1.293 LAYER ME4 ;
END DO62
PIN DI61
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 249.278 0.000 249.598 0.600 ;
  LAYER ME3 ;
  RECT 249.278 0.000 249.598 0.600 ;
  LAYER ME2 ;
  RECT 249.278 0.000 249.598 0.600 ;
  LAYER ME1 ;
  RECT 249.278 0.000 249.598 0.600 ;
 END
 ANTENNAPARTIALMETALAREA                  1.058 LAYER ME2 ;
 ANTENNAGATEAREA                          0.072 LAYER ME2 ;
 ANTENNAGATEAREA                          0.072 LAYER ME3 ;
 ANTENNAGATEAREA                          0.072 LAYER ME4 ;
 ANTENNADIFFAREA                          0.160 LAYER ME2 ;
 ANTENNADIFFAREA                          0.160 LAYER ME3 ;
 ANTENNADIFFAREA                          0.160 LAYER ME4 ;
 ANTENNAMAXAREACAR                       21.782 LAYER ME2 ;
 ANTENNAMAXAREACAR                       24.449 LAYER ME3 ;
 ANTENNAMAXAREACAR                       27.116 LAYER ME4 ;
END DI61
PIN DO61
  DIRECTION OUTPUT ;
 PORT
  LAYER ME4 ;
  RECT 248.716 0.000 249.036 0.600 ;
  LAYER ME3 ;
  RECT 248.716 0.000 249.036 0.600 ;
  LAYER ME2 ;
  RECT 248.716 0.000 249.036 0.600 ;
  LAYER ME1 ;
  RECT 248.716 0.000 249.036 0.600 ;
 END
 ANTENNAPARTIALMETALAREA                  5.273 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME3 ;
 ANTENNADIFFAREA                          1.293 LAYER ME4 ;
END DO61
PIN DI60
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 245.274 0.000 245.594 0.600 ;
  LAYER ME3 ;
  RECT 245.274 0.000 245.594 0.600 ;
  LAYER ME2 ;
  RECT 245.274 0.000 245.594 0.600 ;
  LAYER ME1 ;
  RECT 245.274 0.000 245.594 0.600 ;
 END
 ANTENNAPARTIALMETALAREA                  1.058 LAYER ME2 ;
 ANTENNAGATEAREA                          0.072 LAYER ME2 ;
 ANTENNAGATEAREA                          0.072 LAYER ME3 ;
 ANTENNAGATEAREA                          0.072 LAYER ME4 ;
 ANTENNADIFFAREA                          0.160 LAYER ME2 ;
 ANTENNADIFFAREA                          0.160 LAYER ME3 ;
 ANTENNADIFFAREA                          0.160 LAYER ME4 ;
 ANTENNAMAXAREACAR                       21.782 LAYER ME2 ;
 ANTENNAMAXAREACAR                       24.449 LAYER ME3 ;
 ANTENNAMAXAREACAR                       27.116 LAYER ME4 ;
END DI60
PIN DO60
  DIRECTION OUTPUT ;
 PORT
  LAYER ME4 ;
  RECT 244.712 0.000 245.032 0.600 ;
  LAYER ME3 ;
  RECT 244.712 0.000 245.032 0.600 ;
  LAYER ME2 ;
  RECT 244.712 0.000 245.032 0.600 ;
  LAYER ME1 ;
  RECT 244.712 0.000 245.032 0.600 ;
 END
 ANTENNAPARTIALMETALAREA                  5.273 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME3 ;
 ANTENNADIFFAREA                          1.293 LAYER ME4 ;
END DO60
PIN DI59
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 241.270 0.000 241.590 0.600 ;
  LAYER ME3 ;
  RECT 241.270 0.000 241.590 0.600 ;
  LAYER ME2 ;
  RECT 241.270 0.000 241.590 0.600 ;
  LAYER ME1 ;
  RECT 241.270 0.000 241.590 0.600 ;
 END
 ANTENNAPARTIALMETALAREA                  1.058 LAYER ME2 ;
 ANTENNAGATEAREA                          0.072 LAYER ME2 ;
 ANTENNAGATEAREA                          0.072 LAYER ME3 ;
 ANTENNAGATEAREA                          0.072 LAYER ME4 ;
 ANTENNADIFFAREA                          0.160 LAYER ME2 ;
 ANTENNADIFFAREA                          0.160 LAYER ME3 ;
 ANTENNADIFFAREA                          0.160 LAYER ME4 ;
 ANTENNAMAXAREACAR                       21.782 LAYER ME2 ;
 ANTENNAMAXAREACAR                       24.449 LAYER ME3 ;
 ANTENNAMAXAREACAR                       27.116 LAYER ME4 ;
END DI59
PIN DO59
  DIRECTION OUTPUT ;
 PORT
  LAYER ME4 ;
  RECT 240.708 0.000 241.028 0.600 ;
  LAYER ME3 ;
  RECT 240.708 0.000 241.028 0.600 ;
  LAYER ME2 ;
  RECT 240.708 0.000 241.028 0.600 ;
  LAYER ME1 ;
  RECT 240.708 0.000 241.028 0.600 ;
 END
 ANTENNAPARTIALMETALAREA                  5.273 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME3 ;
 ANTENNADIFFAREA                          1.293 LAYER ME4 ;
END DO59
PIN DI58
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 237.266 0.000 237.586 0.600 ;
  LAYER ME3 ;
  RECT 237.266 0.000 237.586 0.600 ;
  LAYER ME2 ;
  RECT 237.266 0.000 237.586 0.600 ;
  LAYER ME1 ;
  RECT 237.266 0.000 237.586 0.600 ;
 END
 ANTENNAPARTIALMETALAREA                  1.058 LAYER ME2 ;
 ANTENNAGATEAREA                          0.072 LAYER ME2 ;
 ANTENNAGATEAREA                          0.072 LAYER ME3 ;
 ANTENNAGATEAREA                          0.072 LAYER ME4 ;
 ANTENNADIFFAREA                          0.160 LAYER ME2 ;
 ANTENNADIFFAREA                          0.160 LAYER ME3 ;
 ANTENNADIFFAREA                          0.160 LAYER ME4 ;
 ANTENNAMAXAREACAR                       21.782 LAYER ME2 ;
 ANTENNAMAXAREACAR                       24.449 LAYER ME3 ;
 ANTENNAMAXAREACAR                       27.116 LAYER ME4 ;
END DI58
PIN DO58
  DIRECTION OUTPUT ;
 PORT
  LAYER ME4 ;
  RECT 236.704 0.000 237.024 0.600 ;
  LAYER ME3 ;
  RECT 236.704 0.000 237.024 0.600 ;
  LAYER ME2 ;
  RECT 236.704 0.000 237.024 0.600 ;
  LAYER ME1 ;
  RECT 236.704 0.000 237.024 0.600 ;
 END
 ANTENNAPARTIALMETALAREA                  5.273 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME3 ;
 ANTENNADIFFAREA                          1.293 LAYER ME4 ;
END DO58
PIN DI57
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 233.262 0.000 233.582 0.600 ;
  LAYER ME3 ;
  RECT 233.262 0.000 233.582 0.600 ;
  LAYER ME2 ;
  RECT 233.262 0.000 233.582 0.600 ;
  LAYER ME1 ;
  RECT 233.262 0.000 233.582 0.600 ;
 END
 ANTENNAPARTIALMETALAREA                  1.058 LAYER ME2 ;
 ANTENNAGATEAREA                          0.072 LAYER ME2 ;
 ANTENNAGATEAREA                          0.072 LAYER ME3 ;
 ANTENNAGATEAREA                          0.072 LAYER ME4 ;
 ANTENNADIFFAREA                          0.160 LAYER ME2 ;
 ANTENNADIFFAREA                          0.160 LAYER ME3 ;
 ANTENNADIFFAREA                          0.160 LAYER ME4 ;
 ANTENNAMAXAREACAR                       21.782 LAYER ME2 ;
 ANTENNAMAXAREACAR                       24.449 LAYER ME3 ;
 ANTENNAMAXAREACAR                       27.116 LAYER ME4 ;
END DI57
PIN DO57
  DIRECTION OUTPUT ;
 PORT
  LAYER ME4 ;
  RECT 232.700 0.000 233.020 0.600 ;
  LAYER ME3 ;
  RECT 232.700 0.000 233.020 0.600 ;
  LAYER ME2 ;
  RECT 232.700 0.000 233.020 0.600 ;
  LAYER ME1 ;
  RECT 232.700 0.000 233.020 0.600 ;
 END
 ANTENNAPARTIALMETALAREA                  5.273 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME3 ;
 ANTENNADIFFAREA                          1.293 LAYER ME4 ;
END DO57
PIN DI56
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 228.696 0.000 229.016 0.600 ;
  LAYER ME3 ;
  RECT 228.696 0.000 229.016 0.600 ;
  LAYER ME2 ;
  RECT 228.696 0.000 229.016 0.600 ;
  LAYER ME1 ;
  RECT 228.696 0.000 229.016 0.600 ;
 END
 ANTENNAPARTIALMETALAREA                  0.346 LAYER ME1 ;
 ANTENNAPARTIALMETALAREA                  1.466 LAYER ME2 ;
 ANTENNAPARTIALMETALAREA                  0.508 LAYER ME3 ;
 ANTENNAGATEAREA                          0.072 LAYER ME3 ;
 ANTENNAGATEAREA                          0.072 LAYER ME4 ;
 ANTENNADIFFAREA                          0.218 LAYER ME1 ;
 ANTENNADIFFAREA                          0.218 LAYER ME2 ;
 ANTENNADIFFAREA                          0.218 LAYER ME3 ;
 ANTENNADIFFAREA                          0.218 LAYER ME4 ;
 ANTENNAMAXAREACAR                       17.267 LAYER ME3 ;
 ANTENNAMAXAREACAR                       19.933 LAYER ME4 ;
END DI56
PIN DO56
  DIRECTION OUTPUT ;
 PORT
  LAYER ME4 ;
  RECT 229.258 0.000 229.578 0.600 ;
  LAYER ME3 ;
  RECT 229.258 0.000 229.578 0.600 ;
  LAYER ME2 ;
  RECT 229.258 0.000 229.578 0.600 ;
  LAYER ME1 ;
  RECT 229.258 0.000 229.578 0.600 ;
 END
 ANTENNAPARTIALMETALAREA                  5.602 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME3 ;
 ANTENNADIFFAREA                          1.293 LAYER ME4 ;
END DO56
PIN WEB7
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 227.256 0.000 227.576 0.600 ;
  LAYER ME3 ;
  RECT 227.256 0.000 227.576 0.600 ;
  LAYER ME2 ;
  RECT 227.256 0.000 227.576 0.600 ;
  LAYER ME1 ;
  RECT 227.256 0.000 227.576 0.600 ;
 END
 ANTENNAPARTIALMETALAREA                  1.036 LAYER ME2 ;
 ANTENNAGATEAREA                          0.288 LAYER ME2 ;
 ANTENNAGATEAREA                          0.288 LAYER ME3 ;
 ANTENNAGATEAREA                          0.288 LAYER ME4 ;
 ANTENNADIFFAREA                          0.206 LAYER ME2 ;
 ANTENNADIFFAREA                          0.206 LAYER ME3 ;
 ANTENNADIFFAREA                          0.206 LAYER ME4 ;
 ANTENNAMAXAREACAR                        5.844 LAYER ME2 ;
 ANTENNAMAXAREACAR                        6.511 LAYER ME3 ;
 ANTENNAMAXAREACAR                        7.178 LAYER ME4 ;
END WEB7
PIN DI55
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 225.254 0.000 225.574 0.600 ;
  LAYER ME3 ;
  RECT 225.254 0.000 225.574 0.600 ;
  LAYER ME2 ;
  RECT 225.254 0.000 225.574 0.600 ;
  LAYER ME1 ;
  RECT 225.254 0.000 225.574 0.600 ;
 END
 ANTENNAPARTIALMETALAREA                  1.058 LAYER ME2 ;
 ANTENNAGATEAREA                          0.072 LAYER ME2 ;
 ANTENNAGATEAREA                          0.072 LAYER ME3 ;
 ANTENNAGATEAREA                          0.072 LAYER ME4 ;
 ANTENNADIFFAREA                          0.160 LAYER ME2 ;
 ANTENNADIFFAREA                          0.160 LAYER ME3 ;
 ANTENNADIFFAREA                          0.160 LAYER ME4 ;
 ANTENNAMAXAREACAR                       21.782 LAYER ME2 ;
 ANTENNAMAXAREACAR                       24.449 LAYER ME3 ;
 ANTENNAMAXAREACAR                       27.116 LAYER ME4 ;
END DI55
PIN DO55
  DIRECTION OUTPUT ;
 PORT
  LAYER ME4 ;
  RECT 224.692 0.000 225.012 0.600 ;
  LAYER ME3 ;
  RECT 224.692 0.000 225.012 0.600 ;
  LAYER ME2 ;
  RECT 224.692 0.000 225.012 0.600 ;
  LAYER ME1 ;
  RECT 224.692 0.000 225.012 0.600 ;
 END
 ANTENNAPARTIALMETALAREA                  5.273 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME3 ;
 ANTENNADIFFAREA                          1.293 LAYER ME4 ;
END DO55
PIN DI54
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 221.250 0.000 221.570 0.600 ;
  LAYER ME3 ;
  RECT 221.250 0.000 221.570 0.600 ;
  LAYER ME2 ;
  RECT 221.250 0.000 221.570 0.600 ;
  LAYER ME1 ;
  RECT 221.250 0.000 221.570 0.600 ;
 END
 ANTENNAPARTIALMETALAREA                  1.058 LAYER ME2 ;
 ANTENNAGATEAREA                          0.072 LAYER ME2 ;
 ANTENNAGATEAREA                          0.072 LAYER ME3 ;
 ANTENNAGATEAREA                          0.072 LAYER ME4 ;
 ANTENNADIFFAREA                          0.160 LAYER ME2 ;
 ANTENNADIFFAREA                          0.160 LAYER ME3 ;
 ANTENNADIFFAREA                          0.160 LAYER ME4 ;
 ANTENNAMAXAREACAR                       21.782 LAYER ME2 ;
 ANTENNAMAXAREACAR                       24.449 LAYER ME3 ;
 ANTENNAMAXAREACAR                       27.116 LAYER ME4 ;
END DI54
PIN DO54
  DIRECTION OUTPUT ;
 PORT
  LAYER ME4 ;
  RECT 220.688 0.000 221.008 0.600 ;
  LAYER ME3 ;
  RECT 220.688 0.000 221.008 0.600 ;
  LAYER ME2 ;
  RECT 220.688 0.000 221.008 0.600 ;
  LAYER ME1 ;
  RECT 220.688 0.000 221.008 0.600 ;
 END
 ANTENNAPARTIALMETALAREA                  5.273 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME3 ;
 ANTENNADIFFAREA                          1.293 LAYER ME4 ;
END DO54
PIN DI53
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 217.246 0.000 217.566 0.600 ;
  LAYER ME3 ;
  RECT 217.246 0.000 217.566 0.600 ;
  LAYER ME2 ;
  RECT 217.246 0.000 217.566 0.600 ;
  LAYER ME1 ;
  RECT 217.246 0.000 217.566 0.600 ;
 END
 ANTENNAPARTIALMETALAREA                  1.058 LAYER ME2 ;
 ANTENNAGATEAREA                          0.072 LAYER ME2 ;
 ANTENNAGATEAREA                          0.072 LAYER ME3 ;
 ANTENNAGATEAREA                          0.072 LAYER ME4 ;
 ANTENNADIFFAREA                          0.160 LAYER ME2 ;
 ANTENNADIFFAREA                          0.160 LAYER ME3 ;
 ANTENNADIFFAREA                          0.160 LAYER ME4 ;
 ANTENNAMAXAREACAR                       21.782 LAYER ME2 ;
 ANTENNAMAXAREACAR                       24.449 LAYER ME3 ;
 ANTENNAMAXAREACAR                       27.116 LAYER ME4 ;
END DI53
PIN DO53
  DIRECTION OUTPUT ;
 PORT
  LAYER ME4 ;
  RECT 216.684 0.000 217.004 0.600 ;
  LAYER ME3 ;
  RECT 216.684 0.000 217.004 0.600 ;
  LAYER ME2 ;
  RECT 216.684 0.000 217.004 0.600 ;
  LAYER ME1 ;
  RECT 216.684 0.000 217.004 0.600 ;
 END
 ANTENNAPARTIALMETALAREA                  5.273 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME3 ;
 ANTENNADIFFAREA                          1.293 LAYER ME4 ;
END DO53
PIN DI52
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 213.242 0.000 213.562 0.600 ;
  LAYER ME3 ;
  RECT 213.242 0.000 213.562 0.600 ;
  LAYER ME2 ;
  RECT 213.242 0.000 213.562 0.600 ;
  LAYER ME1 ;
  RECT 213.242 0.000 213.562 0.600 ;
 END
 ANTENNAPARTIALMETALAREA                  1.058 LAYER ME2 ;
 ANTENNAGATEAREA                          0.072 LAYER ME2 ;
 ANTENNAGATEAREA                          0.072 LAYER ME3 ;
 ANTENNAGATEAREA                          0.072 LAYER ME4 ;
 ANTENNADIFFAREA                          0.160 LAYER ME2 ;
 ANTENNADIFFAREA                          0.160 LAYER ME3 ;
 ANTENNADIFFAREA                          0.160 LAYER ME4 ;
 ANTENNAMAXAREACAR                       21.782 LAYER ME2 ;
 ANTENNAMAXAREACAR                       24.449 LAYER ME3 ;
 ANTENNAMAXAREACAR                       27.116 LAYER ME4 ;
END DI52
PIN DO52
  DIRECTION OUTPUT ;
 PORT
  LAYER ME4 ;
  RECT 212.680 0.000 213.000 0.600 ;
  LAYER ME3 ;
  RECT 212.680 0.000 213.000 0.600 ;
  LAYER ME2 ;
  RECT 212.680 0.000 213.000 0.600 ;
  LAYER ME1 ;
  RECT 212.680 0.000 213.000 0.600 ;
 END
 ANTENNAPARTIALMETALAREA                  5.273 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME3 ;
 ANTENNADIFFAREA                          1.293 LAYER ME4 ;
END DO52
PIN DI51
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 209.238 0.000 209.558 0.600 ;
  LAYER ME3 ;
  RECT 209.238 0.000 209.558 0.600 ;
  LAYER ME2 ;
  RECT 209.238 0.000 209.558 0.600 ;
  LAYER ME1 ;
  RECT 209.238 0.000 209.558 0.600 ;
 END
 ANTENNAPARTIALMETALAREA                  1.058 LAYER ME2 ;
 ANTENNAGATEAREA                          0.072 LAYER ME2 ;
 ANTENNAGATEAREA                          0.072 LAYER ME3 ;
 ANTENNAGATEAREA                          0.072 LAYER ME4 ;
 ANTENNADIFFAREA                          0.160 LAYER ME2 ;
 ANTENNADIFFAREA                          0.160 LAYER ME3 ;
 ANTENNADIFFAREA                          0.160 LAYER ME4 ;
 ANTENNAMAXAREACAR                       21.782 LAYER ME2 ;
 ANTENNAMAXAREACAR                       24.449 LAYER ME3 ;
 ANTENNAMAXAREACAR                       27.116 LAYER ME4 ;
END DI51
PIN DO51
  DIRECTION OUTPUT ;
 PORT
  LAYER ME4 ;
  RECT 208.676 0.000 208.996 0.600 ;
  LAYER ME3 ;
  RECT 208.676 0.000 208.996 0.600 ;
  LAYER ME2 ;
  RECT 208.676 0.000 208.996 0.600 ;
  LAYER ME1 ;
  RECT 208.676 0.000 208.996 0.600 ;
 END
 ANTENNAPARTIALMETALAREA                  5.273 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME3 ;
 ANTENNADIFFAREA                          1.293 LAYER ME4 ;
END DO51
PIN DI50
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 205.234 0.000 205.554 0.600 ;
  LAYER ME3 ;
  RECT 205.234 0.000 205.554 0.600 ;
  LAYER ME2 ;
  RECT 205.234 0.000 205.554 0.600 ;
  LAYER ME1 ;
  RECT 205.234 0.000 205.554 0.600 ;
 END
 ANTENNAPARTIALMETALAREA                  1.058 LAYER ME2 ;
 ANTENNAGATEAREA                          0.072 LAYER ME2 ;
 ANTENNAGATEAREA                          0.072 LAYER ME3 ;
 ANTENNAGATEAREA                          0.072 LAYER ME4 ;
 ANTENNADIFFAREA                          0.160 LAYER ME2 ;
 ANTENNADIFFAREA                          0.160 LAYER ME3 ;
 ANTENNADIFFAREA                          0.160 LAYER ME4 ;
 ANTENNAMAXAREACAR                       21.782 LAYER ME2 ;
 ANTENNAMAXAREACAR                       24.449 LAYER ME3 ;
 ANTENNAMAXAREACAR                       27.116 LAYER ME4 ;
END DI50
PIN DO50
  DIRECTION OUTPUT ;
 PORT
  LAYER ME4 ;
  RECT 204.672 0.000 204.992 0.600 ;
  LAYER ME3 ;
  RECT 204.672 0.000 204.992 0.600 ;
  LAYER ME2 ;
  RECT 204.672 0.000 204.992 0.600 ;
  LAYER ME1 ;
  RECT 204.672 0.000 204.992 0.600 ;
 END
 ANTENNAPARTIALMETALAREA                  5.273 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME3 ;
 ANTENNADIFFAREA                          1.293 LAYER ME4 ;
END DO50
PIN DI49
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 201.230 0.000 201.550 0.600 ;
  LAYER ME3 ;
  RECT 201.230 0.000 201.550 0.600 ;
  LAYER ME2 ;
  RECT 201.230 0.000 201.550 0.600 ;
  LAYER ME1 ;
  RECT 201.230 0.000 201.550 0.600 ;
 END
 ANTENNAPARTIALMETALAREA                  1.058 LAYER ME2 ;
 ANTENNAGATEAREA                          0.072 LAYER ME2 ;
 ANTENNAGATEAREA                          0.072 LAYER ME3 ;
 ANTENNAGATEAREA                          0.072 LAYER ME4 ;
 ANTENNADIFFAREA                          0.160 LAYER ME2 ;
 ANTENNADIFFAREA                          0.160 LAYER ME3 ;
 ANTENNADIFFAREA                          0.160 LAYER ME4 ;
 ANTENNAMAXAREACAR                       21.782 LAYER ME2 ;
 ANTENNAMAXAREACAR                       24.449 LAYER ME3 ;
 ANTENNAMAXAREACAR                       27.116 LAYER ME4 ;
END DI49
PIN DO49
  DIRECTION OUTPUT ;
 PORT
  LAYER ME4 ;
  RECT 200.668 0.000 200.988 0.600 ;
  LAYER ME3 ;
  RECT 200.668 0.000 200.988 0.600 ;
  LAYER ME2 ;
  RECT 200.668 0.000 200.988 0.600 ;
  LAYER ME1 ;
  RECT 200.668 0.000 200.988 0.600 ;
 END
 ANTENNAPARTIALMETALAREA                  5.273 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME3 ;
 ANTENNADIFFAREA                          1.293 LAYER ME4 ;
END DO49
PIN DI48
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 196.664 0.000 196.984 0.600 ;
  LAYER ME3 ;
  RECT 196.664 0.000 196.984 0.600 ;
  LAYER ME2 ;
  RECT 196.664 0.000 196.984 0.600 ;
  LAYER ME1 ;
  RECT 196.664 0.000 196.984 0.600 ;
 END
 ANTENNAPARTIALMETALAREA                  0.346 LAYER ME1 ;
 ANTENNAPARTIALMETALAREA                  1.466 LAYER ME2 ;
 ANTENNAPARTIALMETALAREA                  0.508 LAYER ME3 ;
 ANTENNAGATEAREA                          0.072 LAYER ME3 ;
 ANTENNAGATEAREA                          0.072 LAYER ME4 ;
 ANTENNADIFFAREA                          0.218 LAYER ME1 ;
 ANTENNADIFFAREA                          0.218 LAYER ME2 ;
 ANTENNADIFFAREA                          0.218 LAYER ME3 ;
 ANTENNADIFFAREA                          0.218 LAYER ME4 ;
 ANTENNAMAXAREACAR                       17.267 LAYER ME3 ;
 ANTENNAMAXAREACAR                       19.933 LAYER ME4 ;
END DI48
PIN DO48
  DIRECTION OUTPUT ;
 PORT
  LAYER ME4 ;
  RECT 197.226 0.000 197.546 0.600 ;
  LAYER ME3 ;
  RECT 197.226 0.000 197.546 0.600 ;
  LAYER ME2 ;
  RECT 197.226 0.000 197.546 0.600 ;
  LAYER ME1 ;
  RECT 197.226 0.000 197.546 0.600 ;
 END
 ANTENNAPARTIALMETALAREA                  5.602 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME3 ;
 ANTENNADIFFAREA                          1.293 LAYER ME4 ;
END DO48
PIN WEB6
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 195.224 0.000 195.544 0.600 ;
  LAYER ME3 ;
  RECT 195.224 0.000 195.544 0.600 ;
  LAYER ME2 ;
  RECT 195.224 0.000 195.544 0.600 ;
  LAYER ME1 ;
  RECT 195.224 0.000 195.544 0.600 ;
 END
 ANTENNAPARTIALMETALAREA                  1.036 LAYER ME2 ;
 ANTENNAGATEAREA                          0.288 LAYER ME2 ;
 ANTENNAGATEAREA                          0.288 LAYER ME3 ;
 ANTENNAGATEAREA                          0.288 LAYER ME4 ;
 ANTENNADIFFAREA                          0.206 LAYER ME2 ;
 ANTENNADIFFAREA                          0.206 LAYER ME3 ;
 ANTENNADIFFAREA                          0.206 LAYER ME4 ;
 ANTENNAMAXAREACAR                        5.844 LAYER ME2 ;
 ANTENNAMAXAREACAR                        6.511 LAYER ME3 ;
 ANTENNAMAXAREACAR                        7.178 LAYER ME4 ;
END WEB6
PIN DI47
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 193.222 0.000 193.542 0.600 ;
  LAYER ME3 ;
  RECT 193.222 0.000 193.542 0.600 ;
  LAYER ME2 ;
  RECT 193.222 0.000 193.542 0.600 ;
  LAYER ME1 ;
  RECT 193.222 0.000 193.542 0.600 ;
 END
 ANTENNAPARTIALMETALAREA                  1.058 LAYER ME2 ;
 ANTENNAGATEAREA                          0.072 LAYER ME2 ;
 ANTENNAGATEAREA                          0.072 LAYER ME3 ;
 ANTENNAGATEAREA                          0.072 LAYER ME4 ;
 ANTENNADIFFAREA                          0.160 LAYER ME2 ;
 ANTENNADIFFAREA                          0.160 LAYER ME3 ;
 ANTENNADIFFAREA                          0.160 LAYER ME4 ;
 ANTENNAMAXAREACAR                       21.782 LAYER ME2 ;
 ANTENNAMAXAREACAR                       24.449 LAYER ME3 ;
 ANTENNAMAXAREACAR                       27.116 LAYER ME4 ;
END DI47
PIN DO47
  DIRECTION OUTPUT ;
 PORT
  LAYER ME4 ;
  RECT 192.660 0.000 192.980 0.600 ;
  LAYER ME3 ;
  RECT 192.660 0.000 192.980 0.600 ;
  LAYER ME2 ;
  RECT 192.660 0.000 192.980 0.600 ;
  LAYER ME1 ;
  RECT 192.660 0.000 192.980 0.600 ;
 END
 ANTENNAPARTIALMETALAREA                  5.273 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME3 ;
 ANTENNADIFFAREA                          1.293 LAYER ME4 ;
END DO47
PIN DI46
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 189.218 0.000 189.538 0.600 ;
  LAYER ME3 ;
  RECT 189.218 0.000 189.538 0.600 ;
  LAYER ME2 ;
  RECT 189.218 0.000 189.538 0.600 ;
  LAYER ME1 ;
  RECT 189.218 0.000 189.538 0.600 ;
 END
 ANTENNAPARTIALMETALAREA                  1.058 LAYER ME2 ;
 ANTENNAGATEAREA                          0.072 LAYER ME2 ;
 ANTENNAGATEAREA                          0.072 LAYER ME3 ;
 ANTENNAGATEAREA                          0.072 LAYER ME4 ;
 ANTENNADIFFAREA                          0.160 LAYER ME2 ;
 ANTENNADIFFAREA                          0.160 LAYER ME3 ;
 ANTENNADIFFAREA                          0.160 LAYER ME4 ;
 ANTENNAMAXAREACAR                       21.782 LAYER ME2 ;
 ANTENNAMAXAREACAR                       24.449 LAYER ME3 ;
 ANTENNAMAXAREACAR                       27.116 LAYER ME4 ;
END DI46
PIN DO46
  DIRECTION OUTPUT ;
 PORT
  LAYER ME4 ;
  RECT 188.656 0.000 188.976 0.600 ;
  LAYER ME3 ;
  RECT 188.656 0.000 188.976 0.600 ;
  LAYER ME2 ;
  RECT 188.656 0.000 188.976 0.600 ;
  LAYER ME1 ;
  RECT 188.656 0.000 188.976 0.600 ;
 END
 ANTENNAPARTIALMETALAREA                  5.273 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME3 ;
 ANTENNADIFFAREA                          1.293 LAYER ME4 ;
END DO46
PIN DI45
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 185.214 0.000 185.534 0.600 ;
  LAYER ME3 ;
  RECT 185.214 0.000 185.534 0.600 ;
  LAYER ME2 ;
  RECT 185.214 0.000 185.534 0.600 ;
  LAYER ME1 ;
  RECT 185.214 0.000 185.534 0.600 ;
 END
 ANTENNAPARTIALMETALAREA                  1.058 LAYER ME2 ;
 ANTENNAGATEAREA                          0.072 LAYER ME2 ;
 ANTENNAGATEAREA                          0.072 LAYER ME3 ;
 ANTENNAGATEAREA                          0.072 LAYER ME4 ;
 ANTENNADIFFAREA                          0.160 LAYER ME2 ;
 ANTENNADIFFAREA                          0.160 LAYER ME3 ;
 ANTENNADIFFAREA                          0.160 LAYER ME4 ;
 ANTENNAMAXAREACAR                       21.782 LAYER ME2 ;
 ANTENNAMAXAREACAR                       24.449 LAYER ME3 ;
 ANTENNAMAXAREACAR                       27.116 LAYER ME4 ;
END DI45
PIN DO45
  DIRECTION OUTPUT ;
 PORT
  LAYER ME4 ;
  RECT 184.652 0.000 184.972 0.600 ;
  LAYER ME3 ;
  RECT 184.652 0.000 184.972 0.600 ;
  LAYER ME2 ;
  RECT 184.652 0.000 184.972 0.600 ;
  LAYER ME1 ;
  RECT 184.652 0.000 184.972 0.600 ;
 END
 ANTENNAPARTIALMETALAREA                  5.273 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME3 ;
 ANTENNADIFFAREA                          1.293 LAYER ME4 ;
END DO45
PIN DI44
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 181.210 0.000 181.530 0.600 ;
  LAYER ME3 ;
  RECT 181.210 0.000 181.530 0.600 ;
  LAYER ME2 ;
  RECT 181.210 0.000 181.530 0.600 ;
  LAYER ME1 ;
  RECT 181.210 0.000 181.530 0.600 ;
 END
 ANTENNAPARTIALMETALAREA                  1.058 LAYER ME2 ;
 ANTENNAGATEAREA                          0.072 LAYER ME2 ;
 ANTENNAGATEAREA                          0.072 LAYER ME3 ;
 ANTENNAGATEAREA                          0.072 LAYER ME4 ;
 ANTENNADIFFAREA                          0.160 LAYER ME2 ;
 ANTENNADIFFAREA                          0.160 LAYER ME3 ;
 ANTENNADIFFAREA                          0.160 LAYER ME4 ;
 ANTENNAMAXAREACAR                       21.782 LAYER ME2 ;
 ANTENNAMAXAREACAR                       24.449 LAYER ME3 ;
 ANTENNAMAXAREACAR                       27.116 LAYER ME4 ;
END DI44
PIN DO44
  DIRECTION OUTPUT ;
 PORT
  LAYER ME4 ;
  RECT 180.648 0.000 180.968 0.600 ;
  LAYER ME3 ;
  RECT 180.648 0.000 180.968 0.600 ;
  LAYER ME2 ;
  RECT 180.648 0.000 180.968 0.600 ;
  LAYER ME1 ;
  RECT 180.648 0.000 180.968 0.600 ;
 END
 ANTENNAPARTIALMETALAREA                  5.273 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME3 ;
 ANTENNADIFFAREA                          1.293 LAYER ME4 ;
END DO44
PIN DI43
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 177.206 0.000 177.526 0.600 ;
  LAYER ME3 ;
  RECT 177.206 0.000 177.526 0.600 ;
  LAYER ME2 ;
  RECT 177.206 0.000 177.526 0.600 ;
  LAYER ME1 ;
  RECT 177.206 0.000 177.526 0.600 ;
 END
 ANTENNAPARTIALMETALAREA                  1.058 LAYER ME2 ;
 ANTENNAGATEAREA                          0.072 LAYER ME2 ;
 ANTENNAGATEAREA                          0.072 LAYER ME3 ;
 ANTENNAGATEAREA                          0.072 LAYER ME4 ;
 ANTENNADIFFAREA                          0.160 LAYER ME2 ;
 ANTENNADIFFAREA                          0.160 LAYER ME3 ;
 ANTENNADIFFAREA                          0.160 LAYER ME4 ;
 ANTENNAMAXAREACAR                       21.782 LAYER ME2 ;
 ANTENNAMAXAREACAR                       24.449 LAYER ME3 ;
 ANTENNAMAXAREACAR                       27.116 LAYER ME4 ;
END DI43
PIN DO43
  DIRECTION OUTPUT ;
 PORT
  LAYER ME4 ;
  RECT 176.644 0.000 176.964 0.600 ;
  LAYER ME3 ;
  RECT 176.644 0.000 176.964 0.600 ;
  LAYER ME2 ;
  RECT 176.644 0.000 176.964 0.600 ;
  LAYER ME1 ;
  RECT 176.644 0.000 176.964 0.600 ;
 END
 ANTENNAPARTIALMETALAREA                  5.273 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME3 ;
 ANTENNADIFFAREA                          1.293 LAYER ME4 ;
END DO43
PIN DI42
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 173.202 0.000 173.522 0.600 ;
  LAYER ME3 ;
  RECT 173.202 0.000 173.522 0.600 ;
  LAYER ME2 ;
  RECT 173.202 0.000 173.522 0.600 ;
  LAYER ME1 ;
  RECT 173.202 0.000 173.522 0.600 ;
 END
 ANTENNAPARTIALMETALAREA                  1.058 LAYER ME2 ;
 ANTENNAGATEAREA                          0.072 LAYER ME2 ;
 ANTENNAGATEAREA                          0.072 LAYER ME3 ;
 ANTENNAGATEAREA                          0.072 LAYER ME4 ;
 ANTENNADIFFAREA                          0.160 LAYER ME2 ;
 ANTENNADIFFAREA                          0.160 LAYER ME3 ;
 ANTENNADIFFAREA                          0.160 LAYER ME4 ;
 ANTENNAMAXAREACAR                       21.782 LAYER ME2 ;
 ANTENNAMAXAREACAR                       24.449 LAYER ME3 ;
 ANTENNAMAXAREACAR                       27.116 LAYER ME4 ;
END DI42
PIN DO42
  DIRECTION OUTPUT ;
 PORT
  LAYER ME4 ;
  RECT 172.640 0.000 172.960 0.600 ;
  LAYER ME3 ;
  RECT 172.640 0.000 172.960 0.600 ;
  LAYER ME2 ;
  RECT 172.640 0.000 172.960 0.600 ;
  LAYER ME1 ;
  RECT 172.640 0.000 172.960 0.600 ;
 END
 ANTENNAPARTIALMETALAREA                  5.273 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME3 ;
 ANTENNADIFFAREA                          1.293 LAYER ME4 ;
END DO42
PIN DI41
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 169.198 0.000 169.518 0.600 ;
  LAYER ME3 ;
  RECT 169.198 0.000 169.518 0.600 ;
  LAYER ME2 ;
  RECT 169.198 0.000 169.518 0.600 ;
  LAYER ME1 ;
  RECT 169.198 0.000 169.518 0.600 ;
 END
 ANTENNAPARTIALMETALAREA                  1.058 LAYER ME2 ;
 ANTENNAGATEAREA                          0.072 LAYER ME2 ;
 ANTENNAGATEAREA                          0.072 LAYER ME3 ;
 ANTENNAGATEAREA                          0.072 LAYER ME4 ;
 ANTENNADIFFAREA                          0.160 LAYER ME2 ;
 ANTENNADIFFAREA                          0.160 LAYER ME3 ;
 ANTENNADIFFAREA                          0.160 LAYER ME4 ;
 ANTENNAMAXAREACAR                       21.782 LAYER ME2 ;
 ANTENNAMAXAREACAR                       24.449 LAYER ME3 ;
 ANTENNAMAXAREACAR                       27.116 LAYER ME4 ;
END DI41
PIN DO41
  DIRECTION OUTPUT ;
 PORT
  LAYER ME4 ;
  RECT 168.636 0.000 168.956 0.600 ;
  LAYER ME3 ;
  RECT 168.636 0.000 168.956 0.600 ;
  LAYER ME2 ;
  RECT 168.636 0.000 168.956 0.600 ;
  LAYER ME1 ;
  RECT 168.636 0.000 168.956 0.600 ;
 END
 ANTENNAPARTIALMETALAREA                  5.273 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME3 ;
 ANTENNADIFFAREA                          1.293 LAYER ME4 ;
END DO41
PIN DI40
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 164.632 0.000 164.952 0.600 ;
  LAYER ME3 ;
  RECT 164.632 0.000 164.952 0.600 ;
  LAYER ME2 ;
  RECT 164.632 0.000 164.952 0.600 ;
  LAYER ME1 ;
  RECT 164.632 0.000 164.952 0.600 ;
 END
 ANTENNAPARTIALMETALAREA                  0.346 LAYER ME1 ;
 ANTENNAPARTIALMETALAREA                  1.466 LAYER ME2 ;
 ANTENNAPARTIALMETALAREA                  0.508 LAYER ME3 ;
 ANTENNAGATEAREA                          0.072 LAYER ME3 ;
 ANTENNAGATEAREA                          0.072 LAYER ME4 ;
 ANTENNADIFFAREA                          0.218 LAYER ME1 ;
 ANTENNADIFFAREA                          0.218 LAYER ME2 ;
 ANTENNADIFFAREA                          0.218 LAYER ME3 ;
 ANTENNADIFFAREA                          0.218 LAYER ME4 ;
 ANTENNAMAXAREACAR                       17.267 LAYER ME3 ;
 ANTENNAMAXAREACAR                       19.933 LAYER ME4 ;
END DI40
PIN DO40
  DIRECTION OUTPUT ;
 PORT
  LAYER ME4 ;
  RECT 165.194 0.000 165.514 0.600 ;
  LAYER ME3 ;
  RECT 165.194 0.000 165.514 0.600 ;
  LAYER ME2 ;
  RECT 165.194 0.000 165.514 0.600 ;
  LAYER ME1 ;
  RECT 165.194 0.000 165.514 0.600 ;
 END
 ANTENNAPARTIALMETALAREA                  5.602 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME3 ;
 ANTENNADIFFAREA                          1.293 LAYER ME4 ;
END DO40
PIN WEB5
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 163.192 0.000 163.512 0.600 ;
  LAYER ME3 ;
  RECT 163.192 0.000 163.512 0.600 ;
  LAYER ME2 ;
  RECT 163.192 0.000 163.512 0.600 ;
  LAYER ME1 ;
  RECT 163.192 0.000 163.512 0.600 ;
 END
 ANTENNAPARTIALMETALAREA                  1.036 LAYER ME2 ;
 ANTENNAGATEAREA                          0.288 LAYER ME2 ;
 ANTENNAGATEAREA                          0.288 LAYER ME3 ;
 ANTENNAGATEAREA                          0.288 LAYER ME4 ;
 ANTENNADIFFAREA                          0.206 LAYER ME2 ;
 ANTENNADIFFAREA                          0.206 LAYER ME3 ;
 ANTENNADIFFAREA                          0.206 LAYER ME4 ;
 ANTENNAMAXAREACAR                        5.844 LAYER ME2 ;
 ANTENNAMAXAREACAR                        6.511 LAYER ME3 ;
 ANTENNAMAXAREACAR                        7.178 LAYER ME4 ;
END WEB5
PIN DI39
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 161.190 0.000 161.510 0.600 ;
  LAYER ME3 ;
  RECT 161.190 0.000 161.510 0.600 ;
  LAYER ME2 ;
  RECT 161.190 0.000 161.510 0.600 ;
  LAYER ME1 ;
  RECT 161.190 0.000 161.510 0.600 ;
 END
 ANTENNAPARTIALMETALAREA                  1.058 LAYER ME2 ;
 ANTENNAGATEAREA                          0.072 LAYER ME2 ;
 ANTENNAGATEAREA                          0.072 LAYER ME3 ;
 ANTENNAGATEAREA                          0.072 LAYER ME4 ;
 ANTENNADIFFAREA                          0.160 LAYER ME2 ;
 ANTENNADIFFAREA                          0.160 LAYER ME3 ;
 ANTENNADIFFAREA                          0.160 LAYER ME4 ;
 ANTENNAMAXAREACAR                       21.782 LAYER ME2 ;
 ANTENNAMAXAREACAR                       24.449 LAYER ME3 ;
 ANTENNAMAXAREACAR                       27.116 LAYER ME4 ;
END DI39
PIN DO39
  DIRECTION OUTPUT ;
 PORT
  LAYER ME4 ;
  RECT 160.628 0.000 160.948 0.600 ;
  LAYER ME3 ;
  RECT 160.628 0.000 160.948 0.600 ;
  LAYER ME2 ;
  RECT 160.628 0.000 160.948 0.600 ;
  LAYER ME1 ;
  RECT 160.628 0.000 160.948 0.600 ;
 END
 ANTENNAPARTIALMETALAREA                  5.273 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME3 ;
 ANTENNADIFFAREA                          1.293 LAYER ME4 ;
END DO39
PIN DI38
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 157.186 0.000 157.506 0.600 ;
  LAYER ME3 ;
  RECT 157.186 0.000 157.506 0.600 ;
  LAYER ME2 ;
  RECT 157.186 0.000 157.506 0.600 ;
  LAYER ME1 ;
  RECT 157.186 0.000 157.506 0.600 ;
 END
 ANTENNAPARTIALMETALAREA                  1.058 LAYER ME2 ;
 ANTENNAGATEAREA                          0.072 LAYER ME2 ;
 ANTENNAGATEAREA                          0.072 LAYER ME3 ;
 ANTENNAGATEAREA                          0.072 LAYER ME4 ;
 ANTENNADIFFAREA                          0.160 LAYER ME2 ;
 ANTENNADIFFAREA                          0.160 LAYER ME3 ;
 ANTENNADIFFAREA                          0.160 LAYER ME4 ;
 ANTENNAMAXAREACAR                       21.782 LAYER ME2 ;
 ANTENNAMAXAREACAR                       24.449 LAYER ME3 ;
 ANTENNAMAXAREACAR                       27.116 LAYER ME4 ;
END DI38
PIN DO38
  DIRECTION OUTPUT ;
 PORT
  LAYER ME4 ;
  RECT 156.624 0.000 156.944 0.600 ;
  LAYER ME3 ;
  RECT 156.624 0.000 156.944 0.600 ;
  LAYER ME2 ;
  RECT 156.624 0.000 156.944 0.600 ;
  LAYER ME1 ;
  RECT 156.624 0.000 156.944 0.600 ;
 END
 ANTENNAPARTIALMETALAREA                  5.273 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME3 ;
 ANTENNADIFFAREA                          1.293 LAYER ME4 ;
END DO38
PIN DI37
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 153.182 0.000 153.502 0.600 ;
  LAYER ME3 ;
  RECT 153.182 0.000 153.502 0.600 ;
  LAYER ME2 ;
  RECT 153.182 0.000 153.502 0.600 ;
  LAYER ME1 ;
  RECT 153.182 0.000 153.502 0.600 ;
 END
 ANTENNAPARTIALMETALAREA                  1.058 LAYER ME2 ;
 ANTENNAGATEAREA                          0.072 LAYER ME2 ;
 ANTENNAGATEAREA                          0.072 LAYER ME3 ;
 ANTENNAGATEAREA                          0.072 LAYER ME4 ;
 ANTENNADIFFAREA                          0.160 LAYER ME2 ;
 ANTENNADIFFAREA                          0.160 LAYER ME3 ;
 ANTENNADIFFAREA                          0.160 LAYER ME4 ;
 ANTENNAMAXAREACAR                       21.782 LAYER ME2 ;
 ANTENNAMAXAREACAR                       24.449 LAYER ME3 ;
 ANTENNAMAXAREACAR                       27.116 LAYER ME4 ;
END DI37
PIN DO37
  DIRECTION OUTPUT ;
 PORT
  LAYER ME4 ;
  RECT 152.620 0.000 152.940 0.600 ;
  LAYER ME3 ;
  RECT 152.620 0.000 152.940 0.600 ;
  LAYER ME2 ;
  RECT 152.620 0.000 152.940 0.600 ;
  LAYER ME1 ;
  RECT 152.620 0.000 152.940 0.600 ;
 END
 ANTENNAPARTIALMETALAREA                  5.273 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME3 ;
 ANTENNADIFFAREA                          1.293 LAYER ME4 ;
END DO37
PIN DI36
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 149.178 0.000 149.498 0.600 ;
  LAYER ME3 ;
  RECT 149.178 0.000 149.498 0.600 ;
  LAYER ME2 ;
  RECT 149.178 0.000 149.498 0.600 ;
  LAYER ME1 ;
  RECT 149.178 0.000 149.498 0.600 ;
 END
 ANTENNAPARTIALMETALAREA                  1.058 LAYER ME2 ;
 ANTENNAGATEAREA                          0.072 LAYER ME2 ;
 ANTENNAGATEAREA                          0.072 LAYER ME3 ;
 ANTENNAGATEAREA                          0.072 LAYER ME4 ;
 ANTENNADIFFAREA                          0.160 LAYER ME2 ;
 ANTENNADIFFAREA                          0.160 LAYER ME3 ;
 ANTENNADIFFAREA                          0.160 LAYER ME4 ;
 ANTENNAMAXAREACAR                       21.782 LAYER ME2 ;
 ANTENNAMAXAREACAR                       24.449 LAYER ME3 ;
 ANTENNAMAXAREACAR                       27.116 LAYER ME4 ;
END DI36
PIN DO36
  DIRECTION OUTPUT ;
 PORT
  LAYER ME4 ;
  RECT 148.616 0.000 148.936 0.600 ;
  LAYER ME3 ;
  RECT 148.616 0.000 148.936 0.600 ;
  LAYER ME2 ;
  RECT 148.616 0.000 148.936 0.600 ;
  LAYER ME1 ;
  RECT 148.616 0.000 148.936 0.600 ;
 END
 ANTENNAPARTIALMETALAREA                  5.273 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME3 ;
 ANTENNADIFFAREA                          1.293 LAYER ME4 ;
END DO36
PIN DI35
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 145.174 0.000 145.494 0.600 ;
  LAYER ME3 ;
  RECT 145.174 0.000 145.494 0.600 ;
  LAYER ME2 ;
  RECT 145.174 0.000 145.494 0.600 ;
  LAYER ME1 ;
  RECT 145.174 0.000 145.494 0.600 ;
 END
 ANTENNAPARTIALMETALAREA                  1.058 LAYER ME2 ;
 ANTENNAGATEAREA                          0.072 LAYER ME2 ;
 ANTENNAGATEAREA                          0.072 LAYER ME3 ;
 ANTENNAGATEAREA                          0.072 LAYER ME4 ;
 ANTENNADIFFAREA                          0.160 LAYER ME2 ;
 ANTENNADIFFAREA                          0.160 LAYER ME3 ;
 ANTENNADIFFAREA                          0.160 LAYER ME4 ;
 ANTENNAMAXAREACAR                       21.782 LAYER ME2 ;
 ANTENNAMAXAREACAR                       24.449 LAYER ME3 ;
 ANTENNAMAXAREACAR                       27.116 LAYER ME4 ;
END DI35
PIN DO35
  DIRECTION OUTPUT ;
 PORT
  LAYER ME4 ;
  RECT 144.612 0.000 144.932 0.600 ;
  LAYER ME3 ;
  RECT 144.612 0.000 144.932 0.600 ;
  LAYER ME2 ;
  RECT 144.612 0.000 144.932 0.600 ;
  LAYER ME1 ;
  RECT 144.612 0.000 144.932 0.600 ;
 END
 ANTENNAPARTIALMETALAREA                  5.273 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME3 ;
 ANTENNADIFFAREA                          1.293 LAYER ME4 ;
END DO35
PIN DI34
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 141.170 0.000 141.490 0.600 ;
  LAYER ME3 ;
  RECT 141.170 0.000 141.490 0.600 ;
  LAYER ME2 ;
  RECT 141.170 0.000 141.490 0.600 ;
  LAYER ME1 ;
  RECT 141.170 0.000 141.490 0.600 ;
 END
 ANTENNAPARTIALMETALAREA                  1.058 LAYER ME2 ;
 ANTENNAGATEAREA                          0.072 LAYER ME2 ;
 ANTENNAGATEAREA                          0.072 LAYER ME3 ;
 ANTENNAGATEAREA                          0.072 LAYER ME4 ;
 ANTENNADIFFAREA                          0.160 LAYER ME2 ;
 ANTENNADIFFAREA                          0.160 LAYER ME3 ;
 ANTENNADIFFAREA                          0.160 LAYER ME4 ;
 ANTENNAMAXAREACAR                       21.782 LAYER ME2 ;
 ANTENNAMAXAREACAR                       24.449 LAYER ME3 ;
 ANTENNAMAXAREACAR                       27.116 LAYER ME4 ;
END DI34
PIN DO34
  DIRECTION OUTPUT ;
 PORT
  LAYER ME4 ;
  RECT 140.608 0.000 140.928 0.600 ;
  LAYER ME3 ;
  RECT 140.608 0.000 140.928 0.600 ;
  LAYER ME2 ;
  RECT 140.608 0.000 140.928 0.600 ;
  LAYER ME1 ;
  RECT 140.608 0.000 140.928 0.600 ;
 END
 ANTENNAPARTIALMETALAREA                  5.273 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME3 ;
 ANTENNADIFFAREA                          1.293 LAYER ME4 ;
END DO34
PIN DI33
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 137.166 0.000 137.486 0.600 ;
  LAYER ME3 ;
  RECT 137.166 0.000 137.486 0.600 ;
  LAYER ME2 ;
  RECT 137.166 0.000 137.486 0.600 ;
  LAYER ME1 ;
  RECT 137.166 0.000 137.486 0.600 ;
 END
 ANTENNAPARTIALMETALAREA                  1.058 LAYER ME2 ;
 ANTENNAGATEAREA                          0.072 LAYER ME2 ;
 ANTENNAGATEAREA                          0.072 LAYER ME3 ;
 ANTENNAGATEAREA                          0.072 LAYER ME4 ;
 ANTENNADIFFAREA                          0.160 LAYER ME2 ;
 ANTENNADIFFAREA                          0.160 LAYER ME3 ;
 ANTENNADIFFAREA                          0.160 LAYER ME4 ;
 ANTENNAMAXAREACAR                       21.782 LAYER ME2 ;
 ANTENNAMAXAREACAR                       24.449 LAYER ME3 ;
 ANTENNAMAXAREACAR                       27.116 LAYER ME4 ;
END DI33
PIN DO33
  DIRECTION OUTPUT ;
 PORT
  LAYER ME4 ;
  RECT 136.604 0.000 136.924 0.600 ;
  LAYER ME3 ;
  RECT 136.604 0.000 136.924 0.600 ;
  LAYER ME2 ;
  RECT 136.604 0.000 136.924 0.600 ;
  LAYER ME1 ;
  RECT 136.604 0.000 136.924 0.600 ;
 END
 ANTENNAPARTIALMETALAREA                  5.273 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME3 ;
 ANTENNADIFFAREA                          1.293 LAYER ME4 ;
END DO33
PIN DI32
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 132.600 0.000 132.920 0.600 ;
  LAYER ME3 ;
  RECT 132.600 0.000 132.920 0.600 ;
  LAYER ME2 ;
  RECT 132.600 0.000 132.920 0.600 ;
  LAYER ME1 ;
  RECT 132.600 0.000 132.920 0.600 ;
 END
 ANTENNAPARTIALMETALAREA                  0.346 LAYER ME1 ;
 ANTENNAPARTIALMETALAREA                  1.466 LAYER ME2 ;
 ANTENNAPARTIALMETALAREA                  0.508 LAYER ME3 ;
 ANTENNAGATEAREA                          0.072 LAYER ME3 ;
 ANTENNAGATEAREA                          0.072 LAYER ME4 ;
 ANTENNADIFFAREA                          0.218 LAYER ME1 ;
 ANTENNADIFFAREA                          0.218 LAYER ME2 ;
 ANTENNADIFFAREA                          0.218 LAYER ME3 ;
 ANTENNADIFFAREA                          0.218 LAYER ME4 ;
 ANTENNAMAXAREACAR                       17.267 LAYER ME3 ;
 ANTENNAMAXAREACAR                       19.933 LAYER ME4 ;
END DI32
PIN DO32
  DIRECTION OUTPUT ;
 PORT
  LAYER ME4 ;
  RECT 133.162 0.000 133.482 0.600 ;
  LAYER ME3 ;
  RECT 133.162 0.000 133.482 0.600 ;
  LAYER ME2 ;
  RECT 133.162 0.000 133.482 0.600 ;
  LAYER ME1 ;
  RECT 133.162 0.000 133.482 0.600 ;
 END
 ANTENNAPARTIALMETALAREA                  5.602 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME3 ;
 ANTENNADIFFAREA                          1.293 LAYER ME4 ;
END DO32
PIN WEB4
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 131.160 0.000 131.480 0.600 ;
  LAYER ME3 ;
  RECT 131.160 0.000 131.480 0.600 ;
  LAYER ME2 ;
  RECT 131.160 0.000 131.480 0.600 ;
  LAYER ME1 ;
  RECT 131.160 0.000 131.480 0.600 ;
 END
 ANTENNAPARTIALMETALAREA                  1.036 LAYER ME2 ;
 ANTENNAGATEAREA                          0.288 LAYER ME2 ;
 ANTENNAGATEAREA                          0.288 LAYER ME3 ;
 ANTENNAGATEAREA                          0.288 LAYER ME4 ;
 ANTENNADIFFAREA                          0.206 LAYER ME2 ;
 ANTENNADIFFAREA                          0.206 LAYER ME3 ;
 ANTENNADIFFAREA                          0.206 LAYER ME4 ;
 ANTENNAMAXAREACAR                        5.844 LAYER ME2 ;
 ANTENNAMAXAREACAR                        6.511 LAYER ME3 ;
 ANTENNAMAXAREACAR                        7.178 LAYER ME4 ;
END WEB4
PIN DI31
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 129.158 0.000 129.478 0.600 ;
  LAYER ME3 ;
  RECT 129.158 0.000 129.478 0.600 ;
  LAYER ME2 ;
  RECT 129.158 0.000 129.478 0.600 ;
  LAYER ME1 ;
  RECT 129.158 0.000 129.478 0.600 ;
 END
 ANTENNAPARTIALMETALAREA                  1.058 LAYER ME2 ;
 ANTENNAGATEAREA                          0.072 LAYER ME2 ;
 ANTENNAGATEAREA                          0.072 LAYER ME3 ;
 ANTENNAGATEAREA                          0.072 LAYER ME4 ;
 ANTENNADIFFAREA                          0.160 LAYER ME2 ;
 ANTENNADIFFAREA                          0.160 LAYER ME3 ;
 ANTENNADIFFAREA                          0.160 LAYER ME4 ;
 ANTENNAMAXAREACAR                       21.782 LAYER ME2 ;
 ANTENNAMAXAREACAR                       24.449 LAYER ME3 ;
 ANTENNAMAXAREACAR                       27.116 LAYER ME4 ;
END DI31
PIN DO31
  DIRECTION OUTPUT ;
 PORT
  LAYER ME4 ;
  RECT 128.596 0.000 128.916 0.600 ;
  LAYER ME3 ;
  RECT 128.596 0.000 128.916 0.600 ;
  LAYER ME2 ;
  RECT 128.596 0.000 128.916 0.600 ;
  LAYER ME1 ;
  RECT 128.596 0.000 128.916 0.600 ;
 END
 ANTENNAPARTIALMETALAREA                  5.273 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME3 ;
 ANTENNADIFFAREA                          1.293 LAYER ME4 ;
END DO31
PIN DI30
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 125.154 0.000 125.474 0.600 ;
  LAYER ME3 ;
  RECT 125.154 0.000 125.474 0.600 ;
  LAYER ME2 ;
  RECT 125.154 0.000 125.474 0.600 ;
  LAYER ME1 ;
  RECT 125.154 0.000 125.474 0.600 ;
 END
 ANTENNAPARTIALMETALAREA                  1.058 LAYER ME2 ;
 ANTENNAGATEAREA                          0.072 LAYER ME2 ;
 ANTENNAGATEAREA                          0.072 LAYER ME3 ;
 ANTENNAGATEAREA                          0.072 LAYER ME4 ;
 ANTENNADIFFAREA                          0.160 LAYER ME2 ;
 ANTENNADIFFAREA                          0.160 LAYER ME3 ;
 ANTENNADIFFAREA                          0.160 LAYER ME4 ;
 ANTENNAMAXAREACAR                       21.782 LAYER ME2 ;
 ANTENNAMAXAREACAR                       24.449 LAYER ME3 ;
 ANTENNAMAXAREACAR                       27.116 LAYER ME4 ;
END DI30
PIN DO30
  DIRECTION OUTPUT ;
 PORT
  LAYER ME4 ;
  RECT 124.592 0.000 124.912 0.600 ;
  LAYER ME3 ;
  RECT 124.592 0.000 124.912 0.600 ;
  LAYER ME2 ;
  RECT 124.592 0.000 124.912 0.600 ;
  LAYER ME1 ;
  RECT 124.592 0.000 124.912 0.600 ;
 END
 ANTENNAPARTIALMETALAREA                  5.273 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME3 ;
 ANTENNADIFFAREA                          1.293 LAYER ME4 ;
END DO30
PIN DI29
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 121.150 0.000 121.470 0.600 ;
  LAYER ME3 ;
  RECT 121.150 0.000 121.470 0.600 ;
  LAYER ME2 ;
  RECT 121.150 0.000 121.470 0.600 ;
  LAYER ME1 ;
  RECT 121.150 0.000 121.470 0.600 ;
 END
 ANTENNAPARTIALMETALAREA                  1.058 LAYER ME2 ;
 ANTENNAGATEAREA                          0.072 LAYER ME2 ;
 ANTENNAGATEAREA                          0.072 LAYER ME3 ;
 ANTENNAGATEAREA                          0.072 LAYER ME4 ;
 ANTENNADIFFAREA                          0.160 LAYER ME2 ;
 ANTENNADIFFAREA                          0.160 LAYER ME3 ;
 ANTENNADIFFAREA                          0.160 LAYER ME4 ;
 ANTENNAMAXAREACAR                       21.782 LAYER ME2 ;
 ANTENNAMAXAREACAR                       24.449 LAYER ME3 ;
 ANTENNAMAXAREACAR                       27.116 LAYER ME4 ;
END DI29
PIN DO29
  DIRECTION OUTPUT ;
 PORT
  LAYER ME4 ;
  RECT 120.588 0.000 120.908 0.600 ;
  LAYER ME3 ;
  RECT 120.588 0.000 120.908 0.600 ;
  LAYER ME2 ;
  RECT 120.588 0.000 120.908 0.600 ;
  LAYER ME1 ;
  RECT 120.588 0.000 120.908 0.600 ;
 END
 ANTENNAPARTIALMETALAREA                  5.273 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME3 ;
 ANTENNADIFFAREA                          1.293 LAYER ME4 ;
END DO29
PIN DI28
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 117.146 0.000 117.466 0.600 ;
  LAYER ME3 ;
  RECT 117.146 0.000 117.466 0.600 ;
  LAYER ME2 ;
  RECT 117.146 0.000 117.466 0.600 ;
  LAYER ME1 ;
  RECT 117.146 0.000 117.466 0.600 ;
 END
 ANTENNAPARTIALMETALAREA                  1.058 LAYER ME2 ;
 ANTENNAGATEAREA                          0.072 LAYER ME2 ;
 ANTENNAGATEAREA                          0.072 LAYER ME3 ;
 ANTENNAGATEAREA                          0.072 LAYER ME4 ;
 ANTENNADIFFAREA                          0.160 LAYER ME2 ;
 ANTENNADIFFAREA                          0.160 LAYER ME3 ;
 ANTENNADIFFAREA                          0.160 LAYER ME4 ;
 ANTENNAMAXAREACAR                       21.782 LAYER ME2 ;
 ANTENNAMAXAREACAR                       24.449 LAYER ME3 ;
 ANTENNAMAXAREACAR                       27.116 LAYER ME4 ;
END DI28
PIN DO28
  DIRECTION OUTPUT ;
 PORT
  LAYER ME4 ;
  RECT 116.584 0.000 116.904 0.600 ;
  LAYER ME3 ;
  RECT 116.584 0.000 116.904 0.600 ;
  LAYER ME2 ;
  RECT 116.584 0.000 116.904 0.600 ;
  LAYER ME1 ;
  RECT 116.584 0.000 116.904 0.600 ;
 END
 ANTENNAPARTIALMETALAREA                  5.273 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME3 ;
 ANTENNADIFFAREA                          1.293 LAYER ME4 ;
END DO28
PIN DI27
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 113.142 0.000 113.462 0.600 ;
  LAYER ME3 ;
  RECT 113.142 0.000 113.462 0.600 ;
  LAYER ME2 ;
  RECT 113.142 0.000 113.462 0.600 ;
  LAYER ME1 ;
  RECT 113.142 0.000 113.462 0.600 ;
 END
 ANTENNAPARTIALMETALAREA                  1.058 LAYER ME2 ;
 ANTENNAGATEAREA                          0.072 LAYER ME2 ;
 ANTENNAGATEAREA                          0.072 LAYER ME3 ;
 ANTENNAGATEAREA                          0.072 LAYER ME4 ;
 ANTENNADIFFAREA                          0.160 LAYER ME2 ;
 ANTENNADIFFAREA                          0.160 LAYER ME3 ;
 ANTENNADIFFAREA                          0.160 LAYER ME4 ;
 ANTENNAMAXAREACAR                       21.782 LAYER ME2 ;
 ANTENNAMAXAREACAR                       24.449 LAYER ME3 ;
 ANTENNAMAXAREACAR                       27.116 LAYER ME4 ;
END DI27
PIN DO27
  DIRECTION OUTPUT ;
 PORT
  LAYER ME4 ;
  RECT 112.580 0.000 112.900 0.600 ;
  LAYER ME3 ;
  RECT 112.580 0.000 112.900 0.600 ;
  LAYER ME2 ;
  RECT 112.580 0.000 112.900 0.600 ;
  LAYER ME1 ;
  RECT 112.580 0.000 112.900 0.600 ;
 END
 ANTENNAPARTIALMETALAREA                  5.273 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME3 ;
 ANTENNADIFFAREA                          1.293 LAYER ME4 ;
END DO27
PIN DI26
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 109.138 0.000 109.458 0.600 ;
  LAYER ME3 ;
  RECT 109.138 0.000 109.458 0.600 ;
  LAYER ME2 ;
  RECT 109.138 0.000 109.458 0.600 ;
  LAYER ME1 ;
  RECT 109.138 0.000 109.458 0.600 ;
 END
 ANTENNAPARTIALMETALAREA                  1.058 LAYER ME2 ;
 ANTENNAGATEAREA                          0.072 LAYER ME2 ;
 ANTENNAGATEAREA                          0.072 LAYER ME3 ;
 ANTENNAGATEAREA                          0.072 LAYER ME4 ;
 ANTENNADIFFAREA                          0.160 LAYER ME2 ;
 ANTENNADIFFAREA                          0.160 LAYER ME3 ;
 ANTENNADIFFAREA                          0.160 LAYER ME4 ;
 ANTENNAMAXAREACAR                       21.782 LAYER ME2 ;
 ANTENNAMAXAREACAR                       24.449 LAYER ME3 ;
 ANTENNAMAXAREACAR                       27.116 LAYER ME4 ;
END DI26
PIN DO26
  DIRECTION OUTPUT ;
 PORT
  LAYER ME4 ;
  RECT 108.576 0.000 108.896 0.600 ;
  LAYER ME3 ;
  RECT 108.576 0.000 108.896 0.600 ;
  LAYER ME2 ;
  RECT 108.576 0.000 108.896 0.600 ;
  LAYER ME1 ;
  RECT 108.576 0.000 108.896 0.600 ;
 END
 ANTENNAPARTIALMETALAREA                  5.273 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME3 ;
 ANTENNADIFFAREA                          1.293 LAYER ME4 ;
END DO26
PIN DI25
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 105.134 0.000 105.454 0.600 ;
  LAYER ME3 ;
  RECT 105.134 0.000 105.454 0.600 ;
  LAYER ME2 ;
  RECT 105.134 0.000 105.454 0.600 ;
  LAYER ME1 ;
  RECT 105.134 0.000 105.454 0.600 ;
 END
 ANTENNAPARTIALMETALAREA                  1.058 LAYER ME2 ;
 ANTENNAGATEAREA                          0.072 LAYER ME2 ;
 ANTENNAGATEAREA                          0.072 LAYER ME3 ;
 ANTENNAGATEAREA                          0.072 LAYER ME4 ;
 ANTENNADIFFAREA                          0.160 LAYER ME2 ;
 ANTENNADIFFAREA                          0.160 LAYER ME3 ;
 ANTENNADIFFAREA                          0.160 LAYER ME4 ;
 ANTENNAMAXAREACAR                       21.782 LAYER ME2 ;
 ANTENNAMAXAREACAR                       24.449 LAYER ME3 ;
 ANTENNAMAXAREACAR                       27.116 LAYER ME4 ;
END DI25
PIN DO25
  DIRECTION OUTPUT ;
 PORT
  LAYER ME4 ;
  RECT 104.572 0.000 104.892 0.600 ;
  LAYER ME3 ;
  RECT 104.572 0.000 104.892 0.600 ;
  LAYER ME2 ;
  RECT 104.572 0.000 104.892 0.600 ;
  LAYER ME1 ;
  RECT 104.572 0.000 104.892 0.600 ;
 END
 ANTENNAPARTIALMETALAREA                  5.273 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME3 ;
 ANTENNADIFFAREA                          1.293 LAYER ME4 ;
END DO25
PIN DI24
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 100.568 0.000 100.888 0.600 ;
  LAYER ME3 ;
  RECT 100.568 0.000 100.888 0.600 ;
  LAYER ME2 ;
  RECT 100.568 0.000 100.888 0.600 ;
  LAYER ME1 ;
  RECT 100.568 0.000 100.888 0.600 ;
 END
 ANTENNAPARTIALMETALAREA                  0.346 LAYER ME1 ;
 ANTENNAPARTIALMETALAREA                  1.466 LAYER ME2 ;
 ANTENNAPARTIALMETALAREA                  0.508 LAYER ME3 ;
 ANTENNAGATEAREA                          0.072 LAYER ME3 ;
 ANTENNAGATEAREA                          0.072 LAYER ME4 ;
 ANTENNADIFFAREA                          0.218 LAYER ME1 ;
 ANTENNADIFFAREA                          0.218 LAYER ME2 ;
 ANTENNADIFFAREA                          0.218 LAYER ME3 ;
 ANTENNADIFFAREA                          0.218 LAYER ME4 ;
 ANTENNAMAXAREACAR                       17.267 LAYER ME3 ;
 ANTENNAMAXAREACAR                       19.933 LAYER ME4 ;
END DI24
PIN DO24
  DIRECTION OUTPUT ;
 PORT
  LAYER ME4 ;
  RECT 101.130 0.000 101.450 0.600 ;
  LAYER ME3 ;
  RECT 101.130 0.000 101.450 0.600 ;
  LAYER ME2 ;
  RECT 101.130 0.000 101.450 0.600 ;
  LAYER ME1 ;
  RECT 101.130 0.000 101.450 0.600 ;
 END
 ANTENNAPARTIALMETALAREA                  5.602 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME3 ;
 ANTENNADIFFAREA                          1.293 LAYER ME4 ;
END DO24
PIN WEB3
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 99.128 0.000 99.448 0.600 ;
  LAYER ME3 ;
  RECT 99.128 0.000 99.448 0.600 ;
  LAYER ME2 ;
  RECT 99.128 0.000 99.448 0.600 ;
  LAYER ME1 ;
  RECT 99.128 0.000 99.448 0.600 ;
 END
 ANTENNAPARTIALMETALAREA                  1.036 LAYER ME2 ;
 ANTENNAGATEAREA                          0.288 LAYER ME2 ;
 ANTENNAGATEAREA                          0.288 LAYER ME3 ;
 ANTENNAGATEAREA                          0.288 LAYER ME4 ;
 ANTENNADIFFAREA                          0.206 LAYER ME2 ;
 ANTENNADIFFAREA                          0.206 LAYER ME3 ;
 ANTENNADIFFAREA                          0.206 LAYER ME4 ;
 ANTENNAMAXAREACAR                        5.844 LAYER ME2 ;
 ANTENNAMAXAREACAR                        6.511 LAYER ME3 ;
 ANTENNAMAXAREACAR                        7.178 LAYER ME4 ;
END WEB3
PIN DI23
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 97.126 0.000 97.446 0.600 ;
  LAYER ME3 ;
  RECT 97.126 0.000 97.446 0.600 ;
  LAYER ME2 ;
  RECT 97.126 0.000 97.446 0.600 ;
  LAYER ME1 ;
  RECT 97.126 0.000 97.446 0.600 ;
 END
 ANTENNAPARTIALMETALAREA                  1.058 LAYER ME2 ;
 ANTENNAGATEAREA                          0.072 LAYER ME2 ;
 ANTENNAGATEAREA                          0.072 LAYER ME3 ;
 ANTENNAGATEAREA                          0.072 LAYER ME4 ;
 ANTENNADIFFAREA                          0.160 LAYER ME2 ;
 ANTENNADIFFAREA                          0.160 LAYER ME3 ;
 ANTENNADIFFAREA                          0.160 LAYER ME4 ;
 ANTENNAMAXAREACAR                       21.782 LAYER ME2 ;
 ANTENNAMAXAREACAR                       24.449 LAYER ME3 ;
 ANTENNAMAXAREACAR                       27.116 LAYER ME4 ;
END DI23
PIN DO23
  DIRECTION OUTPUT ;
 PORT
  LAYER ME4 ;
  RECT 96.564 0.000 96.884 0.600 ;
  LAYER ME3 ;
  RECT 96.564 0.000 96.884 0.600 ;
  LAYER ME2 ;
  RECT 96.564 0.000 96.884 0.600 ;
  LAYER ME1 ;
  RECT 96.564 0.000 96.884 0.600 ;
 END
 ANTENNAPARTIALMETALAREA                  5.273 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME3 ;
 ANTENNADIFFAREA                          1.293 LAYER ME4 ;
END DO23
PIN DI22
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 93.122 0.000 93.442 0.600 ;
  LAYER ME3 ;
  RECT 93.122 0.000 93.442 0.600 ;
  LAYER ME2 ;
  RECT 93.122 0.000 93.442 0.600 ;
  LAYER ME1 ;
  RECT 93.122 0.000 93.442 0.600 ;
 END
 ANTENNAPARTIALMETALAREA                  1.058 LAYER ME2 ;
 ANTENNAGATEAREA                          0.072 LAYER ME2 ;
 ANTENNAGATEAREA                          0.072 LAYER ME3 ;
 ANTENNAGATEAREA                          0.072 LAYER ME4 ;
 ANTENNADIFFAREA                          0.160 LAYER ME2 ;
 ANTENNADIFFAREA                          0.160 LAYER ME3 ;
 ANTENNADIFFAREA                          0.160 LAYER ME4 ;
 ANTENNAMAXAREACAR                       21.782 LAYER ME2 ;
 ANTENNAMAXAREACAR                       24.449 LAYER ME3 ;
 ANTENNAMAXAREACAR                       27.116 LAYER ME4 ;
END DI22
PIN DO22
  DIRECTION OUTPUT ;
 PORT
  LAYER ME4 ;
  RECT 92.560 0.000 92.880 0.600 ;
  LAYER ME3 ;
  RECT 92.560 0.000 92.880 0.600 ;
  LAYER ME2 ;
  RECT 92.560 0.000 92.880 0.600 ;
  LAYER ME1 ;
  RECT 92.560 0.000 92.880 0.600 ;
 END
 ANTENNAPARTIALMETALAREA                  5.273 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME3 ;
 ANTENNADIFFAREA                          1.293 LAYER ME4 ;
END DO22
PIN DI21
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 89.118 0.000 89.438 0.600 ;
  LAYER ME3 ;
  RECT 89.118 0.000 89.438 0.600 ;
  LAYER ME2 ;
  RECT 89.118 0.000 89.438 0.600 ;
  LAYER ME1 ;
  RECT 89.118 0.000 89.438 0.600 ;
 END
 ANTENNAPARTIALMETALAREA                  1.058 LAYER ME2 ;
 ANTENNAGATEAREA                          0.072 LAYER ME2 ;
 ANTENNAGATEAREA                          0.072 LAYER ME3 ;
 ANTENNAGATEAREA                          0.072 LAYER ME4 ;
 ANTENNADIFFAREA                          0.160 LAYER ME2 ;
 ANTENNADIFFAREA                          0.160 LAYER ME3 ;
 ANTENNADIFFAREA                          0.160 LAYER ME4 ;
 ANTENNAMAXAREACAR                       21.782 LAYER ME2 ;
 ANTENNAMAXAREACAR                       24.449 LAYER ME3 ;
 ANTENNAMAXAREACAR                       27.116 LAYER ME4 ;
END DI21
PIN DO21
  DIRECTION OUTPUT ;
 PORT
  LAYER ME4 ;
  RECT 88.556 0.000 88.876 0.600 ;
  LAYER ME3 ;
  RECT 88.556 0.000 88.876 0.600 ;
  LAYER ME2 ;
  RECT 88.556 0.000 88.876 0.600 ;
  LAYER ME1 ;
  RECT 88.556 0.000 88.876 0.600 ;
 END
 ANTENNAPARTIALMETALAREA                  5.273 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME3 ;
 ANTENNADIFFAREA                          1.293 LAYER ME4 ;
END DO21
PIN DI20
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 85.114 0.000 85.434 0.600 ;
  LAYER ME3 ;
  RECT 85.114 0.000 85.434 0.600 ;
  LAYER ME2 ;
  RECT 85.114 0.000 85.434 0.600 ;
  LAYER ME1 ;
  RECT 85.114 0.000 85.434 0.600 ;
 END
 ANTENNAPARTIALMETALAREA                  1.058 LAYER ME2 ;
 ANTENNAGATEAREA                          0.072 LAYER ME2 ;
 ANTENNAGATEAREA                          0.072 LAYER ME3 ;
 ANTENNAGATEAREA                          0.072 LAYER ME4 ;
 ANTENNADIFFAREA                          0.160 LAYER ME2 ;
 ANTENNADIFFAREA                          0.160 LAYER ME3 ;
 ANTENNADIFFAREA                          0.160 LAYER ME4 ;
 ANTENNAMAXAREACAR                       21.782 LAYER ME2 ;
 ANTENNAMAXAREACAR                       24.449 LAYER ME3 ;
 ANTENNAMAXAREACAR                       27.116 LAYER ME4 ;
END DI20
PIN DO20
  DIRECTION OUTPUT ;
 PORT
  LAYER ME4 ;
  RECT 84.552 0.000 84.872 0.600 ;
  LAYER ME3 ;
  RECT 84.552 0.000 84.872 0.600 ;
  LAYER ME2 ;
  RECT 84.552 0.000 84.872 0.600 ;
  LAYER ME1 ;
  RECT 84.552 0.000 84.872 0.600 ;
 END
 ANTENNAPARTIALMETALAREA                  5.273 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME3 ;
 ANTENNADIFFAREA                          1.293 LAYER ME4 ;
END DO20
PIN DI19
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 81.110 0.000 81.430 0.600 ;
  LAYER ME3 ;
  RECT 81.110 0.000 81.430 0.600 ;
  LAYER ME2 ;
  RECT 81.110 0.000 81.430 0.600 ;
  LAYER ME1 ;
  RECT 81.110 0.000 81.430 0.600 ;
 END
 ANTENNAPARTIALMETALAREA                  1.058 LAYER ME2 ;
 ANTENNAGATEAREA                          0.072 LAYER ME2 ;
 ANTENNAGATEAREA                          0.072 LAYER ME3 ;
 ANTENNAGATEAREA                          0.072 LAYER ME4 ;
 ANTENNADIFFAREA                          0.160 LAYER ME2 ;
 ANTENNADIFFAREA                          0.160 LAYER ME3 ;
 ANTENNADIFFAREA                          0.160 LAYER ME4 ;
 ANTENNAMAXAREACAR                       21.782 LAYER ME2 ;
 ANTENNAMAXAREACAR                       24.449 LAYER ME3 ;
 ANTENNAMAXAREACAR                       27.116 LAYER ME4 ;
END DI19
PIN DO19
  DIRECTION OUTPUT ;
 PORT
  LAYER ME4 ;
  RECT 80.548 0.000 80.868 0.600 ;
  LAYER ME3 ;
  RECT 80.548 0.000 80.868 0.600 ;
  LAYER ME2 ;
  RECT 80.548 0.000 80.868 0.600 ;
  LAYER ME1 ;
  RECT 80.548 0.000 80.868 0.600 ;
 END
 ANTENNAPARTIALMETALAREA                  5.273 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME3 ;
 ANTENNADIFFAREA                          1.293 LAYER ME4 ;
END DO19
PIN DI18
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 77.106 0.000 77.426 0.600 ;
  LAYER ME3 ;
  RECT 77.106 0.000 77.426 0.600 ;
  LAYER ME2 ;
  RECT 77.106 0.000 77.426 0.600 ;
  LAYER ME1 ;
  RECT 77.106 0.000 77.426 0.600 ;
 END
 ANTENNAPARTIALMETALAREA                  1.058 LAYER ME2 ;
 ANTENNAGATEAREA                          0.072 LAYER ME2 ;
 ANTENNAGATEAREA                          0.072 LAYER ME3 ;
 ANTENNAGATEAREA                          0.072 LAYER ME4 ;
 ANTENNADIFFAREA                          0.160 LAYER ME2 ;
 ANTENNADIFFAREA                          0.160 LAYER ME3 ;
 ANTENNADIFFAREA                          0.160 LAYER ME4 ;
 ANTENNAMAXAREACAR                       21.782 LAYER ME2 ;
 ANTENNAMAXAREACAR                       24.449 LAYER ME3 ;
 ANTENNAMAXAREACAR                       27.116 LAYER ME4 ;
END DI18
PIN DO18
  DIRECTION OUTPUT ;
 PORT
  LAYER ME4 ;
  RECT 76.544 0.000 76.864 0.600 ;
  LAYER ME3 ;
  RECT 76.544 0.000 76.864 0.600 ;
  LAYER ME2 ;
  RECT 76.544 0.000 76.864 0.600 ;
  LAYER ME1 ;
  RECT 76.544 0.000 76.864 0.600 ;
 END
 ANTENNAPARTIALMETALAREA                  5.273 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME3 ;
 ANTENNADIFFAREA                          1.293 LAYER ME4 ;
END DO18
PIN DI17
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 73.102 0.000 73.422 0.600 ;
  LAYER ME3 ;
  RECT 73.102 0.000 73.422 0.600 ;
  LAYER ME2 ;
  RECT 73.102 0.000 73.422 0.600 ;
  LAYER ME1 ;
  RECT 73.102 0.000 73.422 0.600 ;
 END
 ANTENNAPARTIALMETALAREA                  1.058 LAYER ME2 ;
 ANTENNAGATEAREA                          0.072 LAYER ME2 ;
 ANTENNAGATEAREA                          0.072 LAYER ME3 ;
 ANTENNAGATEAREA                          0.072 LAYER ME4 ;
 ANTENNADIFFAREA                          0.160 LAYER ME2 ;
 ANTENNADIFFAREA                          0.160 LAYER ME3 ;
 ANTENNADIFFAREA                          0.160 LAYER ME4 ;
 ANTENNAMAXAREACAR                       21.782 LAYER ME2 ;
 ANTENNAMAXAREACAR                       24.449 LAYER ME3 ;
 ANTENNAMAXAREACAR                       27.116 LAYER ME4 ;
END DI17
PIN DO17
  DIRECTION OUTPUT ;
 PORT
  LAYER ME4 ;
  RECT 72.540 0.000 72.860 0.600 ;
  LAYER ME3 ;
  RECT 72.540 0.000 72.860 0.600 ;
  LAYER ME2 ;
  RECT 72.540 0.000 72.860 0.600 ;
  LAYER ME1 ;
  RECT 72.540 0.000 72.860 0.600 ;
 END
 ANTENNAPARTIALMETALAREA                  5.273 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME3 ;
 ANTENNADIFFAREA                          1.293 LAYER ME4 ;
END DO17
PIN DI16
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 68.536 0.000 68.856 0.600 ;
  LAYER ME3 ;
  RECT 68.536 0.000 68.856 0.600 ;
  LAYER ME2 ;
  RECT 68.536 0.000 68.856 0.600 ;
  LAYER ME1 ;
  RECT 68.536 0.000 68.856 0.600 ;
 END
 ANTENNAPARTIALMETALAREA                  0.346 LAYER ME1 ;
 ANTENNAPARTIALMETALAREA                  1.466 LAYER ME2 ;
 ANTENNAPARTIALMETALAREA                  0.508 LAYER ME3 ;
 ANTENNAGATEAREA                          0.072 LAYER ME3 ;
 ANTENNAGATEAREA                          0.072 LAYER ME4 ;
 ANTENNADIFFAREA                          0.218 LAYER ME1 ;
 ANTENNADIFFAREA                          0.218 LAYER ME2 ;
 ANTENNADIFFAREA                          0.218 LAYER ME3 ;
 ANTENNADIFFAREA                          0.218 LAYER ME4 ;
 ANTENNAMAXAREACAR                       17.267 LAYER ME3 ;
 ANTENNAMAXAREACAR                       19.933 LAYER ME4 ;
END DI16
PIN DO16
  DIRECTION OUTPUT ;
 PORT
  LAYER ME4 ;
  RECT 69.098 0.000 69.418 0.600 ;
  LAYER ME3 ;
  RECT 69.098 0.000 69.418 0.600 ;
  LAYER ME2 ;
  RECT 69.098 0.000 69.418 0.600 ;
  LAYER ME1 ;
  RECT 69.098 0.000 69.418 0.600 ;
 END
 ANTENNAPARTIALMETALAREA                  5.602 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME3 ;
 ANTENNADIFFAREA                          1.293 LAYER ME4 ;
END DO16
PIN WEB2
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 67.096 0.000 67.416 0.600 ;
  LAYER ME3 ;
  RECT 67.096 0.000 67.416 0.600 ;
  LAYER ME2 ;
  RECT 67.096 0.000 67.416 0.600 ;
  LAYER ME1 ;
  RECT 67.096 0.000 67.416 0.600 ;
 END
 ANTENNAPARTIALMETALAREA                  1.036 LAYER ME2 ;
 ANTENNAGATEAREA                          0.288 LAYER ME2 ;
 ANTENNAGATEAREA                          0.288 LAYER ME3 ;
 ANTENNAGATEAREA                          0.288 LAYER ME4 ;
 ANTENNADIFFAREA                          0.206 LAYER ME2 ;
 ANTENNADIFFAREA                          0.206 LAYER ME3 ;
 ANTENNADIFFAREA                          0.206 LAYER ME4 ;
 ANTENNAMAXAREACAR                        5.844 LAYER ME2 ;
 ANTENNAMAXAREACAR                        6.511 LAYER ME3 ;
 ANTENNAMAXAREACAR                        7.178 LAYER ME4 ;
END WEB2
PIN DI15
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 65.094 0.000 65.414 0.600 ;
  LAYER ME3 ;
  RECT 65.094 0.000 65.414 0.600 ;
  LAYER ME2 ;
  RECT 65.094 0.000 65.414 0.600 ;
  LAYER ME1 ;
  RECT 65.094 0.000 65.414 0.600 ;
 END
 ANTENNAPARTIALMETALAREA                  1.058 LAYER ME2 ;
 ANTENNAGATEAREA                          0.072 LAYER ME2 ;
 ANTENNAGATEAREA                          0.072 LAYER ME3 ;
 ANTENNAGATEAREA                          0.072 LAYER ME4 ;
 ANTENNADIFFAREA                          0.160 LAYER ME2 ;
 ANTENNADIFFAREA                          0.160 LAYER ME3 ;
 ANTENNADIFFAREA                          0.160 LAYER ME4 ;
 ANTENNAMAXAREACAR                       21.782 LAYER ME2 ;
 ANTENNAMAXAREACAR                       24.449 LAYER ME3 ;
 ANTENNAMAXAREACAR                       27.116 LAYER ME4 ;
END DI15
PIN DO15
  DIRECTION OUTPUT ;
 PORT
  LAYER ME4 ;
  RECT 64.532 0.000 64.852 0.600 ;
  LAYER ME3 ;
  RECT 64.532 0.000 64.852 0.600 ;
  LAYER ME2 ;
  RECT 64.532 0.000 64.852 0.600 ;
  LAYER ME1 ;
  RECT 64.532 0.000 64.852 0.600 ;
 END
 ANTENNAPARTIALMETALAREA                  5.273 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME3 ;
 ANTENNADIFFAREA                          1.293 LAYER ME4 ;
END DO15
PIN DI14
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 61.090 0.000 61.410 0.600 ;
  LAYER ME3 ;
  RECT 61.090 0.000 61.410 0.600 ;
  LAYER ME2 ;
  RECT 61.090 0.000 61.410 0.600 ;
  LAYER ME1 ;
  RECT 61.090 0.000 61.410 0.600 ;
 END
 ANTENNAPARTIALMETALAREA                  1.058 LAYER ME2 ;
 ANTENNAGATEAREA                          0.072 LAYER ME2 ;
 ANTENNAGATEAREA                          0.072 LAYER ME3 ;
 ANTENNAGATEAREA                          0.072 LAYER ME4 ;
 ANTENNADIFFAREA                          0.160 LAYER ME2 ;
 ANTENNADIFFAREA                          0.160 LAYER ME3 ;
 ANTENNADIFFAREA                          0.160 LAYER ME4 ;
 ANTENNAMAXAREACAR                       21.782 LAYER ME2 ;
 ANTENNAMAXAREACAR                       24.449 LAYER ME3 ;
 ANTENNAMAXAREACAR                       27.116 LAYER ME4 ;
END DI14
PIN DO14
  DIRECTION OUTPUT ;
 PORT
  LAYER ME4 ;
  RECT 60.528 0.000 60.848 0.600 ;
  LAYER ME3 ;
  RECT 60.528 0.000 60.848 0.600 ;
  LAYER ME2 ;
  RECT 60.528 0.000 60.848 0.600 ;
  LAYER ME1 ;
  RECT 60.528 0.000 60.848 0.600 ;
 END
 ANTENNAPARTIALMETALAREA                  5.273 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME3 ;
 ANTENNADIFFAREA                          1.293 LAYER ME4 ;
END DO14
PIN DI13
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 57.086 0.000 57.406 0.600 ;
  LAYER ME3 ;
  RECT 57.086 0.000 57.406 0.600 ;
  LAYER ME2 ;
  RECT 57.086 0.000 57.406 0.600 ;
  LAYER ME1 ;
  RECT 57.086 0.000 57.406 0.600 ;
 END
 ANTENNAPARTIALMETALAREA                  1.058 LAYER ME2 ;
 ANTENNAGATEAREA                          0.072 LAYER ME2 ;
 ANTENNAGATEAREA                          0.072 LAYER ME3 ;
 ANTENNAGATEAREA                          0.072 LAYER ME4 ;
 ANTENNADIFFAREA                          0.160 LAYER ME2 ;
 ANTENNADIFFAREA                          0.160 LAYER ME3 ;
 ANTENNADIFFAREA                          0.160 LAYER ME4 ;
 ANTENNAMAXAREACAR                       21.782 LAYER ME2 ;
 ANTENNAMAXAREACAR                       24.449 LAYER ME3 ;
 ANTENNAMAXAREACAR                       27.116 LAYER ME4 ;
END DI13
PIN DO13
  DIRECTION OUTPUT ;
 PORT
  LAYER ME4 ;
  RECT 56.524 0.000 56.844 0.600 ;
  LAYER ME3 ;
  RECT 56.524 0.000 56.844 0.600 ;
  LAYER ME2 ;
  RECT 56.524 0.000 56.844 0.600 ;
  LAYER ME1 ;
  RECT 56.524 0.000 56.844 0.600 ;
 END
 ANTENNAPARTIALMETALAREA                  5.273 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME3 ;
 ANTENNADIFFAREA                          1.293 LAYER ME4 ;
END DO13
PIN DI12
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 53.082 0.000 53.402 0.600 ;
  LAYER ME3 ;
  RECT 53.082 0.000 53.402 0.600 ;
  LAYER ME2 ;
  RECT 53.082 0.000 53.402 0.600 ;
  LAYER ME1 ;
  RECT 53.082 0.000 53.402 0.600 ;
 END
 ANTENNAPARTIALMETALAREA                  1.058 LAYER ME2 ;
 ANTENNAGATEAREA                          0.072 LAYER ME2 ;
 ANTENNAGATEAREA                          0.072 LAYER ME3 ;
 ANTENNAGATEAREA                          0.072 LAYER ME4 ;
 ANTENNADIFFAREA                          0.160 LAYER ME2 ;
 ANTENNADIFFAREA                          0.160 LAYER ME3 ;
 ANTENNADIFFAREA                          0.160 LAYER ME4 ;
 ANTENNAMAXAREACAR                       21.782 LAYER ME2 ;
 ANTENNAMAXAREACAR                       24.449 LAYER ME3 ;
 ANTENNAMAXAREACAR                       27.116 LAYER ME4 ;
END DI12
PIN DO12
  DIRECTION OUTPUT ;
 PORT
  LAYER ME4 ;
  RECT 52.520 0.000 52.840 0.600 ;
  LAYER ME3 ;
  RECT 52.520 0.000 52.840 0.600 ;
  LAYER ME2 ;
  RECT 52.520 0.000 52.840 0.600 ;
  LAYER ME1 ;
  RECT 52.520 0.000 52.840 0.600 ;
 END
 ANTENNAPARTIALMETALAREA                  5.273 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME3 ;
 ANTENNADIFFAREA                          1.293 LAYER ME4 ;
END DO12
PIN DI11
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 49.078 0.000 49.398 0.600 ;
  LAYER ME3 ;
  RECT 49.078 0.000 49.398 0.600 ;
  LAYER ME2 ;
  RECT 49.078 0.000 49.398 0.600 ;
  LAYER ME1 ;
  RECT 49.078 0.000 49.398 0.600 ;
 END
 ANTENNAPARTIALMETALAREA                  1.058 LAYER ME2 ;
 ANTENNAGATEAREA                          0.072 LAYER ME2 ;
 ANTENNAGATEAREA                          0.072 LAYER ME3 ;
 ANTENNAGATEAREA                          0.072 LAYER ME4 ;
 ANTENNADIFFAREA                          0.160 LAYER ME2 ;
 ANTENNADIFFAREA                          0.160 LAYER ME3 ;
 ANTENNADIFFAREA                          0.160 LAYER ME4 ;
 ANTENNAMAXAREACAR                       21.782 LAYER ME2 ;
 ANTENNAMAXAREACAR                       24.449 LAYER ME3 ;
 ANTENNAMAXAREACAR                       27.116 LAYER ME4 ;
END DI11
PIN DO11
  DIRECTION OUTPUT ;
 PORT
  LAYER ME4 ;
  RECT 48.516 0.000 48.836 0.600 ;
  LAYER ME3 ;
  RECT 48.516 0.000 48.836 0.600 ;
  LAYER ME2 ;
  RECT 48.516 0.000 48.836 0.600 ;
  LAYER ME1 ;
  RECT 48.516 0.000 48.836 0.600 ;
 END
 ANTENNAPARTIALMETALAREA                  5.273 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME3 ;
 ANTENNADIFFAREA                          1.293 LAYER ME4 ;
END DO11
PIN DI10
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 45.074 0.000 45.394 0.600 ;
  LAYER ME3 ;
  RECT 45.074 0.000 45.394 0.600 ;
  LAYER ME2 ;
  RECT 45.074 0.000 45.394 0.600 ;
  LAYER ME1 ;
  RECT 45.074 0.000 45.394 0.600 ;
 END
 ANTENNAPARTIALMETALAREA                  1.058 LAYER ME2 ;
 ANTENNAGATEAREA                          0.072 LAYER ME2 ;
 ANTENNAGATEAREA                          0.072 LAYER ME3 ;
 ANTENNAGATEAREA                          0.072 LAYER ME4 ;
 ANTENNADIFFAREA                          0.160 LAYER ME2 ;
 ANTENNADIFFAREA                          0.160 LAYER ME3 ;
 ANTENNADIFFAREA                          0.160 LAYER ME4 ;
 ANTENNAMAXAREACAR                       21.782 LAYER ME2 ;
 ANTENNAMAXAREACAR                       24.449 LAYER ME3 ;
 ANTENNAMAXAREACAR                       27.116 LAYER ME4 ;
END DI10
PIN DO10
  DIRECTION OUTPUT ;
 PORT
  LAYER ME4 ;
  RECT 44.512 0.000 44.832 0.600 ;
  LAYER ME3 ;
  RECT 44.512 0.000 44.832 0.600 ;
  LAYER ME2 ;
  RECT 44.512 0.000 44.832 0.600 ;
  LAYER ME1 ;
  RECT 44.512 0.000 44.832 0.600 ;
 END
 ANTENNAPARTIALMETALAREA                  5.273 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME3 ;
 ANTENNADIFFAREA                          1.293 LAYER ME4 ;
END DO10
PIN DI9
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 41.070 0.000 41.390 0.600 ;
  LAYER ME3 ;
  RECT 41.070 0.000 41.390 0.600 ;
  LAYER ME2 ;
  RECT 41.070 0.000 41.390 0.600 ;
  LAYER ME1 ;
  RECT 41.070 0.000 41.390 0.600 ;
 END
 ANTENNAPARTIALMETALAREA                  1.058 LAYER ME2 ;
 ANTENNAGATEAREA                          0.072 LAYER ME2 ;
 ANTENNAGATEAREA                          0.072 LAYER ME3 ;
 ANTENNAGATEAREA                          0.072 LAYER ME4 ;
 ANTENNADIFFAREA                          0.160 LAYER ME2 ;
 ANTENNADIFFAREA                          0.160 LAYER ME3 ;
 ANTENNADIFFAREA                          0.160 LAYER ME4 ;
 ANTENNAMAXAREACAR                       21.782 LAYER ME2 ;
 ANTENNAMAXAREACAR                       24.449 LAYER ME3 ;
 ANTENNAMAXAREACAR                       27.116 LAYER ME4 ;
END DI9
PIN DO9
  DIRECTION OUTPUT ;
 PORT
  LAYER ME4 ;
  RECT 40.508 0.000 40.828 0.600 ;
  LAYER ME3 ;
  RECT 40.508 0.000 40.828 0.600 ;
  LAYER ME2 ;
  RECT 40.508 0.000 40.828 0.600 ;
  LAYER ME1 ;
  RECT 40.508 0.000 40.828 0.600 ;
 END
 ANTENNAPARTIALMETALAREA                  5.273 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME3 ;
 ANTENNADIFFAREA                          1.293 LAYER ME4 ;
END DO9
PIN DI8
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 36.504 0.000 36.824 0.600 ;
  LAYER ME3 ;
  RECT 36.504 0.000 36.824 0.600 ;
  LAYER ME2 ;
  RECT 36.504 0.000 36.824 0.600 ;
  LAYER ME1 ;
  RECT 36.504 0.000 36.824 0.600 ;
 END
 ANTENNAPARTIALMETALAREA                  0.346 LAYER ME1 ;
 ANTENNAPARTIALMETALAREA                  1.466 LAYER ME2 ;
 ANTENNAPARTIALMETALAREA                  0.508 LAYER ME3 ;
 ANTENNAGATEAREA                          0.072 LAYER ME3 ;
 ANTENNAGATEAREA                          0.072 LAYER ME4 ;
 ANTENNADIFFAREA                          0.218 LAYER ME1 ;
 ANTENNADIFFAREA                          0.218 LAYER ME2 ;
 ANTENNADIFFAREA                          0.218 LAYER ME3 ;
 ANTENNADIFFAREA                          0.218 LAYER ME4 ;
 ANTENNAMAXAREACAR                       17.267 LAYER ME3 ;
 ANTENNAMAXAREACAR                       19.933 LAYER ME4 ;
END DI8
PIN DO8
  DIRECTION OUTPUT ;
 PORT
  LAYER ME4 ;
  RECT 37.066 0.000 37.386 0.600 ;
  LAYER ME3 ;
  RECT 37.066 0.000 37.386 0.600 ;
  LAYER ME2 ;
  RECT 37.066 0.000 37.386 0.600 ;
  LAYER ME1 ;
  RECT 37.066 0.000 37.386 0.600 ;
 END
 ANTENNAPARTIALMETALAREA                  5.602 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME3 ;
 ANTENNADIFFAREA                          1.293 LAYER ME4 ;
END DO8
PIN WEB1
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 35.064 0.000 35.384 0.600 ;
  LAYER ME3 ;
  RECT 35.064 0.000 35.384 0.600 ;
  LAYER ME2 ;
  RECT 35.064 0.000 35.384 0.600 ;
  LAYER ME1 ;
  RECT 35.064 0.000 35.384 0.600 ;
 END
 ANTENNAPARTIALMETALAREA                  1.036 LAYER ME2 ;
 ANTENNAGATEAREA                          0.288 LAYER ME2 ;
 ANTENNAGATEAREA                          0.288 LAYER ME3 ;
 ANTENNAGATEAREA                          0.288 LAYER ME4 ;
 ANTENNADIFFAREA                          0.206 LAYER ME2 ;
 ANTENNADIFFAREA                          0.206 LAYER ME3 ;
 ANTENNADIFFAREA                          0.206 LAYER ME4 ;
 ANTENNAMAXAREACAR                        5.844 LAYER ME2 ;
 ANTENNAMAXAREACAR                        6.511 LAYER ME3 ;
 ANTENNAMAXAREACAR                        7.178 LAYER ME4 ;
END WEB1
PIN DI7
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 33.062 0.000 33.382 0.600 ;
  LAYER ME3 ;
  RECT 33.062 0.000 33.382 0.600 ;
  LAYER ME2 ;
  RECT 33.062 0.000 33.382 0.600 ;
  LAYER ME1 ;
  RECT 33.062 0.000 33.382 0.600 ;
 END
 ANTENNAPARTIALMETALAREA                  1.058 LAYER ME2 ;
 ANTENNAGATEAREA                          0.072 LAYER ME2 ;
 ANTENNAGATEAREA                          0.072 LAYER ME3 ;
 ANTENNAGATEAREA                          0.072 LAYER ME4 ;
 ANTENNADIFFAREA                          0.160 LAYER ME2 ;
 ANTENNADIFFAREA                          0.160 LAYER ME3 ;
 ANTENNADIFFAREA                          0.160 LAYER ME4 ;
 ANTENNAMAXAREACAR                       21.782 LAYER ME2 ;
 ANTENNAMAXAREACAR                       24.449 LAYER ME3 ;
 ANTENNAMAXAREACAR                       27.116 LAYER ME4 ;
END DI7
PIN DO7
  DIRECTION OUTPUT ;
 PORT
  LAYER ME4 ;
  RECT 32.500 0.000 32.820 0.600 ;
  LAYER ME3 ;
  RECT 32.500 0.000 32.820 0.600 ;
  LAYER ME2 ;
  RECT 32.500 0.000 32.820 0.600 ;
  LAYER ME1 ;
  RECT 32.500 0.000 32.820 0.600 ;
 END
 ANTENNAPARTIALMETALAREA                  5.273 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME3 ;
 ANTENNADIFFAREA                          1.293 LAYER ME4 ;
END DO7
PIN DI6
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 29.058 0.000 29.378 0.600 ;
  LAYER ME3 ;
  RECT 29.058 0.000 29.378 0.600 ;
  LAYER ME2 ;
  RECT 29.058 0.000 29.378 0.600 ;
  LAYER ME1 ;
  RECT 29.058 0.000 29.378 0.600 ;
 END
 ANTENNAPARTIALMETALAREA                  1.058 LAYER ME2 ;
 ANTENNAGATEAREA                          0.072 LAYER ME2 ;
 ANTENNAGATEAREA                          0.072 LAYER ME3 ;
 ANTENNAGATEAREA                          0.072 LAYER ME4 ;
 ANTENNADIFFAREA                          0.160 LAYER ME2 ;
 ANTENNADIFFAREA                          0.160 LAYER ME3 ;
 ANTENNADIFFAREA                          0.160 LAYER ME4 ;
 ANTENNAMAXAREACAR                       21.782 LAYER ME2 ;
 ANTENNAMAXAREACAR                       24.449 LAYER ME3 ;
 ANTENNAMAXAREACAR                       27.116 LAYER ME4 ;
END DI6
PIN DO6
  DIRECTION OUTPUT ;
 PORT
  LAYER ME4 ;
  RECT 28.496 0.000 28.816 0.600 ;
  LAYER ME3 ;
  RECT 28.496 0.000 28.816 0.600 ;
  LAYER ME2 ;
  RECT 28.496 0.000 28.816 0.600 ;
  LAYER ME1 ;
  RECT 28.496 0.000 28.816 0.600 ;
 END
 ANTENNAPARTIALMETALAREA                  5.273 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME3 ;
 ANTENNADIFFAREA                          1.293 LAYER ME4 ;
END DO6
PIN DI5
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 25.054 0.000 25.374 0.600 ;
  LAYER ME3 ;
  RECT 25.054 0.000 25.374 0.600 ;
  LAYER ME2 ;
  RECT 25.054 0.000 25.374 0.600 ;
  LAYER ME1 ;
  RECT 25.054 0.000 25.374 0.600 ;
 END
 ANTENNAPARTIALMETALAREA                  1.058 LAYER ME2 ;
 ANTENNAGATEAREA                          0.072 LAYER ME2 ;
 ANTENNAGATEAREA                          0.072 LAYER ME3 ;
 ANTENNAGATEAREA                          0.072 LAYER ME4 ;
 ANTENNADIFFAREA                          0.160 LAYER ME2 ;
 ANTENNADIFFAREA                          0.160 LAYER ME3 ;
 ANTENNADIFFAREA                          0.160 LAYER ME4 ;
 ANTENNAMAXAREACAR                       21.782 LAYER ME2 ;
 ANTENNAMAXAREACAR                       24.449 LAYER ME3 ;
 ANTENNAMAXAREACAR                       27.116 LAYER ME4 ;
END DI5
PIN DO5
  DIRECTION OUTPUT ;
 PORT
  LAYER ME4 ;
  RECT 24.492 0.000 24.812 0.600 ;
  LAYER ME3 ;
  RECT 24.492 0.000 24.812 0.600 ;
  LAYER ME2 ;
  RECT 24.492 0.000 24.812 0.600 ;
  LAYER ME1 ;
  RECT 24.492 0.000 24.812 0.600 ;
 END
 ANTENNAPARTIALMETALAREA                  5.273 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME3 ;
 ANTENNADIFFAREA                          1.293 LAYER ME4 ;
END DO5
PIN DI4
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 21.050 0.000 21.370 0.600 ;
  LAYER ME3 ;
  RECT 21.050 0.000 21.370 0.600 ;
  LAYER ME2 ;
  RECT 21.050 0.000 21.370 0.600 ;
  LAYER ME1 ;
  RECT 21.050 0.000 21.370 0.600 ;
 END
 ANTENNAPARTIALMETALAREA                  1.058 LAYER ME2 ;
 ANTENNAGATEAREA                          0.072 LAYER ME2 ;
 ANTENNAGATEAREA                          0.072 LAYER ME3 ;
 ANTENNAGATEAREA                          0.072 LAYER ME4 ;
 ANTENNADIFFAREA                          0.160 LAYER ME2 ;
 ANTENNADIFFAREA                          0.160 LAYER ME3 ;
 ANTENNADIFFAREA                          0.160 LAYER ME4 ;
 ANTENNAMAXAREACAR                       21.782 LAYER ME2 ;
 ANTENNAMAXAREACAR                       24.449 LAYER ME3 ;
 ANTENNAMAXAREACAR                       27.116 LAYER ME4 ;
END DI4
PIN DO4
  DIRECTION OUTPUT ;
 PORT
  LAYER ME4 ;
  RECT 20.488 0.000 20.808 0.600 ;
  LAYER ME3 ;
  RECT 20.488 0.000 20.808 0.600 ;
  LAYER ME2 ;
  RECT 20.488 0.000 20.808 0.600 ;
  LAYER ME1 ;
  RECT 20.488 0.000 20.808 0.600 ;
 END
 ANTENNAPARTIALMETALAREA                  5.273 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME3 ;
 ANTENNADIFFAREA                          1.293 LAYER ME4 ;
END DO4
PIN DI3
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 17.046 0.000 17.366 0.600 ;
  LAYER ME3 ;
  RECT 17.046 0.000 17.366 0.600 ;
  LAYER ME2 ;
  RECT 17.046 0.000 17.366 0.600 ;
  LAYER ME1 ;
  RECT 17.046 0.000 17.366 0.600 ;
 END
 ANTENNAPARTIALMETALAREA                  1.058 LAYER ME2 ;
 ANTENNAGATEAREA                          0.072 LAYER ME2 ;
 ANTENNAGATEAREA                          0.072 LAYER ME3 ;
 ANTENNAGATEAREA                          0.072 LAYER ME4 ;
 ANTENNADIFFAREA                          0.160 LAYER ME2 ;
 ANTENNADIFFAREA                          0.160 LAYER ME3 ;
 ANTENNADIFFAREA                          0.160 LAYER ME4 ;
 ANTENNAMAXAREACAR                       21.782 LAYER ME2 ;
 ANTENNAMAXAREACAR                       24.449 LAYER ME3 ;
 ANTENNAMAXAREACAR                       27.116 LAYER ME4 ;
END DI3
PIN DO3
  DIRECTION OUTPUT ;
 PORT
  LAYER ME4 ;
  RECT 16.484 0.000 16.804 0.600 ;
  LAYER ME3 ;
  RECT 16.484 0.000 16.804 0.600 ;
  LAYER ME2 ;
  RECT 16.484 0.000 16.804 0.600 ;
  LAYER ME1 ;
  RECT 16.484 0.000 16.804 0.600 ;
 END
 ANTENNAPARTIALMETALAREA                  5.273 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME3 ;
 ANTENNADIFFAREA                          1.293 LAYER ME4 ;
END DO3
PIN DI2
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 13.042 0.000 13.362 0.600 ;
  LAYER ME3 ;
  RECT 13.042 0.000 13.362 0.600 ;
  LAYER ME2 ;
  RECT 13.042 0.000 13.362 0.600 ;
  LAYER ME1 ;
  RECT 13.042 0.000 13.362 0.600 ;
 END
 ANTENNAPARTIALMETALAREA                  1.058 LAYER ME2 ;
 ANTENNAGATEAREA                          0.072 LAYER ME2 ;
 ANTENNAGATEAREA                          0.072 LAYER ME3 ;
 ANTENNAGATEAREA                          0.072 LAYER ME4 ;
 ANTENNADIFFAREA                          0.160 LAYER ME2 ;
 ANTENNADIFFAREA                          0.160 LAYER ME3 ;
 ANTENNADIFFAREA                          0.160 LAYER ME4 ;
 ANTENNAMAXAREACAR                       21.782 LAYER ME2 ;
 ANTENNAMAXAREACAR                       24.449 LAYER ME3 ;
 ANTENNAMAXAREACAR                       27.116 LAYER ME4 ;
END DI2
PIN DO2
  DIRECTION OUTPUT ;
 PORT
  LAYER ME4 ;
  RECT 12.480 0.000 12.800 0.600 ;
  LAYER ME3 ;
  RECT 12.480 0.000 12.800 0.600 ;
  LAYER ME2 ;
  RECT 12.480 0.000 12.800 0.600 ;
  LAYER ME1 ;
  RECT 12.480 0.000 12.800 0.600 ;
 END
 ANTENNAPARTIALMETALAREA                  5.273 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME3 ;
 ANTENNADIFFAREA                          1.293 LAYER ME4 ;
END DO2
PIN DI1
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 9.038 0.000 9.358 0.600 ;
  LAYER ME3 ;
  RECT 9.038 0.000 9.358 0.600 ;
  LAYER ME2 ;
  RECT 9.038 0.000 9.358 0.600 ;
  LAYER ME1 ;
  RECT 9.038 0.000 9.358 0.600 ;
 END
 ANTENNAPARTIALMETALAREA                  1.058 LAYER ME2 ;
 ANTENNAGATEAREA                          0.072 LAYER ME2 ;
 ANTENNAGATEAREA                          0.072 LAYER ME3 ;
 ANTENNAGATEAREA                          0.072 LAYER ME4 ;
 ANTENNADIFFAREA                          0.160 LAYER ME2 ;
 ANTENNADIFFAREA                          0.160 LAYER ME3 ;
 ANTENNADIFFAREA                          0.160 LAYER ME4 ;
 ANTENNAMAXAREACAR                       21.782 LAYER ME2 ;
 ANTENNAMAXAREACAR                       24.449 LAYER ME3 ;
 ANTENNAMAXAREACAR                       27.116 LAYER ME4 ;
END DI1
PIN DO1
  DIRECTION OUTPUT ;
 PORT
  LAYER ME4 ;
  RECT 8.476 0.000 8.796 0.600 ;
  LAYER ME3 ;
  RECT 8.476 0.000 8.796 0.600 ;
  LAYER ME2 ;
  RECT 8.476 0.000 8.796 0.600 ;
  LAYER ME1 ;
  RECT 8.476 0.000 8.796 0.600 ;
 END
 ANTENNAPARTIALMETALAREA                  5.273 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME3 ;
 ANTENNADIFFAREA                          1.293 LAYER ME4 ;
END DO1
PIN DI0
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 4.472 0.000 4.792 0.600 ;
  LAYER ME3 ;
  RECT 4.472 0.000 4.792 0.600 ;
  LAYER ME2 ;
  RECT 4.472 0.000 4.792 0.600 ;
  LAYER ME1 ;
  RECT 4.472 0.000 4.792 0.600 ;
 END
 ANTENNAPARTIALMETALAREA                  0.346 LAYER ME1 ;
 ANTENNAPARTIALMETALAREA                  1.466 LAYER ME2 ;
 ANTENNAPARTIALMETALAREA                  0.508 LAYER ME3 ;
 ANTENNAGATEAREA                          0.072 LAYER ME3 ;
 ANTENNAGATEAREA                          0.072 LAYER ME4 ;
 ANTENNADIFFAREA                          0.218 LAYER ME1 ;
 ANTENNADIFFAREA                          0.218 LAYER ME2 ;
 ANTENNADIFFAREA                          0.218 LAYER ME3 ;
 ANTENNADIFFAREA                          0.218 LAYER ME4 ;
 ANTENNAMAXAREACAR                       17.267 LAYER ME3 ;
 ANTENNAMAXAREACAR                       19.933 LAYER ME4 ;
END DI0
PIN DO0
  DIRECTION OUTPUT ;
 PORT
  LAYER ME4 ;
  RECT 5.034 0.000 5.354 0.600 ;
  LAYER ME3 ;
  RECT 5.034 0.000 5.354 0.600 ;
  LAYER ME2 ;
  RECT 5.034 0.000 5.354 0.600 ;
  LAYER ME1 ;
  RECT 5.034 0.000 5.354 0.600 ;
 END
 ANTENNAPARTIALMETALAREA                  5.602 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME3 ;
 ANTENNADIFFAREA                          1.293 LAYER ME4 ;
END DO0
PIN WEB0
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 3.032 0.000 3.352 0.600 ;
  LAYER ME3 ;
  RECT 3.032 0.000 3.352 0.600 ;
  LAYER ME2 ;
  RECT 3.032 0.000 3.352 0.600 ;
  LAYER ME1 ;
  RECT 3.032 0.000 3.352 0.600 ;
 END
 ANTENNAPARTIALMETALAREA                  1.036 LAYER ME2 ;
 ANTENNAGATEAREA                          0.288 LAYER ME2 ;
 ANTENNAGATEAREA                          0.288 LAYER ME3 ;
 ANTENNAGATEAREA                          0.288 LAYER ME4 ;
 ANTENNADIFFAREA                          0.206 LAYER ME2 ;
 ANTENNADIFFAREA                          0.206 LAYER ME3 ;
 ANTENNADIFFAREA                          0.206 LAYER ME4 ;
 ANTENNAMAXAREACAR                        5.844 LAYER ME2 ;
 ANTENNAMAXAREACAR                        6.511 LAYER ME3 ;
 ANTENNAMAXAREACAR                        7.178 LAYER ME4 ;
END WEB0
PIN A1
  DIRECTION INPUT ;
 PORT
  LAYER ME3 ;
  RECT 273.536 0.000 273.856 0.720 ;
  LAYER ME2 ;
  RECT 273.536 0.000 273.856 0.720 ;
  LAYER ME1 ;
  RECT 273.536 0.000 273.856 0.720 ;
 END
 ANTENNAPARTIALMETALAREA                  3.547 LAYER ME2 ;
 ANTENNAGATEAREA                          0.144 LAYER ME2 ;
 ANTENNAGATEAREA                          0.144 LAYER ME3 ;
 ANTENNADIFFAREA                          0.218 LAYER ME2 ;
 ANTENNADIFFAREA                          0.218 LAYER ME3 ;
 ANTENNAMAXAREACAR                       27.235 LAYER ME2 ;
 ANTENNAMAXAREACAR                       28.835 LAYER ME3 ;
END A1
PIN A2
  DIRECTION INPUT ;
 PORT
  LAYER ME3 ;
  RECT 274.106 0.000 274.426 0.720 ;
  LAYER ME2 ;
  RECT 274.106 0.000 274.426 0.720 ;
  LAYER ME1 ;
  RECT 274.106 0.000 274.426 0.720 ;
 END
 ANTENNAPARTIALMETALAREA                  3.688 LAYER ME2 ;
 ANTENNAGATEAREA                          0.144 LAYER ME2 ;
 ANTENNAGATEAREA                          0.144 LAYER ME3 ;
 ANTENNADIFFAREA                          0.218 LAYER ME2 ;
 ANTENNADIFFAREA                          0.218 LAYER ME3 ;
 ANTENNAMAXAREACAR                       28.214 LAYER ME2 ;
 ANTENNAMAXAREACAR                       29.814 LAYER ME3 ;
END A2
PIN A3
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 267.288 0.000 267.608 0.720 ;
  LAYER ME3 ;
  RECT 267.288 0.000 267.608 0.720 ;
  LAYER ME2 ;
  RECT 267.288 0.000 267.608 0.720 ;
  LAYER ME1 ;
  RECT 267.288 0.000 267.608 0.720 ;
 END
 ANTENNAPARTIALMETALAREA                  4.391 LAYER ME2 ;
 ANTENNAGATEAREA                          0.180 LAYER ME2 ;
 ANTENNAGATEAREA                          0.180 LAYER ME3 ;
 ANTENNAGATEAREA                          0.180 LAYER ME4 ;
 ANTENNADIFFAREA                          0.218 LAYER ME2 ;
 ANTENNADIFFAREA                          0.218 LAYER ME3 ;
 ANTENNADIFFAREA                          0.218 LAYER ME4 ;
 ANTENNAMAXAREACAR                       27.451 LAYER ME2 ;
 ANTENNAMAXAREACAR                       28.731 LAYER ME3 ;
 ANTENNAMAXAREACAR                       30.011 LAYER ME4 ;
END A3
PIN A4
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 266.608 0.000 266.928 0.720 ;
  LAYER ME3 ;
  RECT 266.608 0.000 266.928 0.720 ;
  LAYER ME2 ;
  RECT 266.608 0.000 266.928 0.720 ;
  LAYER ME1 ;
  RECT 266.608 0.000 266.928 0.720 ;
 END
 ANTENNAPARTIALMETALAREA                  3.928 LAYER ME2 ;
 ANTENNAGATEAREA                          0.180 LAYER ME2 ;
 ANTENNAGATEAREA                          0.180 LAYER ME3 ;
 ANTENNAGATEAREA                          0.180 LAYER ME4 ;
 ANTENNADIFFAREA                          0.218 LAYER ME2 ;
 ANTENNADIFFAREA                          0.218 LAYER ME3 ;
 ANTENNADIFFAREA                          0.218 LAYER ME4 ;
 ANTENNAMAXAREACAR                       26.813 LAYER ME2 ;
 ANTENNAMAXAREACAR                       28.093 LAYER ME3 ;
 ANTENNAMAXAREACAR                       29.373 LAYER ME4 ;
END A4
PIN A0
  DIRECTION INPUT ;
 PORT
  LAYER ME3 ;
  RECT 284.122 0.000 284.442 0.662 ;
  LAYER ME2 ;
  RECT 284.122 0.000 284.442 0.662 ;
  LAYER ME1 ;
  RECT 284.122 0.000 284.442 0.662 ;
 END
 ANTENNAPARTIALMETALAREA                  5.907 LAYER ME2 ;
 ANTENNAGATEAREA                          0.108 LAYER ME2 ;
 ANTENNAGATEAREA                          0.108 LAYER ME3 ;
 ANTENNADIFFAREA                          0.218 LAYER ME2 ;
 ANTENNADIFFAREA                          0.218 LAYER ME3 ;
 ANTENNAMAXAREACAR                       58.521 LAYER ME2 ;
 ANTENNAMAXAREACAR                       60.482 LAYER ME3 ;
END A0
PIN DVSE
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 293.713 0.000 294.033 0.720 ;
  LAYER ME3 ;
  RECT 293.713 0.000 294.033 0.720 ;
  LAYER ME3 ;
  RECT 293.713 0.000 294.033 0.720 ;
  LAYER ME2 ;
  RECT 293.713 0.000 294.033 0.720 ;
  LAYER ME2 ;
  RECT 293.713 0.000 294.033 0.720 ;
  LAYER ME1 ;
  RECT 293.713 0.000 294.033 0.720 ;
  LAYER ME1 ;
  RECT 293.713 0.000 294.033 0.720 ;
 END
 ANTENNAPARTIALMETALAREA                  7.809 LAYER ME2 ;
 ANTENNAGATEAREA                          0.612 LAYER ME2 ;
 ANTENNAGATEAREA                          0.612 LAYER ME3 ;
 ANTENNAGATEAREA                          0.612 LAYER ME4 ;
 ANTENNADIFFAREA                          0.218 LAYER ME2 ;
 ANTENNADIFFAREA                          0.218 LAYER ME3 ;
 ANTENNADIFFAREA                          0.218 LAYER ME4 ;
 ANTENNAMAXAREACAR                       76.330 LAYER ME2 ;
 ANTENNAMAXAREACAR                       78.463 LAYER ME3 ;
 ANTENNAMAXAREACAR                       80.596 LAYER ME4 ;
END DVSE
PIN DVS3
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 293.193 0.000 293.513 0.720 ;
  LAYER ME3 ;
  RECT 293.193 0.000 293.513 0.720 ;
  LAYER ME3 ;
  RECT 293.193 0.000 293.513 0.720 ;
  LAYER ME2 ;
  RECT 293.193 0.000 293.513 0.720 ;
  LAYER ME2 ;
  RECT 293.193 0.000 293.513 0.720 ;
  LAYER ME1 ;
  RECT 293.193 0.000 293.513 0.720 ;
  LAYER ME1 ;
  RECT 293.193 0.000 293.513 0.720 ;
 END
 ANTENNAPARTIALMETALAREA                  6.179 LAYER ME2 ;
 ANTENNAGATEAREA                          0.108 LAYER ME2 ;
 ANTENNAGATEAREA                          0.108 LAYER ME3 ;
 ANTENNAGATEAREA                          0.108 LAYER ME4 ;
 ANTENNADIFFAREA                          0.218 LAYER ME2 ;
 ANTENNADIFFAREA                          0.218 LAYER ME3 ;
 ANTENNADIFFAREA                          0.218 LAYER ME4 ;
 ANTENNAMAXAREACAR                       68.823 LAYER ME2 ;
 ANTENNAMAXAREACAR                       70.956 LAYER ME3 ;
 ANTENNAMAXAREACAR                       73.089 LAYER ME4 ;
END DVS3
PIN DVS2
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 294.233 0.000 294.553 0.720 ;
  LAYER ME3 ;
  RECT 294.233 0.000 294.553 0.720 ;
  LAYER ME3 ;
  RECT 294.233 0.000 294.553 0.720 ;
  LAYER ME2 ;
  RECT 294.233 0.000 294.553 0.720 ;
  LAYER ME2 ;
  RECT 294.233 0.000 294.553 0.720 ;
  LAYER ME1 ;
  RECT 294.233 0.000 294.553 0.720 ;
  LAYER ME1 ;
  RECT 294.233 0.000 294.553 0.720 ;
 END
 ANTENNAPARTIALMETALAREA                  7.876 LAYER ME2 ;
 ANTENNAGATEAREA                          0.108 LAYER ME2 ;
 ANTENNAGATEAREA                          0.108 LAYER ME3 ;
 ANTENNAGATEAREA                          0.108 LAYER ME4 ;
 ANTENNADIFFAREA                          0.218 LAYER ME2 ;
 ANTENNADIFFAREA                          0.218 LAYER ME3 ;
 ANTENNADIFFAREA                          0.218 LAYER ME4 ;
 ANTENNAMAXAREACAR                       83.257 LAYER ME2 ;
 ANTENNAMAXAREACAR                       85.391 LAYER ME3 ;
 ANTENNAMAXAREACAR                       87.524 LAYER ME4 ;
END DVS2
PIN DVS1
  DIRECTION INPUT ;
 PORT
  LAYER ME3 ;
  RECT 290.577 0.000 290.897 0.720 ;
  LAYER ME2 ;
  RECT 290.577 0.000 290.897 0.720 ;
  LAYER ME1 ;
  RECT 290.577 0.000 290.897 0.720 ;
 END
 ANTENNAPARTIALMETALAREA                  6.247 LAYER ME2 ;
 ANTENNAGATEAREA                          0.108 LAYER ME2 ;
 ANTENNAGATEAREA                          0.108 LAYER ME3 ;
 ANTENNADIFFAREA                          0.218 LAYER ME2 ;
 ANTENNADIFFAREA                          0.218 LAYER ME3 ;
 ANTENNAMAXAREACAR                       69.294 LAYER ME2 ;
 ANTENNAMAXAREACAR                       71.427 LAYER ME3 ;
END DVS1
PIN DVS0
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 294.753 0.000 295.073 0.720 ;
  LAYER ME3 ;
  RECT 294.753 0.000 295.073 0.720 ;
  LAYER ME3 ;
  RECT 294.753 0.000 295.073 0.720 ;
  LAYER ME2 ;
  RECT 294.753 0.000 295.073 0.720 ;
  LAYER ME2 ;
  RECT 294.753 0.000 295.073 0.720 ;
  LAYER ME1 ;
  RECT 294.753 0.000 295.073 0.720 ;
  LAYER ME1 ;
  RECT 294.753 0.000 295.073 0.720 ;
 END
 ANTENNAPARTIALMETALAREA                  7.119 LAYER ME2 ;
 ANTENNAGATEAREA                          0.108 LAYER ME2 ;
 ANTENNAGATEAREA                          0.108 LAYER ME3 ;
 ANTENNAGATEAREA                          0.108 LAYER ME4 ;
 ANTENNADIFFAREA                          0.218 LAYER ME2 ;
 ANTENNADIFFAREA                          0.218 LAYER ME3 ;
 ANTENNADIFFAREA                          0.218 LAYER ME4 ;
 ANTENNAMAXAREACAR                       77.987 LAYER ME2 ;
 ANTENNAMAXAREACAR                       80.120 LAYER ME3 ;
 ANTENNAMAXAREACAR                       82.254 LAYER ME4 ;
END DVS0
PIN CK
  DIRECTION INPUT ;
 PORT
  LAYER ME3 ;
  RECT 286.661 0.000 286.981 0.720 ;
  LAYER ME2 ;
  RECT 286.661 0.000 286.981 0.720 ;
  LAYER ME1 ;
  RECT 286.661 0.000 286.981 0.720 ;
 END
 ANTENNAPARTIALMETALAREA                  5.257 LAYER ME2 ;
 ANTENNAPARTIALMETALAREA                  6.084 LAYER ME3 ;
 ANTENNAGATEAREA                          0.072 LAYER ME2 ;
 ANTENNAGATEAREA                          0.792 LAYER ME3 ;
 ANTENNADIFFAREA                          0.218 LAYER ME2 ;
 ANTENNADIFFAREA                          0.218 LAYER ME3 ;
 ANTENNAMAXAREACAR                       86.308 LAYER ME2 ;
 ANTENNAMAXAREACAR                      174.014 LAYER ME3 ;
END CK
PIN CSB
  DIRECTION INPUT ;
 PORT
  LAYER ME3 ;
  RECT 278.047 0.000 278.367 0.720 ;
  LAYER ME2 ;
  RECT 278.047 0.000 278.367 0.720 ;
  LAYER ME1 ;
  RECT 278.047 0.000 278.367 0.720 ;
 END
 ANTENNAPARTIALMETALAREA                  5.788 LAYER ME2 ;
 ANTENNAPARTIALMETALAREA                  6.164 LAYER ME3 ;
 ANTENNAGATEAREA                          2.508 LAYER ME2 ;
 ANTENNAGATEAREA                          3.228 LAYER ME3 ;
 ANTENNADIFFAREA                          0.218 LAYER ME2 ;
 ANTENNADIFFAREA                          0.218 LAYER ME3 ;
 ANTENNAMAXAREACAR                        3.046 LAYER ME2 ;
 ANTENNAMAXAREACAR                       32.772 LAYER ME3 ;
END CSB
PIN DI127
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 549.619 0.000 549.939 0.600 ;
  LAYER ME3 ;
  RECT 549.619 0.000 549.939 0.600 ;
  LAYER ME2 ;
  RECT 549.619 0.000 549.939 0.600 ;
  LAYER ME1 ;
  RECT 549.619 0.000 549.939 0.600 ;
 END
 ANTENNAPARTIALMETALAREA                  1.058 LAYER ME2 ;
 ANTENNAGATEAREA                          0.072 LAYER ME2 ;
 ANTENNAGATEAREA                          0.072 LAYER ME3 ;
 ANTENNAGATEAREA                          0.072 LAYER ME4 ;
 ANTENNADIFFAREA                          0.160 LAYER ME2 ;
 ANTENNADIFFAREA                          0.160 LAYER ME3 ;
 ANTENNADIFFAREA                          0.160 LAYER ME4 ;
 ANTENNAMAXAREACAR                       21.782 LAYER ME2 ;
 ANTENNAMAXAREACAR                       24.449 LAYER ME3 ;
 ANTENNAMAXAREACAR                       27.116 LAYER ME4 ;
END DI127
PIN DO127
  DIRECTION OUTPUT ;
 PORT
  LAYER ME4 ;
  RECT 549.057 0.000 549.377 0.600 ;
  LAYER ME3 ;
  RECT 549.057 0.000 549.377 0.600 ;
  LAYER ME2 ;
  RECT 549.057 0.000 549.377 0.600 ;
  LAYER ME1 ;
  RECT 549.057 0.000 549.377 0.600 ;
 END
 ANTENNAPARTIALMETALAREA                  5.273 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME3 ;
 ANTENNADIFFAREA                          1.293 LAYER ME4 ;
END DO127
PIN DI126
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 545.615 0.000 545.935 0.600 ;
  LAYER ME3 ;
  RECT 545.615 0.000 545.935 0.600 ;
  LAYER ME2 ;
  RECT 545.615 0.000 545.935 0.600 ;
  LAYER ME1 ;
  RECT 545.615 0.000 545.935 0.600 ;
 END
 ANTENNAPARTIALMETALAREA                  1.058 LAYER ME2 ;
 ANTENNAGATEAREA                          0.072 LAYER ME2 ;
 ANTENNAGATEAREA                          0.072 LAYER ME3 ;
 ANTENNAGATEAREA                          0.072 LAYER ME4 ;
 ANTENNADIFFAREA                          0.160 LAYER ME2 ;
 ANTENNADIFFAREA                          0.160 LAYER ME3 ;
 ANTENNADIFFAREA                          0.160 LAYER ME4 ;
 ANTENNAMAXAREACAR                       21.782 LAYER ME2 ;
 ANTENNAMAXAREACAR                       24.449 LAYER ME3 ;
 ANTENNAMAXAREACAR                       27.116 LAYER ME4 ;
END DI126
PIN DO126
  DIRECTION OUTPUT ;
 PORT
  LAYER ME4 ;
  RECT 545.053 0.000 545.373 0.600 ;
  LAYER ME3 ;
  RECT 545.053 0.000 545.373 0.600 ;
  LAYER ME2 ;
  RECT 545.053 0.000 545.373 0.600 ;
  LAYER ME1 ;
  RECT 545.053 0.000 545.373 0.600 ;
 END
 ANTENNAPARTIALMETALAREA                  5.273 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME3 ;
 ANTENNADIFFAREA                          1.293 LAYER ME4 ;
END DO126
PIN DI125
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 541.611 0.000 541.931 0.600 ;
  LAYER ME3 ;
  RECT 541.611 0.000 541.931 0.600 ;
  LAYER ME2 ;
  RECT 541.611 0.000 541.931 0.600 ;
  LAYER ME1 ;
  RECT 541.611 0.000 541.931 0.600 ;
 END
 ANTENNAPARTIALMETALAREA                  1.058 LAYER ME2 ;
 ANTENNAGATEAREA                          0.072 LAYER ME2 ;
 ANTENNAGATEAREA                          0.072 LAYER ME3 ;
 ANTENNAGATEAREA                          0.072 LAYER ME4 ;
 ANTENNADIFFAREA                          0.160 LAYER ME2 ;
 ANTENNADIFFAREA                          0.160 LAYER ME3 ;
 ANTENNADIFFAREA                          0.160 LAYER ME4 ;
 ANTENNAMAXAREACAR                       21.782 LAYER ME2 ;
 ANTENNAMAXAREACAR                       24.449 LAYER ME3 ;
 ANTENNAMAXAREACAR                       27.116 LAYER ME4 ;
END DI125
PIN DO125
  DIRECTION OUTPUT ;
 PORT
  LAYER ME4 ;
  RECT 541.049 0.000 541.369 0.600 ;
  LAYER ME3 ;
  RECT 541.049 0.000 541.369 0.600 ;
  LAYER ME2 ;
  RECT 541.049 0.000 541.369 0.600 ;
  LAYER ME1 ;
  RECT 541.049 0.000 541.369 0.600 ;
 END
 ANTENNAPARTIALMETALAREA                  5.273 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME3 ;
 ANTENNADIFFAREA                          1.293 LAYER ME4 ;
END DO125
PIN DI124
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 537.607 0.000 537.927 0.600 ;
  LAYER ME3 ;
  RECT 537.607 0.000 537.927 0.600 ;
  LAYER ME2 ;
  RECT 537.607 0.000 537.927 0.600 ;
  LAYER ME1 ;
  RECT 537.607 0.000 537.927 0.600 ;
 END
 ANTENNAPARTIALMETALAREA                  1.058 LAYER ME2 ;
 ANTENNAGATEAREA                          0.072 LAYER ME2 ;
 ANTENNAGATEAREA                          0.072 LAYER ME3 ;
 ANTENNAGATEAREA                          0.072 LAYER ME4 ;
 ANTENNADIFFAREA                          0.160 LAYER ME2 ;
 ANTENNADIFFAREA                          0.160 LAYER ME3 ;
 ANTENNADIFFAREA                          0.160 LAYER ME4 ;
 ANTENNAMAXAREACAR                       21.782 LAYER ME2 ;
 ANTENNAMAXAREACAR                       24.449 LAYER ME3 ;
 ANTENNAMAXAREACAR                       27.116 LAYER ME4 ;
END DI124
PIN DO124
  DIRECTION OUTPUT ;
 PORT
  LAYER ME4 ;
  RECT 537.045 0.000 537.365 0.600 ;
  LAYER ME3 ;
  RECT 537.045 0.000 537.365 0.600 ;
  LAYER ME2 ;
  RECT 537.045 0.000 537.365 0.600 ;
  LAYER ME1 ;
  RECT 537.045 0.000 537.365 0.600 ;
 END
 ANTENNAPARTIALMETALAREA                  5.273 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME3 ;
 ANTENNADIFFAREA                          1.293 LAYER ME4 ;
END DO124
PIN DI123
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 533.603 0.000 533.923 0.600 ;
  LAYER ME3 ;
  RECT 533.603 0.000 533.923 0.600 ;
  LAYER ME2 ;
  RECT 533.603 0.000 533.923 0.600 ;
  LAYER ME1 ;
  RECT 533.603 0.000 533.923 0.600 ;
 END
 ANTENNAPARTIALMETALAREA                  1.058 LAYER ME2 ;
 ANTENNAGATEAREA                          0.072 LAYER ME2 ;
 ANTENNAGATEAREA                          0.072 LAYER ME3 ;
 ANTENNAGATEAREA                          0.072 LAYER ME4 ;
 ANTENNADIFFAREA                          0.160 LAYER ME2 ;
 ANTENNADIFFAREA                          0.160 LAYER ME3 ;
 ANTENNADIFFAREA                          0.160 LAYER ME4 ;
 ANTENNAMAXAREACAR                       21.782 LAYER ME2 ;
 ANTENNAMAXAREACAR                       24.449 LAYER ME3 ;
 ANTENNAMAXAREACAR                       27.116 LAYER ME4 ;
END DI123
PIN DO123
  DIRECTION OUTPUT ;
 PORT
  LAYER ME4 ;
  RECT 533.041 0.000 533.361 0.600 ;
  LAYER ME3 ;
  RECT 533.041 0.000 533.361 0.600 ;
  LAYER ME2 ;
  RECT 533.041 0.000 533.361 0.600 ;
  LAYER ME1 ;
  RECT 533.041 0.000 533.361 0.600 ;
 END
 ANTENNAPARTIALMETALAREA                  5.273 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME3 ;
 ANTENNADIFFAREA                          1.293 LAYER ME4 ;
END DO123
PIN DI122
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 529.599 0.000 529.919 0.600 ;
  LAYER ME3 ;
  RECT 529.599 0.000 529.919 0.600 ;
  LAYER ME2 ;
  RECT 529.599 0.000 529.919 0.600 ;
  LAYER ME1 ;
  RECT 529.599 0.000 529.919 0.600 ;
 END
 ANTENNAPARTIALMETALAREA                  1.058 LAYER ME2 ;
 ANTENNAGATEAREA                          0.072 LAYER ME2 ;
 ANTENNAGATEAREA                          0.072 LAYER ME3 ;
 ANTENNAGATEAREA                          0.072 LAYER ME4 ;
 ANTENNADIFFAREA                          0.160 LAYER ME2 ;
 ANTENNADIFFAREA                          0.160 LAYER ME3 ;
 ANTENNADIFFAREA                          0.160 LAYER ME4 ;
 ANTENNAMAXAREACAR                       21.782 LAYER ME2 ;
 ANTENNAMAXAREACAR                       24.449 LAYER ME3 ;
 ANTENNAMAXAREACAR                       27.116 LAYER ME4 ;
END DI122
PIN DO122
  DIRECTION OUTPUT ;
 PORT
  LAYER ME4 ;
  RECT 529.037 0.000 529.357 0.600 ;
  LAYER ME3 ;
  RECT 529.037 0.000 529.357 0.600 ;
  LAYER ME2 ;
  RECT 529.037 0.000 529.357 0.600 ;
  LAYER ME1 ;
  RECT 529.037 0.000 529.357 0.600 ;
 END
 ANTENNAPARTIALMETALAREA                  5.273 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME3 ;
 ANTENNADIFFAREA                          1.293 LAYER ME4 ;
END DO122
PIN DI121
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 525.595 0.000 525.915 0.600 ;
  LAYER ME3 ;
  RECT 525.595 0.000 525.915 0.600 ;
  LAYER ME2 ;
  RECT 525.595 0.000 525.915 0.600 ;
  LAYER ME1 ;
  RECT 525.595 0.000 525.915 0.600 ;
 END
 ANTENNAPARTIALMETALAREA                  1.058 LAYER ME2 ;
 ANTENNAGATEAREA                          0.072 LAYER ME2 ;
 ANTENNAGATEAREA                          0.072 LAYER ME3 ;
 ANTENNAGATEAREA                          0.072 LAYER ME4 ;
 ANTENNADIFFAREA                          0.160 LAYER ME2 ;
 ANTENNADIFFAREA                          0.160 LAYER ME3 ;
 ANTENNADIFFAREA                          0.160 LAYER ME4 ;
 ANTENNAMAXAREACAR                       21.782 LAYER ME2 ;
 ANTENNAMAXAREACAR                       24.449 LAYER ME3 ;
 ANTENNAMAXAREACAR                       27.116 LAYER ME4 ;
END DI121
PIN DO121
  DIRECTION OUTPUT ;
 PORT
  LAYER ME4 ;
  RECT 525.033 0.000 525.353 0.600 ;
  LAYER ME3 ;
  RECT 525.033 0.000 525.353 0.600 ;
  LAYER ME2 ;
  RECT 525.033 0.000 525.353 0.600 ;
  LAYER ME1 ;
  RECT 525.033 0.000 525.353 0.600 ;
 END
 ANTENNAPARTIALMETALAREA                  5.273 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME3 ;
 ANTENNADIFFAREA                          1.293 LAYER ME4 ;
END DO121
PIN DI120
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 521.029 0.000 521.349 0.600 ;
  LAYER ME3 ;
  RECT 521.029 0.000 521.349 0.600 ;
  LAYER ME2 ;
  RECT 521.029 0.000 521.349 0.600 ;
  LAYER ME1 ;
  RECT 521.029 0.000 521.349 0.600 ;
 END
 ANTENNAPARTIALMETALAREA                  0.346 LAYER ME1 ;
 ANTENNAPARTIALMETALAREA                  1.466 LAYER ME2 ;
 ANTENNAPARTIALMETALAREA                  0.508 LAYER ME3 ;
 ANTENNAGATEAREA                          0.072 LAYER ME3 ;
 ANTENNAGATEAREA                          0.072 LAYER ME4 ;
 ANTENNADIFFAREA                          0.218 LAYER ME1 ;
 ANTENNADIFFAREA                          0.218 LAYER ME2 ;
 ANTENNADIFFAREA                          0.218 LAYER ME3 ;
 ANTENNADIFFAREA                          0.218 LAYER ME4 ;
 ANTENNAMAXAREACAR                       17.267 LAYER ME3 ;
 ANTENNAMAXAREACAR                       19.933 LAYER ME4 ;
END DI120
PIN DO120
  DIRECTION OUTPUT ;
 PORT
  LAYER ME4 ;
  RECT 521.591 0.000 521.911 0.600 ;
  LAYER ME3 ;
  RECT 521.591 0.000 521.911 0.600 ;
  LAYER ME2 ;
  RECT 521.591 0.000 521.911 0.600 ;
  LAYER ME1 ;
  RECT 521.591 0.000 521.911 0.600 ;
 END
 ANTENNAPARTIALMETALAREA                  5.602 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME3 ;
 ANTENNADIFFAREA                          1.293 LAYER ME4 ;
END DO120
PIN WEB15
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 519.589 0.000 519.909 0.600 ;
  LAYER ME3 ;
  RECT 519.589 0.000 519.909 0.600 ;
  LAYER ME2 ;
  RECT 519.589 0.000 519.909 0.600 ;
  LAYER ME1 ;
  RECT 519.589 0.000 519.909 0.600 ;
 END
 ANTENNAPARTIALMETALAREA                  1.036 LAYER ME2 ;
 ANTENNAGATEAREA                          0.288 LAYER ME2 ;
 ANTENNAGATEAREA                          0.288 LAYER ME3 ;
 ANTENNAGATEAREA                          0.288 LAYER ME4 ;
 ANTENNADIFFAREA                          0.206 LAYER ME2 ;
 ANTENNADIFFAREA                          0.206 LAYER ME3 ;
 ANTENNADIFFAREA                          0.206 LAYER ME4 ;
 ANTENNAMAXAREACAR                        5.844 LAYER ME2 ;
 ANTENNAMAXAREACAR                        6.511 LAYER ME3 ;
 ANTENNAMAXAREACAR                        7.178 LAYER ME4 ;
END WEB15
PIN DI119
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 517.587 0.000 517.907 0.600 ;
  LAYER ME3 ;
  RECT 517.587 0.000 517.907 0.600 ;
  LAYER ME2 ;
  RECT 517.587 0.000 517.907 0.600 ;
  LAYER ME1 ;
  RECT 517.587 0.000 517.907 0.600 ;
 END
 ANTENNAPARTIALMETALAREA                  1.058 LAYER ME2 ;
 ANTENNAGATEAREA                          0.072 LAYER ME2 ;
 ANTENNAGATEAREA                          0.072 LAYER ME3 ;
 ANTENNAGATEAREA                          0.072 LAYER ME4 ;
 ANTENNADIFFAREA                          0.160 LAYER ME2 ;
 ANTENNADIFFAREA                          0.160 LAYER ME3 ;
 ANTENNADIFFAREA                          0.160 LAYER ME4 ;
 ANTENNAMAXAREACAR                       21.782 LAYER ME2 ;
 ANTENNAMAXAREACAR                       24.449 LAYER ME3 ;
 ANTENNAMAXAREACAR                       27.116 LAYER ME4 ;
END DI119
PIN DO119
  DIRECTION OUTPUT ;
 PORT
  LAYER ME4 ;
  RECT 517.025 0.000 517.345 0.600 ;
  LAYER ME3 ;
  RECT 517.025 0.000 517.345 0.600 ;
  LAYER ME2 ;
  RECT 517.025 0.000 517.345 0.600 ;
  LAYER ME1 ;
  RECT 517.025 0.000 517.345 0.600 ;
 END
 ANTENNAPARTIALMETALAREA                  5.273 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME3 ;
 ANTENNADIFFAREA                          1.293 LAYER ME4 ;
END DO119
PIN DI118
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 513.583 0.000 513.903 0.600 ;
  LAYER ME3 ;
  RECT 513.583 0.000 513.903 0.600 ;
  LAYER ME2 ;
  RECT 513.583 0.000 513.903 0.600 ;
  LAYER ME1 ;
  RECT 513.583 0.000 513.903 0.600 ;
 END
 ANTENNAPARTIALMETALAREA                  1.058 LAYER ME2 ;
 ANTENNAGATEAREA                          0.072 LAYER ME2 ;
 ANTENNAGATEAREA                          0.072 LAYER ME3 ;
 ANTENNAGATEAREA                          0.072 LAYER ME4 ;
 ANTENNADIFFAREA                          0.160 LAYER ME2 ;
 ANTENNADIFFAREA                          0.160 LAYER ME3 ;
 ANTENNADIFFAREA                          0.160 LAYER ME4 ;
 ANTENNAMAXAREACAR                       21.782 LAYER ME2 ;
 ANTENNAMAXAREACAR                       24.449 LAYER ME3 ;
 ANTENNAMAXAREACAR                       27.116 LAYER ME4 ;
END DI118
PIN DO118
  DIRECTION OUTPUT ;
 PORT
  LAYER ME4 ;
  RECT 513.021 0.000 513.341 0.600 ;
  LAYER ME3 ;
  RECT 513.021 0.000 513.341 0.600 ;
  LAYER ME2 ;
  RECT 513.021 0.000 513.341 0.600 ;
  LAYER ME1 ;
  RECT 513.021 0.000 513.341 0.600 ;
 END
 ANTENNAPARTIALMETALAREA                  5.273 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME3 ;
 ANTENNADIFFAREA                          1.293 LAYER ME4 ;
END DO118
PIN DI117
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 509.579 0.000 509.899 0.600 ;
  LAYER ME3 ;
  RECT 509.579 0.000 509.899 0.600 ;
  LAYER ME2 ;
  RECT 509.579 0.000 509.899 0.600 ;
  LAYER ME1 ;
  RECT 509.579 0.000 509.899 0.600 ;
 END
 ANTENNAPARTIALMETALAREA                  1.058 LAYER ME2 ;
 ANTENNAGATEAREA                          0.072 LAYER ME2 ;
 ANTENNAGATEAREA                          0.072 LAYER ME3 ;
 ANTENNAGATEAREA                          0.072 LAYER ME4 ;
 ANTENNADIFFAREA                          0.160 LAYER ME2 ;
 ANTENNADIFFAREA                          0.160 LAYER ME3 ;
 ANTENNADIFFAREA                          0.160 LAYER ME4 ;
 ANTENNAMAXAREACAR                       21.782 LAYER ME2 ;
 ANTENNAMAXAREACAR                       24.449 LAYER ME3 ;
 ANTENNAMAXAREACAR                       27.116 LAYER ME4 ;
END DI117
PIN DO117
  DIRECTION OUTPUT ;
 PORT
  LAYER ME4 ;
  RECT 509.017 0.000 509.337 0.600 ;
  LAYER ME3 ;
  RECT 509.017 0.000 509.337 0.600 ;
  LAYER ME2 ;
  RECT 509.017 0.000 509.337 0.600 ;
  LAYER ME1 ;
  RECT 509.017 0.000 509.337 0.600 ;
 END
 ANTENNAPARTIALMETALAREA                  5.273 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME3 ;
 ANTENNADIFFAREA                          1.293 LAYER ME4 ;
END DO117
PIN DI116
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 505.575 0.000 505.895 0.600 ;
  LAYER ME3 ;
  RECT 505.575 0.000 505.895 0.600 ;
  LAYER ME2 ;
  RECT 505.575 0.000 505.895 0.600 ;
  LAYER ME1 ;
  RECT 505.575 0.000 505.895 0.600 ;
 END
 ANTENNAPARTIALMETALAREA                  1.058 LAYER ME2 ;
 ANTENNAGATEAREA                          0.072 LAYER ME2 ;
 ANTENNAGATEAREA                          0.072 LAYER ME3 ;
 ANTENNAGATEAREA                          0.072 LAYER ME4 ;
 ANTENNADIFFAREA                          0.160 LAYER ME2 ;
 ANTENNADIFFAREA                          0.160 LAYER ME3 ;
 ANTENNADIFFAREA                          0.160 LAYER ME4 ;
 ANTENNAMAXAREACAR                       21.782 LAYER ME2 ;
 ANTENNAMAXAREACAR                       24.449 LAYER ME3 ;
 ANTENNAMAXAREACAR                       27.116 LAYER ME4 ;
END DI116
PIN DO116
  DIRECTION OUTPUT ;
 PORT
  LAYER ME4 ;
  RECT 505.013 0.000 505.333 0.600 ;
  LAYER ME3 ;
  RECT 505.013 0.000 505.333 0.600 ;
  LAYER ME2 ;
  RECT 505.013 0.000 505.333 0.600 ;
  LAYER ME1 ;
  RECT 505.013 0.000 505.333 0.600 ;
 END
 ANTENNAPARTIALMETALAREA                  5.273 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME3 ;
 ANTENNADIFFAREA                          1.293 LAYER ME4 ;
END DO116
PIN DI115
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 501.571 0.000 501.891 0.600 ;
  LAYER ME3 ;
  RECT 501.571 0.000 501.891 0.600 ;
  LAYER ME2 ;
  RECT 501.571 0.000 501.891 0.600 ;
  LAYER ME1 ;
  RECT 501.571 0.000 501.891 0.600 ;
 END
 ANTENNAPARTIALMETALAREA                  1.058 LAYER ME2 ;
 ANTENNAGATEAREA                          0.072 LAYER ME2 ;
 ANTENNAGATEAREA                          0.072 LAYER ME3 ;
 ANTENNAGATEAREA                          0.072 LAYER ME4 ;
 ANTENNADIFFAREA                          0.160 LAYER ME2 ;
 ANTENNADIFFAREA                          0.160 LAYER ME3 ;
 ANTENNADIFFAREA                          0.160 LAYER ME4 ;
 ANTENNAMAXAREACAR                       21.782 LAYER ME2 ;
 ANTENNAMAXAREACAR                       24.449 LAYER ME3 ;
 ANTENNAMAXAREACAR                       27.116 LAYER ME4 ;
END DI115
PIN DO115
  DIRECTION OUTPUT ;
 PORT
  LAYER ME4 ;
  RECT 501.009 0.000 501.329 0.600 ;
  LAYER ME3 ;
  RECT 501.009 0.000 501.329 0.600 ;
  LAYER ME2 ;
  RECT 501.009 0.000 501.329 0.600 ;
  LAYER ME1 ;
  RECT 501.009 0.000 501.329 0.600 ;
 END
 ANTENNAPARTIALMETALAREA                  5.273 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME3 ;
 ANTENNADIFFAREA                          1.293 LAYER ME4 ;
END DO115
PIN DI114
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 497.567 0.000 497.887 0.600 ;
  LAYER ME3 ;
  RECT 497.567 0.000 497.887 0.600 ;
  LAYER ME2 ;
  RECT 497.567 0.000 497.887 0.600 ;
  LAYER ME1 ;
  RECT 497.567 0.000 497.887 0.600 ;
 END
 ANTENNAPARTIALMETALAREA                  1.058 LAYER ME2 ;
 ANTENNAGATEAREA                          0.072 LAYER ME2 ;
 ANTENNAGATEAREA                          0.072 LAYER ME3 ;
 ANTENNAGATEAREA                          0.072 LAYER ME4 ;
 ANTENNADIFFAREA                          0.160 LAYER ME2 ;
 ANTENNADIFFAREA                          0.160 LAYER ME3 ;
 ANTENNADIFFAREA                          0.160 LAYER ME4 ;
 ANTENNAMAXAREACAR                       21.782 LAYER ME2 ;
 ANTENNAMAXAREACAR                       24.449 LAYER ME3 ;
 ANTENNAMAXAREACAR                       27.116 LAYER ME4 ;
END DI114
PIN DO114
  DIRECTION OUTPUT ;
 PORT
  LAYER ME4 ;
  RECT 497.005 0.000 497.325 0.600 ;
  LAYER ME3 ;
  RECT 497.005 0.000 497.325 0.600 ;
  LAYER ME2 ;
  RECT 497.005 0.000 497.325 0.600 ;
  LAYER ME1 ;
  RECT 497.005 0.000 497.325 0.600 ;
 END
 ANTENNAPARTIALMETALAREA                  5.273 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME3 ;
 ANTENNADIFFAREA                          1.293 LAYER ME4 ;
END DO114
PIN DI113
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 493.563 0.000 493.883 0.600 ;
  LAYER ME3 ;
  RECT 493.563 0.000 493.883 0.600 ;
  LAYER ME2 ;
  RECT 493.563 0.000 493.883 0.600 ;
  LAYER ME1 ;
  RECT 493.563 0.000 493.883 0.600 ;
 END
 ANTENNAPARTIALMETALAREA                  1.058 LAYER ME2 ;
 ANTENNAGATEAREA                          0.072 LAYER ME2 ;
 ANTENNAGATEAREA                          0.072 LAYER ME3 ;
 ANTENNAGATEAREA                          0.072 LAYER ME4 ;
 ANTENNADIFFAREA                          0.160 LAYER ME2 ;
 ANTENNADIFFAREA                          0.160 LAYER ME3 ;
 ANTENNADIFFAREA                          0.160 LAYER ME4 ;
 ANTENNAMAXAREACAR                       21.782 LAYER ME2 ;
 ANTENNAMAXAREACAR                       24.449 LAYER ME3 ;
 ANTENNAMAXAREACAR                       27.116 LAYER ME4 ;
END DI113
PIN DO113
  DIRECTION OUTPUT ;
 PORT
  LAYER ME4 ;
  RECT 493.001 0.000 493.321 0.600 ;
  LAYER ME3 ;
  RECT 493.001 0.000 493.321 0.600 ;
  LAYER ME2 ;
  RECT 493.001 0.000 493.321 0.600 ;
  LAYER ME1 ;
  RECT 493.001 0.000 493.321 0.600 ;
 END
 ANTENNAPARTIALMETALAREA                  5.273 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME3 ;
 ANTENNADIFFAREA                          1.293 LAYER ME4 ;
END DO113
PIN DI112
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 488.997 0.000 489.317 0.600 ;
  LAYER ME3 ;
  RECT 488.997 0.000 489.317 0.600 ;
  LAYER ME2 ;
  RECT 488.997 0.000 489.317 0.600 ;
  LAYER ME1 ;
  RECT 488.997 0.000 489.317 0.600 ;
 END
 ANTENNAPARTIALMETALAREA                  0.346 LAYER ME1 ;
 ANTENNAPARTIALMETALAREA                  1.466 LAYER ME2 ;
 ANTENNAPARTIALMETALAREA                  0.508 LAYER ME3 ;
 ANTENNAGATEAREA                          0.072 LAYER ME3 ;
 ANTENNAGATEAREA                          0.072 LAYER ME4 ;
 ANTENNADIFFAREA                          0.218 LAYER ME1 ;
 ANTENNADIFFAREA                          0.218 LAYER ME2 ;
 ANTENNADIFFAREA                          0.218 LAYER ME3 ;
 ANTENNADIFFAREA                          0.218 LAYER ME4 ;
 ANTENNAMAXAREACAR                       17.267 LAYER ME3 ;
 ANTENNAMAXAREACAR                       19.933 LAYER ME4 ;
END DI112
PIN DO112
  DIRECTION OUTPUT ;
 PORT
  LAYER ME4 ;
  RECT 489.559 0.000 489.879 0.600 ;
  LAYER ME3 ;
  RECT 489.559 0.000 489.879 0.600 ;
  LAYER ME2 ;
  RECT 489.559 0.000 489.879 0.600 ;
  LAYER ME1 ;
  RECT 489.559 0.000 489.879 0.600 ;
 END
 ANTENNAPARTIALMETALAREA                  5.602 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME3 ;
 ANTENNADIFFAREA                          1.293 LAYER ME4 ;
END DO112
PIN WEB14
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 487.557 0.000 487.877 0.600 ;
  LAYER ME3 ;
  RECT 487.557 0.000 487.877 0.600 ;
  LAYER ME2 ;
  RECT 487.557 0.000 487.877 0.600 ;
  LAYER ME1 ;
  RECT 487.557 0.000 487.877 0.600 ;
 END
 ANTENNAPARTIALMETALAREA                  1.036 LAYER ME2 ;
 ANTENNAGATEAREA                          0.288 LAYER ME2 ;
 ANTENNAGATEAREA                          0.288 LAYER ME3 ;
 ANTENNAGATEAREA                          0.288 LAYER ME4 ;
 ANTENNADIFFAREA                          0.206 LAYER ME2 ;
 ANTENNADIFFAREA                          0.206 LAYER ME3 ;
 ANTENNADIFFAREA                          0.206 LAYER ME4 ;
 ANTENNAMAXAREACAR                        5.844 LAYER ME2 ;
 ANTENNAMAXAREACAR                        6.511 LAYER ME3 ;
 ANTENNAMAXAREACAR                        7.178 LAYER ME4 ;
END WEB14
PIN DI111
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 485.555 0.000 485.875 0.600 ;
  LAYER ME3 ;
  RECT 485.555 0.000 485.875 0.600 ;
  LAYER ME2 ;
  RECT 485.555 0.000 485.875 0.600 ;
  LAYER ME1 ;
  RECT 485.555 0.000 485.875 0.600 ;
 END
 ANTENNAPARTIALMETALAREA                  1.058 LAYER ME2 ;
 ANTENNAGATEAREA                          0.072 LAYER ME2 ;
 ANTENNAGATEAREA                          0.072 LAYER ME3 ;
 ANTENNAGATEAREA                          0.072 LAYER ME4 ;
 ANTENNADIFFAREA                          0.160 LAYER ME2 ;
 ANTENNADIFFAREA                          0.160 LAYER ME3 ;
 ANTENNADIFFAREA                          0.160 LAYER ME4 ;
 ANTENNAMAXAREACAR                       21.782 LAYER ME2 ;
 ANTENNAMAXAREACAR                       24.449 LAYER ME3 ;
 ANTENNAMAXAREACAR                       27.116 LAYER ME4 ;
END DI111
PIN DO111
  DIRECTION OUTPUT ;
 PORT
  LAYER ME4 ;
  RECT 484.993 0.000 485.313 0.600 ;
  LAYER ME3 ;
  RECT 484.993 0.000 485.313 0.600 ;
  LAYER ME2 ;
  RECT 484.993 0.000 485.313 0.600 ;
  LAYER ME1 ;
  RECT 484.993 0.000 485.313 0.600 ;
 END
 ANTENNAPARTIALMETALAREA                  5.273 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME3 ;
 ANTENNADIFFAREA                          1.293 LAYER ME4 ;
END DO111
PIN DI110
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 481.551 0.000 481.871 0.600 ;
  LAYER ME3 ;
  RECT 481.551 0.000 481.871 0.600 ;
  LAYER ME2 ;
  RECT 481.551 0.000 481.871 0.600 ;
  LAYER ME1 ;
  RECT 481.551 0.000 481.871 0.600 ;
 END
 ANTENNAPARTIALMETALAREA                  1.058 LAYER ME2 ;
 ANTENNAGATEAREA                          0.072 LAYER ME2 ;
 ANTENNAGATEAREA                          0.072 LAYER ME3 ;
 ANTENNAGATEAREA                          0.072 LAYER ME4 ;
 ANTENNADIFFAREA                          0.160 LAYER ME2 ;
 ANTENNADIFFAREA                          0.160 LAYER ME3 ;
 ANTENNADIFFAREA                          0.160 LAYER ME4 ;
 ANTENNAMAXAREACAR                       21.782 LAYER ME2 ;
 ANTENNAMAXAREACAR                       24.449 LAYER ME3 ;
 ANTENNAMAXAREACAR                       27.116 LAYER ME4 ;
END DI110
PIN DO110
  DIRECTION OUTPUT ;
 PORT
  LAYER ME4 ;
  RECT 480.989 0.000 481.309 0.600 ;
  LAYER ME3 ;
  RECT 480.989 0.000 481.309 0.600 ;
  LAYER ME2 ;
  RECT 480.989 0.000 481.309 0.600 ;
  LAYER ME1 ;
  RECT 480.989 0.000 481.309 0.600 ;
 END
 ANTENNAPARTIALMETALAREA                  5.273 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME3 ;
 ANTENNADIFFAREA                          1.293 LAYER ME4 ;
END DO110
PIN DI109
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 477.547 0.000 477.867 0.600 ;
  LAYER ME3 ;
  RECT 477.547 0.000 477.867 0.600 ;
  LAYER ME2 ;
  RECT 477.547 0.000 477.867 0.600 ;
  LAYER ME1 ;
  RECT 477.547 0.000 477.867 0.600 ;
 END
 ANTENNAPARTIALMETALAREA                  1.058 LAYER ME2 ;
 ANTENNAGATEAREA                          0.072 LAYER ME2 ;
 ANTENNAGATEAREA                          0.072 LAYER ME3 ;
 ANTENNAGATEAREA                          0.072 LAYER ME4 ;
 ANTENNADIFFAREA                          0.160 LAYER ME2 ;
 ANTENNADIFFAREA                          0.160 LAYER ME3 ;
 ANTENNADIFFAREA                          0.160 LAYER ME4 ;
 ANTENNAMAXAREACAR                       21.782 LAYER ME2 ;
 ANTENNAMAXAREACAR                       24.449 LAYER ME3 ;
 ANTENNAMAXAREACAR                       27.116 LAYER ME4 ;
END DI109
PIN DO109
  DIRECTION OUTPUT ;
 PORT
  LAYER ME4 ;
  RECT 476.985 0.000 477.305 0.600 ;
  LAYER ME3 ;
  RECT 476.985 0.000 477.305 0.600 ;
  LAYER ME2 ;
  RECT 476.985 0.000 477.305 0.600 ;
  LAYER ME1 ;
  RECT 476.985 0.000 477.305 0.600 ;
 END
 ANTENNAPARTIALMETALAREA                  5.273 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME3 ;
 ANTENNADIFFAREA                          1.293 LAYER ME4 ;
END DO109
PIN DI108
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 473.543 0.000 473.863 0.600 ;
  LAYER ME3 ;
  RECT 473.543 0.000 473.863 0.600 ;
  LAYER ME2 ;
  RECT 473.543 0.000 473.863 0.600 ;
  LAYER ME1 ;
  RECT 473.543 0.000 473.863 0.600 ;
 END
 ANTENNAPARTIALMETALAREA                  1.058 LAYER ME2 ;
 ANTENNAGATEAREA                          0.072 LAYER ME2 ;
 ANTENNAGATEAREA                          0.072 LAYER ME3 ;
 ANTENNAGATEAREA                          0.072 LAYER ME4 ;
 ANTENNADIFFAREA                          0.160 LAYER ME2 ;
 ANTENNADIFFAREA                          0.160 LAYER ME3 ;
 ANTENNADIFFAREA                          0.160 LAYER ME4 ;
 ANTENNAMAXAREACAR                       21.782 LAYER ME2 ;
 ANTENNAMAXAREACAR                       24.449 LAYER ME3 ;
 ANTENNAMAXAREACAR                       27.116 LAYER ME4 ;
END DI108
PIN DO108
  DIRECTION OUTPUT ;
 PORT
  LAYER ME4 ;
  RECT 472.981 0.000 473.301 0.600 ;
  LAYER ME3 ;
  RECT 472.981 0.000 473.301 0.600 ;
  LAYER ME2 ;
  RECT 472.981 0.000 473.301 0.600 ;
  LAYER ME1 ;
  RECT 472.981 0.000 473.301 0.600 ;
 END
 ANTENNAPARTIALMETALAREA                  5.273 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME3 ;
 ANTENNADIFFAREA                          1.293 LAYER ME4 ;
END DO108
PIN DI107
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 469.539 0.000 469.859 0.600 ;
  LAYER ME3 ;
  RECT 469.539 0.000 469.859 0.600 ;
  LAYER ME2 ;
  RECT 469.539 0.000 469.859 0.600 ;
  LAYER ME1 ;
  RECT 469.539 0.000 469.859 0.600 ;
 END
 ANTENNAPARTIALMETALAREA                  1.058 LAYER ME2 ;
 ANTENNAGATEAREA                          0.072 LAYER ME2 ;
 ANTENNAGATEAREA                          0.072 LAYER ME3 ;
 ANTENNAGATEAREA                          0.072 LAYER ME4 ;
 ANTENNADIFFAREA                          0.160 LAYER ME2 ;
 ANTENNADIFFAREA                          0.160 LAYER ME3 ;
 ANTENNADIFFAREA                          0.160 LAYER ME4 ;
 ANTENNAMAXAREACAR                       21.782 LAYER ME2 ;
 ANTENNAMAXAREACAR                       24.449 LAYER ME3 ;
 ANTENNAMAXAREACAR                       27.116 LAYER ME4 ;
END DI107
PIN DO107
  DIRECTION OUTPUT ;
 PORT
  LAYER ME4 ;
  RECT 468.977 0.000 469.297 0.600 ;
  LAYER ME3 ;
  RECT 468.977 0.000 469.297 0.600 ;
  LAYER ME2 ;
  RECT 468.977 0.000 469.297 0.600 ;
  LAYER ME1 ;
  RECT 468.977 0.000 469.297 0.600 ;
 END
 ANTENNAPARTIALMETALAREA                  5.273 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME3 ;
 ANTENNADIFFAREA                          1.293 LAYER ME4 ;
END DO107
PIN DI106
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 465.535 0.000 465.855 0.600 ;
  LAYER ME3 ;
  RECT 465.535 0.000 465.855 0.600 ;
  LAYER ME2 ;
  RECT 465.535 0.000 465.855 0.600 ;
  LAYER ME1 ;
  RECT 465.535 0.000 465.855 0.600 ;
 END
 ANTENNAPARTIALMETALAREA                  1.058 LAYER ME2 ;
 ANTENNAGATEAREA                          0.072 LAYER ME2 ;
 ANTENNAGATEAREA                          0.072 LAYER ME3 ;
 ANTENNAGATEAREA                          0.072 LAYER ME4 ;
 ANTENNADIFFAREA                          0.160 LAYER ME2 ;
 ANTENNADIFFAREA                          0.160 LAYER ME3 ;
 ANTENNADIFFAREA                          0.160 LAYER ME4 ;
 ANTENNAMAXAREACAR                       21.782 LAYER ME2 ;
 ANTENNAMAXAREACAR                       24.449 LAYER ME3 ;
 ANTENNAMAXAREACAR                       27.116 LAYER ME4 ;
END DI106
PIN DO106
  DIRECTION OUTPUT ;
 PORT
  LAYER ME4 ;
  RECT 464.973 0.000 465.293 0.600 ;
  LAYER ME3 ;
  RECT 464.973 0.000 465.293 0.600 ;
  LAYER ME2 ;
  RECT 464.973 0.000 465.293 0.600 ;
  LAYER ME1 ;
  RECT 464.973 0.000 465.293 0.600 ;
 END
 ANTENNAPARTIALMETALAREA                  5.273 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME3 ;
 ANTENNADIFFAREA                          1.293 LAYER ME4 ;
END DO106
PIN DI105
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 461.531 0.000 461.851 0.600 ;
  LAYER ME3 ;
  RECT 461.531 0.000 461.851 0.600 ;
  LAYER ME2 ;
  RECT 461.531 0.000 461.851 0.600 ;
  LAYER ME1 ;
  RECT 461.531 0.000 461.851 0.600 ;
 END
 ANTENNAPARTIALMETALAREA                  1.058 LAYER ME2 ;
 ANTENNAGATEAREA                          0.072 LAYER ME2 ;
 ANTENNAGATEAREA                          0.072 LAYER ME3 ;
 ANTENNAGATEAREA                          0.072 LAYER ME4 ;
 ANTENNADIFFAREA                          0.160 LAYER ME2 ;
 ANTENNADIFFAREA                          0.160 LAYER ME3 ;
 ANTENNADIFFAREA                          0.160 LAYER ME4 ;
 ANTENNAMAXAREACAR                       21.782 LAYER ME2 ;
 ANTENNAMAXAREACAR                       24.449 LAYER ME3 ;
 ANTENNAMAXAREACAR                       27.116 LAYER ME4 ;
END DI105
PIN DO105
  DIRECTION OUTPUT ;
 PORT
  LAYER ME4 ;
  RECT 460.969 0.000 461.289 0.600 ;
  LAYER ME3 ;
  RECT 460.969 0.000 461.289 0.600 ;
  LAYER ME2 ;
  RECT 460.969 0.000 461.289 0.600 ;
  LAYER ME1 ;
  RECT 460.969 0.000 461.289 0.600 ;
 END
 ANTENNAPARTIALMETALAREA                  5.273 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME3 ;
 ANTENNADIFFAREA                          1.293 LAYER ME4 ;
END DO105
PIN DI104
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 456.965 0.000 457.285 0.600 ;
  LAYER ME3 ;
  RECT 456.965 0.000 457.285 0.600 ;
  LAYER ME2 ;
  RECT 456.965 0.000 457.285 0.600 ;
  LAYER ME1 ;
  RECT 456.965 0.000 457.285 0.600 ;
 END
 ANTENNAPARTIALMETALAREA                  0.346 LAYER ME1 ;
 ANTENNAPARTIALMETALAREA                  1.466 LAYER ME2 ;
 ANTENNAPARTIALMETALAREA                  0.508 LAYER ME3 ;
 ANTENNAGATEAREA                          0.072 LAYER ME3 ;
 ANTENNAGATEAREA                          0.072 LAYER ME4 ;
 ANTENNADIFFAREA                          0.218 LAYER ME1 ;
 ANTENNADIFFAREA                          0.218 LAYER ME2 ;
 ANTENNADIFFAREA                          0.218 LAYER ME3 ;
 ANTENNADIFFAREA                          0.218 LAYER ME4 ;
 ANTENNAMAXAREACAR                       17.267 LAYER ME3 ;
 ANTENNAMAXAREACAR                       19.933 LAYER ME4 ;
END DI104
PIN DO104
  DIRECTION OUTPUT ;
 PORT
  LAYER ME4 ;
  RECT 457.527 0.000 457.847 0.600 ;
  LAYER ME3 ;
  RECT 457.527 0.000 457.847 0.600 ;
  LAYER ME2 ;
  RECT 457.527 0.000 457.847 0.600 ;
  LAYER ME1 ;
  RECT 457.527 0.000 457.847 0.600 ;
 END
 ANTENNAPARTIALMETALAREA                  5.602 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME3 ;
 ANTENNADIFFAREA                          1.293 LAYER ME4 ;
END DO104
PIN WEB13
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 455.525 0.000 455.845 0.600 ;
  LAYER ME3 ;
  RECT 455.525 0.000 455.845 0.600 ;
  LAYER ME2 ;
  RECT 455.525 0.000 455.845 0.600 ;
  LAYER ME1 ;
  RECT 455.525 0.000 455.845 0.600 ;
 END
 ANTENNAPARTIALMETALAREA                  1.036 LAYER ME2 ;
 ANTENNAGATEAREA                          0.288 LAYER ME2 ;
 ANTENNAGATEAREA                          0.288 LAYER ME3 ;
 ANTENNAGATEAREA                          0.288 LAYER ME4 ;
 ANTENNADIFFAREA                          0.206 LAYER ME2 ;
 ANTENNADIFFAREA                          0.206 LAYER ME3 ;
 ANTENNADIFFAREA                          0.206 LAYER ME4 ;
 ANTENNAMAXAREACAR                        5.844 LAYER ME2 ;
 ANTENNAMAXAREACAR                        6.511 LAYER ME3 ;
 ANTENNAMAXAREACAR                        7.178 LAYER ME4 ;
END WEB13
PIN DI103
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 453.523 0.000 453.843 0.600 ;
  LAYER ME3 ;
  RECT 453.523 0.000 453.843 0.600 ;
  LAYER ME2 ;
  RECT 453.523 0.000 453.843 0.600 ;
  LAYER ME1 ;
  RECT 453.523 0.000 453.843 0.600 ;
 END
 ANTENNAPARTIALMETALAREA                  1.058 LAYER ME2 ;
 ANTENNAGATEAREA                          0.072 LAYER ME2 ;
 ANTENNAGATEAREA                          0.072 LAYER ME3 ;
 ANTENNAGATEAREA                          0.072 LAYER ME4 ;
 ANTENNADIFFAREA                          0.160 LAYER ME2 ;
 ANTENNADIFFAREA                          0.160 LAYER ME3 ;
 ANTENNADIFFAREA                          0.160 LAYER ME4 ;
 ANTENNAMAXAREACAR                       21.782 LAYER ME2 ;
 ANTENNAMAXAREACAR                       24.449 LAYER ME3 ;
 ANTENNAMAXAREACAR                       27.116 LAYER ME4 ;
END DI103
PIN DO103
  DIRECTION OUTPUT ;
 PORT
  LAYER ME4 ;
  RECT 452.961 0.000 453.281 0.600 ;
  LAYER ME3 ;
  RECT 452.961 0.000 453.281 0.600 ;
  LAYER ME2 ;
  RECT 452.961 0.000 453.281 0.600 ;
  LAYER ME1 ;
  RECT 452.961 0.000 453.281 0.600 ;
 END
 ANTENNAPARTIALMETALAREA                  5.273 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME3 ;
 ANTENNADIFFAREA                          1.293 LAYER ME4 ;
END DO103
PIN DI102
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 449.519 0.000 449.839 0.600 ;
  LAYER ME3 ;
  RECT 449.519 0.000 449.839 0.600 ;
  LAYER ME2 ;
  RECT 449.519 0.000 449.839 0.600 ;
  LAYER ME1 ;
  RECT 449.519 0.000 449.839 0.600 ;
 END
 ANTENNAPARTIALMETALAREA                  1.058 LAYER ME2 ;
 ANTENNAGATEAREA                          0.072 LAYER ME2 ;
 ANTENNAGATEAREA                          0.072 LAYER ME3 ;
 ANTENNAGATEAREA                          0.072 LAYER ME4 ;
 ANTENNADIFFAREA                          0.160 LAYER ME2 ;
 ANTENNADIFFAREA                          0.160 LAYER ME3 ;
 ANTENNADIFFAREA                          0.160 LAYER ME4 ;
 ANTENNAMAXAREACAR                       21.782 LAYER ME2 ;
 ANTENNAMAXAREACAR                       24.449 LAYER ME3 ;
 ANTENNAMAXAREACAR                       27.116 LAYER ME4 ;
END DI102
PIN DO102
  DIRECTION OUTPUT ;
 PORT
  LAYER ME4 ;
  RECT 448.957 0.000 449.277 0.600 ;
  LAYER ME3 ;
  RECT 448.957 0.000 449.277 0.600 ;
  LAYER ME2 ;
  RECT 448.957 0.000 449.277 0.600 ;
  LAYER ME1 ;
  RECT 448.957 0.000 449.277 0.600 ;
 END
 ANTENNAPARTIALMETALAREA                  5.273 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME3 ;
 ANTENNADIFFAREA                          1.293 LAYER ME4 ;
END DO102
PIN DI101
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 445.515 0.000 445.835 0.600 ;
  LAYER ME3 ;
  RECT 445.515 0.000 445.835 0.600 ;
  LAYER ME2 ;
  RECT 445.515 0.000 445.835 0.600 ;
  LAYER ME1 ;
  RECT 445.515 0.000 445.835 0.600 ;
 END
 ANTENNAPARTIALMETALAREA                  1.058 LAYER ME2 ;
 ANTENNAGATEAREA                          0.072 LAYER ME2 ;
 ANTENNAGATEAREA                          0.072 LAYER ME3 ;
 ANTENNAGATEAREA                          0.072 LAYER ME4 ;
 ANTENNADIFFAREA                          0.160 LAYER ME2 ;
 ANTENNADIFFAREA                          0.160 LAYER ME3 ;
 ANTENNADIFFAREA                          0.160 LAYER ME4 ;
 ANTENNAMAXAREACAR                       21.782 LAYER ME2 ;
 ANTENNAMAXAREACAR                       24.449 LAYER ME3 ;
 ANTENNAMAXAREACAR                       27.116 LAYER ME4 ;
END DI101
PIN DO101
  DIRECTION OUTPUT ;
 PORT
  LAYER ME4 ;
  RECT 444.953 0.000 445.273 0.600 ;
  LAYER ME3 ;
  RECT 444.953 0.000 445.273 0.600 ;
  LAYER ME2 ;
  RECT 444.953 0.000 445.273 0.600 ;
  LAYER ME1 ;
  RECT 444.953 0.000 445.273 0.600 ;
 END
 ANTENNAPARTIALMETALAREA                  5.273 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME3 ;
 ANTENNADIFFAREA                          1.293 LAYER ME4 ;
END DO101
PIN DI100
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 441.511 0.000 441.831 0.600 ;
  LAYER ME3 ;
  RECT 441.511 0.000 441.831 0.600 ;
  LAYER ME2 ;
  RECT 441.511 0.000 441.831 0.600 ;
  LAYER ME1 ;
  RECT 441.511 0.000 441.831 0.600 ;
 END
 ANTENNAPARTIALMETALAREA                  1.058 LAYER ME2 ;
 ANTENNAGATEAREA                          0.072 LAYER ME2 ;
 ANTENNAGATEAREA                          0.072 LAYER ME3 ;
 ANTENNAGATEAREA                          0.072 LAYER ME4 ;
 ANTENNADIFFAREA                          0.160 LAYER ME2 ;
 ANTENNADIFFAREA                          0.160 LAYER ME3 ;
 ANTENNADIFFAREA                          0.160 LAYER ME4 ;
 ANTENNAMAXAREACAR                       21.782 LAYER ME2 ;
 ANTENNAMAXAREACAR                       24.449 LAYER ME3 ;
 ANTENNAMAXAREACAR                       27.116 LAYER ME4 ;
END DI100
PIN DO100
  DIRECTION OUTPUT ;
 PORT
  LAYER ME4 ;
  RECT 440.949 0.000 441.269 0.600 ;
  LAYER ME3 ;
  RECT 440.949 0.000 441.269 0.600 ;
  LAYER ME2 ;
  RECT 440.949 0.000 441.269 0.600 ;
  LAYER ME1 ;
  RECT 440.949 0.000 441.269 0.600 ;
 END
 ANTENNAPARTIALMETALAREA                  5.273 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME3 ;
 ANTENNADIFFAREA                          1.293 LAYER ME4 ;
END DO100
PIN DI99
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 437.507 0.000 437.827 0.600 ;
  LAYER ME3 ;
  RECT 437.507 0.000 437.827 0.600 ;
  LAYER ME2 ;
  RECT 437.507 0.000 437.827 0.600 ;
  LAYER ME1 ;
  RECT 437.507 0.000 437.827 0.600 ;
 END
 ANTENNAPARTIALMETALAREA                  1.058 LAYER ME2 ;
 ANTENNAGATEAREA                          0.072 LAYER ME2 ;
 ANTENNAGATEAREA                          0.072 LAYER ME3 ;
 ANTENNAGATEAREA                          0.072 LAYER ME4 ;
 ANTENNADIFFAREA                          0.160 LAYER ME2 ;
 ANTENNADIFFAREA                          0.160 LAYER ME3 ;
 ANTENNADIFFAREA                          0.160 LAYER ME4 ;
 ANTENNAMAXAREACAR                       21.782 LAYER ME2 ;
 ANTENNAMAXAREACAR                       24.449 LAYER ME3 ;
 ANTENNAMAXAREACAR                       27.116 LAYER ME4 ;
END DI99
PIN DO99
  DIRECTION OUTPUT ;
 PORT
  LAYER ME4 ;
  RECT 436.945 0.000 437.265 0.600 ;
  LAYER ME3 ;
  RECT 436.945 0.000 437.265 0.600 ;
  LAYER ME2 ;
  RECT 436.945 0.000 437.265 0.600 ;
  LAYER ME1 ;
  RECT 436.945 0.000 437.265 0.600 ;
 END
 ANTENNAPARTIALMETALAREA                  5.273 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME3 ;
 ANTENNADIFFAREA                          1.293 LAYER ME4 ;
END DO99
PIN DI98
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 433.503 0.000 433.823 0.600 ;
  LAYER ME3 ;
  RECT 433.503 0.000 433.823 0.600 ;
  LAYER ME2 ;
  RECT 433.503 0.000 433.823 0.600 ;
  LAYER ME1 ;
  RECT 433.503 0.000 433.823 0.600 ;
 END
 ANTENNAPARTIALMETALAREA                  1.058 LAYER ME2 ;
 ANTENNAGATEAREA                          0.072 LAYER ME2 ;
 ANTENNAGATEAREA                          0.072 LAYER ME3 ;
 ANTENNAGATEAREA                          0.072 LAYER ME4 ;
 ANTENNADIFFAREA                          0.160 LAYER ME2 ;
 ANTENNADIFFAREA                          0.160 LAYER ME3 ;
 ANTENNADIFFAREA                          0.160 LAYER ME4 ;
 ANTENNAMAXAREACAR                       21.782 LAYER ME2 ;
 ANTENNAMAXAREACAR                       24.449 LAYER ME3 ;
 ANTENNAMAXAREACAR                       27.116 LAYER ME4 ;
END DI98
PIN DO98
  DIRECTION OUTPUT ;
 PORT
  LAYER ME4 ;
  RECT 432.941 0.000 433.261 0.600 ;
  LAYER ME3 ;
  RECT 432.941 0.000 433.261 0.600 ;
  LAYER ME2 ;
  RECT 432.941 0.000 433.261 0.600 ;
  LAYER ME1 ;
  RECT 432.941 0.000 433.261 0.600 ;
 END
 ANTENNAPARTIALMETALAREA                  5.273 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME3 ;
 ANTENNADIFFAREA                          1.293 LAYER ME4 ;
END DO98
PIN DI97
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 429.499 0.000 429.819 0.600 ;
  LAYER ME3 ;
  RECT 429.499 0.000 429.819 0.600 ;
  LAYER ME2 ;
  RECT 429.499 0.000 429.819 0.600 ;
  LAYER ME1 ;
  RECT 429.499 0.000 429.819 0.600 ;
 END
 ANTENNAPARTIALMETALAREA                  1.058 LAYER ME2 ;
 ANTENNAGATEAREA                          0.072 LAYER ME2 ;
 ANTENNAGATEAREA                          0.072 LAYER ME3 ;
 ANTENNAGATEAREA                          0.072 LAYER ME4 ;
 ANTENNADIFFAREA                          0.160 LAYER ME2 ;
 ANTENNADIFFAREA                          0.160 LAYER ME3 ;
 ANTENNADIFFAREA                          0.160 LAYER ME4 ;
 ANTENNAMAXAREACAR                       21.782 LAYER ME2 ;
 ANTENNAMAXAREACAR                       24.449 LAYER ME3 ;
 ANTENNAMAXAREACAR                       27.116 LAYER ME4 ;
END DI97
PIN DO97
  DIRECTION OUTPUT ;
 PORT
  LAYER ME4 ;
  RECT 428.937 0.000 429.257 0.600 ;
  LAYER ME3 ;
  RECT 428.937 0.000 429.257 0.600 ;
  LAYER ME2 ;
  RECT 428.937 0.000 429.257 0.600 ;
  LAYER ME1 ;
  RECT 428.937 0.000 429.257 0.600 ;
 END
 ANTENNAPARTIALMETALAREA                  5.273 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME3 ;
 ANTENNADIFFAREA                          1.293 LAYER ME4 ;
END DO97
PIN DI96
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 424.933 0.000 425.253 0.600 ;
  LAYER ME3 ;
  RECT 424.933 0.000 425.253 0.600 ;
  LAYER ME2 ;
  RECT 424.933 0.000 425.253 0.600 ;
  LAYER ME1 ;
  RECT 424.933 0.000 425.253 0.600 ;
 END
 ANTENNAPARTIALMETALAREA                  0.346 LAYER ME1 ;
 ANTENNAPARTIALMETALAREA                  1.466 LAYER ME2 ;
 ANTENNAPARTIALMETALAREA                  0.508 LAYER ME3 ;
 ANTENNAGATEAREA                          0.072 LAYER ME3 ;
 ANTENNAGATEAREA                          0.072 LAYER ME4 ;
 ANTENNADIFFAREA                          0.218 LAYER ME1 ;
 ANTENNADIFFAREA                          0.218 LAYER ME2 ;
 ANTENNADIFFAREA                          0.218 LAYER ME3 ;
 ANTENNADIFFAREA                          0.218 LAYER ME4 ;
 ANTENNAMAXAREACAR                       17.267 LAYER ME3 ;
 ANTENNAMAXAREACAR                       19.933 LAYER ME4 ;
END DI96
PIN DO96
  DIRECTION OUTPUT ;
 PORT
  LAYER ME4 ;
  RECT 425.495 0.000 425.815 0.600 ;
  LAYER ME3 ;
  RECT 425.495 0.000 425.815 0.600 ;
  LAYER ME2 ;
  RECT 425.495 0.000 425.815 0.600 ;
  LAYER ME1 ;
  RECT 425.495 0.000 425.815 0.600 ;
 END
 ANTENNAPARTIALMETALAREA                  5.602 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME3 ;
 ANTENNADIFFAREA                          1.293 LAYER ME4 ;
END DO96
PIN WEB12
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 423.493 0.000 423.813 0.600 ;
  LAYER ME3 ;
  RECT 423.493 0.000 423.813 0.600 ;
  LAYER ME2 ;
  RECT 423.493 0.000 423.813 0.600 ;
  LAYER ME1 ;
  RECT 423.493 0.000 423.813 0.600 ;
 END
 ANTENNAPARTIALMETALAREA                  1.036 LAYER ME2 ;
 ANTENNAGATEAREA                          0.288 LAYER ME2 ;
 ANTENNAGATEAREA                          0.288 LAYER ME3 ;
 ANTENNAGATEAREA                          0.288 LAYER ME4 ;
 ANTENNADIFFAREA                          0.206 LAYER ME2 ;
 ANTENNADIFFAREA                          0.206 LAYER ME3 ;
 ANTENNADIFFAREA                          0.206 LAYER ME4 ;
 ANTENNAMAXAREACAR                        5.844 LAYER ME2 ;
 ANTENNAMAXAREACAR                        6.511 LAYER ME3 ;
 ANTENNAMAXAREACAR                        7.178 LAYER ME4 ;
END WEB12
PIN DI95
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 421.491 0.000 421.811 0.600 ;
  LAYER ME3 ;
  RECT 421.491 0.000 421.811 0.600 ;
  LAYER ME2 ;
  RECT 421.491 0.000 421.811 0.600 ;
  LAYER ME1 ;
  RECT 421.491 0.000 421.811 0.600 ;
 END
 ANTENNAPARTIALMETALAREA                  1.058 LAYER ME2 ;
 ANTENNAGATEAREA                          0.072 LAYER ME2 ;
 ANTENNAGATEAREA                          0.072 LAYER ME3 ;
 ANTENNAGATEAREA                          0.072 LAYER ME4 ;
 ANTENNADIFFAREA                          0.160 LAYER ME2 ;
 ANTENNADIFFAREA                          0.160 LAYER ME3 ;
 ANTENNADIFFAREA                          0.160 LAYER ME4 ;
 ANTENNAMAXAREACAR                       21.782 LAYER ME2 ;
 ANTENNAMAXAREACAR                       24.449 LAYER ME3 ;
 ANTENNAMAXAREACAR                       27.116 LAYER ME4 ;
END DI95
PIN DO95
  DIRECTION OUTPUT ;
 PORT
  LAYER ME4 ;
  RECT 420.929 0.000 421.249 0.600 ;
  LAYER ME3 ;
  RECT 420.929 0.000 421.249 0.600 ;
  LAYER ME2 ;
  RECT 420.929 0.000 421.249 0.600 ;
  LAYER ME1 ;
  RECT 420.929 0.000 421.249 0.600 ;
 END
 ANTENNAPARTIALMETALAREA                  5.273 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME3 ;
 ANTENNADIFFAREA                          1.293 LAYER ME4 ;
END DO95
PIN DI94
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 417.487 0.000 417.807 0.600 ;
  LAYER ME3 ;
  RECT 417.487 0.000 417.807 0.600 ;
  LAYER ME2 ;
  RECT 417.487 0.000 417.807 0.600 ;
  LAYER ME1 ;
  RECT 417.487 0.000 417.807 0.600 ;
 END
 ANTENNAPARTIALMETALAREA                  1.058 LAYER ME2 ;
 ANTENNAGATEAREA                          0.072 LAYER ME2 ;
 ANTENNAGATEAREA                          0.072 LAYER ME3 ;
 ANTENNAGATEAREA                          0.072 LAYER ME4 ;
 ANTENNADIFFAREA                          0.160 LAYER ME2 ;
 ANTENNADIFFAREA                          0.160 LAYER ME3 ;
 ANTENNADIFFAREA                          0.160 LAYER ME4 ;
 ANTENNAMAXAREACAR                       21.782 LAYER ME2 ;
 ANTENNAMAXAREACAR                       24.449 LAYER ME3 ;
 ANTENNAMAXAREACAR                       27.116 LAYER ME4 ;
END DI94
PIN DO94
  DIRECTION OUTPUT ;
 PORT
  LAYER ME4 ;
  RECT 416.925 0.000 417.245 0.600 ;
  LAYER ME3 ;
  RECT 416.925 0.000 417.245 0.600 ;
  LAYER ME2 ;
  RECT 416.925 0.000 417.245 0.600 ;
  LAYER ME1 ;
  RECT 416.925 0.000 417.245 0.600 ;
 END
 ANTENNAPARTIALMETALAREA                  5.273 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME3 ;
 ANTENNADIFFAREA                          1.293 LAYER ME4 ;
END DO94
PIN DI93
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 413.483 0.000 413.803 0.600 ;
  LAYER ME3 ;
  RECT 413.483 0.000 413.803 0.600 ;
  LAYER ME2 ;
  RECT 413.483 0.000 413.803 0.600 ;
  LAYER ME1 ;
  RECT 413.483 0.000 413.803 0.600 ;
 END
 ANTENNAPARTIALMETALAREA                  1.058 LAYER ME2 ;
 ANTENNAGATEAREA                          0.072 LAYER ME2 ;
 ANTENNAGATEAREA                          0.072 LAYER ME3 ;
 ANTENNAGATEAREA                          0.072 LAYER ME4 ;
 ANTENNADIFFAREA                          0.160 LAYER ME2 ;
 ANTENNADIFFAREA                          0.160 LAYER ME3 ;
 ANTENNADIFFAREA                          0.160 LAYER ME4 ;
 ANTENNAMAXAREACAR                       21.782 LAYER ME2 ;
 ANTENNAMAXAREACAR                       24.449 LAYER ME3 ;
 ANTENNAMAXAREACAR                       27.116 LAYER ME4 ;
END DI93
PIN DO93
  DIRECTION OUTPUT ;
 PORT
  LAYER ME4 ;
  RECT 412.921 0.000 413.241 0.600 ;
  LAYER ME3 ;
  RECT 412.921 0.000 413.241 0.600 ;
  LAYER ME2 ;
  RECT 412.921 0.000 413.241 0.600 ;
  LAYER ME1 ;
  RECT 412.921 0.000 413.241 0.600 ;
 END
 ANTENNAPARTIALMETALAREA                  5.273 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME3 ;
 ANTENNADIFFAREA                          1.293 LAYER ME4 ;
END DO93
PIN DI92
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 409.479 0.000 409.799 0.600 ;
  LAYER ME3 ;
  RECT 409.479 0.000 409.799 0.600 ;
  LAYER ME2 ;
  RECT 409.479 0.000 409.799 0.600 ;
  LAYER ME1 ;
  RECT 409.479 0.000 409.799 0.600 ;
 END
 ANTENNAPARTIALMETALAREA                  1.058 LAYER ME2 ;
 ANTENNAGATEAREA                          0.072 LAYER ME2 ;
 ANTENNAGATEAREA                          0.072 LAYER ME3 ;
 ANTENNAGATEAREA                          0.072 LAYER ME4 ;
 ANTENNADIFFAREA                          0.160 LAYER ME2 ;
 ANTENNADIFFAREA                          0.160 LAYER ME3 ;
 ANTENNADIFFAREA                          0.160 LAYER ME4 ;
 ANTENNAMAXAREACAR                       21.782 LAYER ME2 ;
 ANTENNAMAXAREACAR                       24.449 LAYER ME3 ;
 ANTENNAMAXAREACAR                       27.116 LAYER ME4 ;
END DI92
PIN DO92
  DIRECTION OUTPUT ;
 PORT
  LAYER ME4 ;
  RECT 408.917 0.000 409.237 0.600 ;
  LAYER ME3 ;
  RECT 408.917 0.000 409.237 0.600 ;
  LAYER ME2 ;
  RECT 408.917 0.000 409.237 0.600 ;
  LAYER ME1 ;
  RECT 408.917 0.000 409.237 0.600 ;
 END
 ANTENNAPARTIALMETALAREA                  5.273 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME3 ;
 ANTENNADIFFAREA                          1.293 LAYER ME4 ;
END DO92
PIN DI91
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 405.475 0.000 405.795 0.600 ;
  LAYER ME3 ;
  RECT 405.475 0.000 405.795 0.600 ;
  LAYER ME2 ;
  RECT 405.475 0.000 405.795 0.600 ;
  LAYER ME1 ;
  RECT 405.475 0.000 405.795 0.600 ;
 END
 ANTENNAPARTIALMETALAREA                  1.058 LAYER ME2 ;
 ANTENNAGATEAREA                          0.072 LAYER ME2 ;
 ANTENNAGATEAREA                          0.072 LAYER ME3 ;
 ANTENNAGATEAREA                          0.072 LAYER ME4 ;
 ANTENNADIFFAREA                          0.160 LAYER ME2 ;
 ANTENNADIFFAREA                          0.160 LAYER ME3 ;
 ANTENNADIFFAREA                          0.160 LAYER ME4 ;
 ANTENNAMAXAREACAR                       21.782 LAYER ME2 ;
 ANTENNAMAXAREACAR                       24.449 LAYER ME3 ;
 ANTENNAMAXAREACAR                       27.116 LAYER ME4 ;
END DI91
PIN DO91
  DIRECTION OUTPUT ;
 PORT
  LAYER ME4 ;
  RECT 404.913 0.000 405.233 0.600 ;
  LAYER ME3 ;
  RECT 404.913 0.000 405.233 0.600 ;
  LAYER ME2 ;
  RECT 404.913 0.000 405.233 0.600 ;
  LAYER ME1 ;
  RECT 404.913 0.000 405.233 0.600 ;
 END
 ANTENNAPARTIALMETALAREA                  5.273 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME3 ;
 ANTENNADIFFAREA                          1.293 LAYER ME4 ;
END DO91
PIN DI90
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 401.471 0.000 401.791 0.600 ;
  LAYER ME3 ;
  RECT 401.471 0.000 401.791 0.600 ;
  LAYER ME2 ;
  RECT 401.471 0.000 401.791 0.600 ;
  LAYER ME1 ;
  RECT 401.471 0.000 401.791 0.600 ;
 END
 ANTENNAPARTIALMETALAREA                  1.058 LAYER ME2 ;
 ANTENNAGATEAREA                          0.072 LAYER ME2 ;
 ANTENNAGATEAREA                          0.072 LAYER ME3 ;
 ANTENNAGATEAREA                          0.072 LAYER ME4 ;
 ANTENNADIFFAREA                          0.160 LAYER ME2 ;
 ANTENNADIFFAREA                          0.160 LAYER ME3 ;
 ANTENNADIFFAREA                          0.160 LAYER ME4 ;
 ANTENNAMAXAREACAR                       21.782 LAYER ME2 ;
 ANTENNAMAXAREACAR                       24.449 LAYER ME3 ;
 ANTENNAMAXAREACAR                       27.116 LAYER ME4 ;
END DI90
PIN DO90
  DIRECTION OUTPUT ;
 PORT
  LAYER ME4 ;
  RECT 400.909 0.000 401.229 0.600 ;
  LAYER ME3 ;
  RECT 400.909 0.000 401.229 0.600 ;
  LAYER ME2 ;
  RECT 400.909 0.000 401.229 0.600 ;
  LAYER ME1 ;
  RECT 400.909 0.000 401.229 0.600 ;
 END
 ANTENNAPARTIALMETALAREA                  5.273 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME3 ;
 ANTENNADIFFAREA                          1.293 LAYER ME4 ;
END DO90
PIN DI89
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 397.467 0.000 397.787 0.600 ;
  LAYER ME3 ;
  RECT 397.467 0.000 397.787 0.600 ;
  LAYER ME2 ;
  RECT 397.467 0.000 397.787 0.600 ;
  LAYER ME1 ;
  RECT 397.467 0.000 397.787 0.600 ;
 END
 ANTENNAPARTIALMETALAREA                  1.058 LAYER ME2 ;
 ANTENNAGATEAREA                          0.072 LAYER ME2 ;
 ANTENNAGATEAREA                          0.072 LAYER ME3 ;
 ANTENNAGATEAREA                          0.072 LAYER ME4 ;
 ANTENNADIFFAREA                          0.160 LAYER ME2 ;
 ANTENNADIFFAREA                          0.160 LAYER ME3 ;
 ANTENNADIFFAREA                          0.160 LAYER ME4 ;
 ANTENNAMAXAREACAR                       21.782 LAYER ME2 ;
 ANTENNAMAXAREACAR                       24.449 LAYER ME3 ;
 ANTENNAMAXAREACAR                       27.116 LAYER ME4 ;
END DI89
PIN DO89
  DIRECTION OUTPUT ;
 PORT
  LAYER ME4 ;
  RECT 396.905 0.000 397.225 0.600 ;
  LAYER ME3 ;
  RECT 396.905 0.000 397.225 0.600 ;
  LAYER ME2 ;
  RECT 396.905 0.000 397.225 0.600 ;
  LAYER ME1 ;
  RECT 396.905 0.000 397.225 0.600 ;
 END
 ANTENNAPARTIALMETALAREA                  5.273 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME3 ;
 ANTENNADIFFAREA                          1.293 LAYER ME4 ;
END DO89
PIN DI88
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 392.901 0.000 393.221 0.600 ;
  LAYER ME3 ;
  RECT 392.901 0.000 393.221 0.600 ;
  LAYER ME2 ;
  RECT 392.901 0.000 393.221 0.600 ;
  LAYER ME1 ;
  RECT 392.901 0.000 393.221 0.600 ;
 END
 ANTENNAPARTIALMETALAREA                  0.346 LAYER ME1 ;
 ANTENNAPARTIALMETALAREA                  1.466 LAYER ME2 ;
 ANTENNAPARTIALMETALAREA                  0.508 LAYER ME3 ;
 ANTENNAGATEAREA                          0.072 LAYER ME3 ;
 ANTENNAGATEAREA                          0.072 LAYER ME4 ;
 ANTENNADIFFAREA                          0.218 LAYER ME1 ;
 ANTENNADIFFAREA                          0.218 LAYER ME2 ;
 ANTENNADIFFAREA                          0.218 LAYER ME3 ;
 ANTENNADIFFAREA                          0.218 LAYER ME4 ;
 ANTENNAMAXAREACAR                       17.267 LAYER ME3 ;
 ANTENNAMAXAREACAR                       19.933 LAYER ME4 ;
END DI88
PIN DO88
  DIRECTION OUTPUT ;
 PORT
  LAYER ME4 ;
  RECT 393.463 0.000 393.783 0.600 ;
  LAYER ME3 ;
  RECT 393.463 0.000 393.783 0.600 ;
  LAYER ME2 ;
  RECT 393.463 0.000 393.783 0.600 ;
  LAYER ME1 ;
  RECT 393.463 0.000 393.783 0.600 ;
 END
 ANTENNAPARTIALMETALAREA                  5.602 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME3 ;
 ANTENNADIFFAREA                          1.293 LAYER ME4 ;
END DO88
PIN WEB11
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 391.461 0.000 391.781 0.600 ;
  LAYER ME3 ;
  RECT 391.461 0.000 391.781 0.600 ;
  LAYER ME2 ;
  RECT 391.461 0.000 391.781 0.600 ;
  LAYER ME1 ;
  RECT 391.461 0.000 391.781 0.600 ;
 END
 ANTENNAPARTIALMETALAREA                  1.036 LAYER ME2 ;
 ANTENNAGATEAREA                          0.288 LAYER ME2 ;
 ANTENNAGATEAREA                          0.288 LAYER ME3 ;
 ANTENNAGATEAREA                          0.288 LAYER ME4 ;
 ANTENNADIFFAREA                          0.206 LAYER ME2 ;
 ANTENNADIFFAREA                          0.206 LAYER ME3 ;
 ANTENNADIFFAREA                          0.206 LAYER ME4 ;
 ANTENNAMAXAREACAR                        5.844 LAYER ME2 ;
 ANTENNAMAXAREACAR                        6.511 LAYER ME3 ;
 ANTENNAMAXAREACAR                        7.178 LAYER ME4 ;
END WEB11
PIN DI87
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 389.459 0.000 389.779 0.600 ;
  LAYER ME3 ;
  RECT 389.459 0.000 389.779 0.600 ;
  LAYER ME2 ;
  RECT 389.459 0.000 389.779 0.600 ;
  LAYER ME1 ;
  RECT 389.459 0.000 389.779 0.600 ;
 END
 ANTENNAPARTIALMETALAREA                  1.058 LAYER ME2 ;
 ANTENNAGATEAREA                          0.072 LAYER ME2 ;
 ANTENNAGATEAREA                          0.072 LAYER ME3 ;
 ANTENNAGATEAREA                          0.072 LAYER ME4 ;
 ANTENNADIFFAREA                          0.160 LAYER ME2 ;
 ANTENNADIFFAREA                          0.160 LAYER ME3 ;
 ANTENNADIFFAREA                          0.160 LAYER ME4 ;
 ANTENNAMAXAREACAR                       21.782 LAYER ME2 ;
 ANTENNAMAXAREACAR                       24.449 LAYER ME3 ;
 ANTENNAMAXAREACAR                       27.116 LAYER ME4 ;
END DI87
PIN DO87
  DIRECTION OUTPUT ;
 PORT
  LAYER ME4 ;
  RECT 388.897 0.000 389.217 0.600 ;
  LAYER ME3 ;
  RECT 388.897 0.000 389.217 0.600 ;
  LAYER ME2 ;
  RECT 388.897 0.000 389.217 0.600 ;
  LAYER ME1 ;
  RECT 388.897 0.000 389.217 0.600 ;
 END
 ANTENNAPARTIALMETALAREA                  5.273 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME3 ;
 ANTENNADIFFAREA                          1.293 LAYER ME4 ;
END DO87
PIN DI86
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 385.455 0.000 385.775 0.600 ;
  LAYER ME3 ;
  RECT 385.455 0.000 385.775 0.600 ;
  LAYER ME2 ;
  RECT 385.455 0.000 385.775 0.600 ;
  LAYER ME1 ;
  RECT 385.455 0.000 385.775 0.600 ;
 END
 ANTENNAPARTIALMETALAREA                  1.058 LAYER ME2 ;
 ANTENNAGATEAREA                          0.072 LAYER ME2 ;
 ANTENNAGATEAREA                          0.072 LAYER ME3 ;
 ANTENNAGATEAREA                          0.072 LAYER ME4 ;
 ANTENNADIFFAREA                          0.160 LAYER ME2 ;
 ANTENNADIFFAREA                          0.160 LAYER ME3 ;
 ANTENNADIFFAREA                          0.160 LAYER ME4 ;
 ANTENNAMAXAREACAR                       21.782 LAYER ME2 ;
 ANTENNAMAXAREACAR                       24.449 LAYER ME3 ;
 ANTENNAMAXAREACAR                       27.116 LAYER ME4 ;
END DI86
PIN DO86
  DIRECTION OUTPUT ;
 PORT
  LAYER ME4 ;
  RECT 384.893 0.000 385.213 0.600 ;
  LAYER ME3 ;
  RECT 384.893 0.000 385.213 0.600 ;
  LAYER ME2 ;
  RECT 384.893 0.000 385.213 0.600 ;
  LAYER ME1 ;
  RECT 384.893 0.000 385.213 0.600 ;
 END
 ANTENNAPARTIALMETALAREA                  5.273 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME3 ;
 ANTENNADIFFAREA                          1.293 LAYER ME4 ;
END DO86
PIN DI85
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 381.451 0.000 381.771 0.600 ;
  LAYER ME3 ;
  RECT 381.451 0.000 381.771 0.600 ;
  LAYER ME2 ;
  RECT 381.451 0.000 381.771 0.600 ;
  LAYER ME1 ;
  RECT 381.451 0.000 381.771 0.600 ;
 END
 ANTENNAPARTIALMETALAREA                  1.058 LAYER ME2 ;
 ANTENNAGATEAREA                          0.072 LAYER ME2 ;
 ANTENNAGATEAREA                          0.072 LAYER ME3 ;
 ANTENNAGATEAREA                          0.072 LAYER ME4 ;
 ANTENNADIFFAREA                          0.160 LAYER ME2 ;
 ANTENNADIFFAREA                          0.160 LAYER ME3 ;
 ANTENNADIFFAREA                          0.160 LAYER ME4 ;
 ANTENNAMAXAREACAR                       21.782 LAYER ME2 ;
 ANTENNAMAXAREACAR                       24.449 LAYER ME3 ;
 ANTENNAMAXAREACAR                       27.116 LAYER ME4 ;
END DI85
PIN DO85
  DIRECTION OUTPUT ;
 PORT
  LAYER ME4 ;
  RECT 380.889 0.000 381.209 0.600 ;
  LAYER ME3 ;
  RECT 380.889 0.000 381.209 0.600 ;
  LAYER ME2 ;
  RECT 380.889 0.000 381.209 0.600 ;
  LAYER ME1 ;
  RECT 380.889 0.000 381.209 0.600 ;
 END
 ANTENNAPARTIALMETALAREA                  5.273 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME3 ;
 ANTENNADIFFAREA                          1.293 LAYER ME4 ;
END DO85
PIN DI84
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 377.447 0.000 377.767 0.600 ;
  LAYER ME3 ;
  RECT 377.447 0.000 377.767 0.600 ;
  LAYER ME2 ;
  RECT 377.447 0.000 377.767 0.600 ;
  LAYER ME1 ;
  RECT 377.447 0.000 377.767 0.600 ;
 END
 ANTENNAPARTIALMETALAREA                  1.058 LAYER ME2 ;
 ANTENNAGATEAREA                          0.072 LAYER ME2 ;
 ANTENNAGATEAREA                          0.072 LAYER ME3 ;
 ANTENNAGATEAREA                          0.072 LAYER ME4 ;
 ANTENNADIFFAREA                          0.160 LAYER ME2 ;
 ANTENNADIFFAREA                          0.160 LAYER ME3 ;
 ANTENNADIFFAREA                          0.160 LAYER ME4 ;
 ANTENNAMAXAREACAR                       21.782 LAYER ME2 ;
 ANTENNAMAXAREACAR                       24.449 LAYER ME3 ;
 ANTENNAMAXAREACAR                       27.116 LAYER ME4 ;
END DI84
PIN DO84
  DIRECTION OUTPUT ;
 PORT
  LAYER ME4 ;
  RECT 376.885 0.000 377.205 0.600 ;
  LAYER ME3 ;
  RECT 376.885 0.000 377.205 0.600 ;
  LAYER ME2 ;
  RECT 376.885 0.000 377.205 0.600 ;
  LAYER ME1 ;
  RECT 376.885 0.000 377.205 0.600 ;
 END
 ANTENNAPARTIALMETALAREA                  5.273 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME3 ;
 ANTENNADIFFAREA                          1.293 LAYER ME4 ;
END DO84
PIN DI83
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 373.443 0.000 373.763 0.600 ;
  LAYER ME3 ;
  RECT 373.443 0.000 373.763 0.600 ;
  LAYER ME2 ;
  RECT 373.443 0.000 373.763 0.600 ;
  LAYER ME1 ;
  RECT 373.443 0.000 373.763 0.600 ;
 END
 ANTENNAPARTIALMETALAREA                  1.058 LAYER ME2 ;
 ANTENNAGATEAREA                          0.072 LAYER ME2 ;
 ANTENNAGATEAREA                          0.072 LAYER ME3 ;
 ANTENNAGATEAREA                          0.072 LAYER ME4 ;
 ANTENNADIFFAREA                          0.160 LAYER ME2 ;
 ANTENNADIFFAREA                          0.160 LAYER ME3 ;
 ANTENNADIFFAREA                          0.160 LAYER ME4 ;
 ANTENNAMAXAREACAR                       21.782 LAYER ME2 ;
 ANTENNAMAXAREACAR                       24.449 LAYER ME3 ;
 ANTENNAMAXAREACAR                       27.116 LAYER ME4 ;
END DI83
PIN DO83
  DIRECTION OUTPUT ;
 PORT
  LAYER ME4 ;
  RECT 372.881 0.000 373.201 0.600 ;
  LAYER ME3 ;
  RECT 372.881 0.000 373.201 0.600 ;
  LAYER ME2 ;
  RECT 372.881 0.000 373.201 0.600 ;
  LAYER ME1 ;
  RECT 372.881 0.000 373.201 0.600 ;
 END
 ANTENNAPARTIALMETALAREA                  5.273 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME3 ;
 ANTENNADIFFAREA                          1.293 LAYER ME4 ;
END DO83
PIN DI82
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 369.439 0.000 369.759 0.600 ;
  LAYER ME3 ;
  RECT 369.439 0.000 369.759 0.600 ;
  LAYER ME2 ;
  RECT 369.439 0.000 369.759 0.600 ;
  LAYER ME1 ;
  RECT 369.439 0.000 369.759 0.600 ;
 END
 ANTENNAPARTIALMETALAREA                  1.058 LAYER ME2 ;
 ANTENNAGATEAREA                          0.072 LAYER ME2 ;
 ANTENNAGATEAREA                          0.072 LAYER ME3 ;
 ANTENNAGATEAREA                          0.072 LAYER ME4 ;
 ANTENNADIFFAREA                          0.160 LAYER ME2 ;
 ANTENNADIFFAREA                          0.160 LAYER ME3 ;
 ANTENNADIFFAREA                          0.160 LAYER ME4 ;
 ANTENNAMAXAREACAR                       21.782 LAYER ME2 ;
 ANTENNAMAXAREACAR                       24.449 LAYER ME3 ;
 ANTENNAMAXAREACAR                       27.116 LAYER ME4 ;
END DI82
PIN DO82
  DIRECTION OUTPUT ;
 PORT
  LAYER ME4 ;
  RECT 368.877 0.000 369.197 0.600 ;
  LAYER ME3 ;
  RECT 368.877 0.000 369.197 0.600 ;
  LAYER ME2 ;
  RECT 368.877 0.000 369.197 0.600 ;
  LAYER ME1 ;
  RECT 368.877 0.000 369.197 0.600 ;
 END
 ANTENNAPARTIALMETALAREA                  5.273 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME3 ;
 ANTENNADIFFAREA                          1.293 LAYER ME4 ;
END DO82
PIN DI81
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 365.435 0.000 365.755 0.600 ;
  LAYER ME3 ;
  RECT 365.435 0.000 365.755 0.600 ;
  LAYER ME2 ;
  RECT 365.435 0.000 365.755 0.600 ;
  LAYER ME1 ;
  RECT 365.435 0.000 365.755 0.600 ;
 END
 ANTENNAPARTIALMETALAREA                  1.058 LAYER ME2 ;
 ANTENNAGATEAREA                          0.072 LAYER ME2 ;
 ANTENNAGATEAREA                          0.072 LAYER ME3 ;
 ANTENNAGATEAREA                          0.072 LAYER ME4 ;
 ANTENNADIFFAREA                          0.160 LAYER ME2 ;
 ANTENNADIFFAREA                          0.160 LAYER ME3 ;
 ANTENNADIFFAREA                          0.160 LAYER ME4 ;
 ANTENNAMAXAREACAR                       21.782 LAYER ME2 ;
 ANTENNAMAXAREACAR                       24.449 LAYER ME3 ;
 ANTENNAMAXAREACAR                       27.116 LAYER ME4 ;
END DI81
PIN DO81
  DIRECTION OUTPUT ;
 PORT
  LAYER ME4 ;
  RECT 364.873 0.000 365.193 0.600 ;
  LAYER ME3 ;
  RECT 364.873 0.000 365.193 0.600 ;
  LAYER ME2 ;
  RECT 364.873 0.000 365.193 0.600 ;
  LAYER ME1 ;
  RECT 364.873 0.000 365.193 0.600 ;
 END
 ANTENNAPARTIALMETALAREA                  5.273 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME3 ;
 ANTENNADIFFAREA                          1.293 LAYER ME4 ;
END DO81
PIN DI80
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 360.869 0.000 361.189 0.600 ;
  LAYER ME3 ;
  RECT 360.869 0.000 361.189 0.600 ;
  LAYER ME2 ;
  RECT 360.869 0.000 361.189 0.600 ;
  LAYER ME1 ;
  RECT 360.869 0.000 361.189 0.600 ;
 END
 ANTENNAPARTIALMETALAREA                  0.346 LAYER ME1 ;
 ANTENNAPARTIALMETALAREA                  1.466 LAYER ME2 ;
 ANTENNAPARTIALMETALAREA                  0.508 LAYER ME3 ;
 ANTENNAGATEAREA                          0.072 LAYER ME3 ;
 ANTENNAGATEAREA                          0.072 LAYER ME4 ;
 ANTENNADIFFAREA                          0.218 LAYER ME1 ;
 ANTENNADIFFAREA                          0.218 LAYER ME2 ;
 ANTENNADIFFAREA                          0.218 LAYER ME3 ;
 ANTENNADIFFAREA                          0.218 LAYER ME4 ;
 ANTENNAMAXAREACAR                       17.267 LAYER ME3 ;
 ANTENNAMAXAREACAR                       19.933 LAYER ME4 ;
END DI80
PIN DO80
  DIRECTION OUTPUT ;
 PORT
  LAYER ME4 ;
  RECT 361.431 0.000 361.751 0.600 ;
  LAYER ME3 ;
  RECT 361.431 0.000 361.751 0.600 ;
  LAYER ME2 ;
  RECT 361.431 0.000 361.751 0.600 ;
  LAYER ME1 ;
  RECT 361.431 0.000 361.751 0.600 ;
 END
 ANTENNAPARTIALMETALAREA                  5.602 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME3 ;
 ANTENNADIFFAREA                          1.293 LAYER ME4 ;
END DO80
PIN WEB10
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 359.429 0.000 359.749 0.600 ;
  LAYER ME3 ;
  RECT 359.429 0.000 359.749 0.600 ;
  LAYER ME2 ;
  RECT 359.429 0.000 359.749 0.600 ;
  LAYER ME1 ;
  RECT 359.429 0.000 359.749 0.600 ;
 END
 ANTENNAPARTIALMETALAREA                  1.036 LAYER ME2 ;
 ANTENNAGATEAREA                          0.288 LAYER ME2 ;
 ANTENNAGATEAREA                          0.288 LAYER ME3 ;
 ANTENNAGATEAREA                          0.288 LAYER ME4 ;
 ANTENNADIFFAREA                          0.206 LAYER ME2 ;
 ANTENNADIFFAREA                          0.206 LAYER ME3 ;
 ANTENNADIFFAREA                          0.206 LAYER ME4 ;
 ANTENNAMAXAREACAR                        5.844 LAYER ME2 ;
 ANTENNAMAXAREACAR                        6.511 LAYER ME3 ;
 ANTENNAMAXAREACAR                        7.178 LAYER ME4 ;
END WEB10
PIN DI79
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 357.427 0.000 357.747 0.600 ;
  LAYER ME3 ;
  RECT 357.427 0.000 357.747 0.600 ;
  LAYER ME2 ;
  RECT 357.427 0.000 357.747 0.600 ;
  LAYER ME1 ;
  RECT 357.427 0.000 357.747 0.600 ;
 END
 ANTENNAPARTIALMETALAREA                  1.058 LAYER ME2 ;
 ANTENNAGATEAREA                          0.072 LAYER ME2 ;
 ANTENNAGATEAREA                          0.072 LAYER ME3 ;
 ANTENNAGATEAREA                          0.072 LAYER ME4 ;
 ANTENNADIFFAREA                          0.160 LAYER ME2 ;
 ANTENNADIFFAREA                          0.160 LAYER ME3 ;
 ANTENNADIFFAREA                          0.160 LAYER ME4 ;
 ANTENNAMAXAREACAR                       21.782 LAYER ME2 ;
 ANTENNAMAXAREACAR                       24.449 LAYER ME3 ;
 ANTENNAMAXAREACAR                       27.116 LAYER ME4 ;
END DI79
PIN DO79
  DIRECTION OUTPUT ;
 PORT
  LAYER ME4 ;
  RECT 356.865 0.000 357.185 0.600 ;
  LAYER ME3 ;
  RECT 356.865 0.000 357.185 0.600 ;
  LAYER ME2 ;
  RECT 356.865 0.000 357.185 0.600 ;
  LAYER ME1 ;
  RECT 356.865 0.000 357.185 0.600 ;
 END
 ANTENNAPARTIALMETALAREA                  5.273 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME3 ;
 ANTENNADIFFAREA                          1.293 LAYER ME4 ;
END DO79
PIN DI78
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 353.423 0.000 353.743 0.600 ;
  LAYER ME3 ;
  RECT 353.423 0.000 353.743 0.600 ;
  LAYER ME2 ;
  RECT 353.423 0.000 353.743 0.600 ;
  LAYER ME1 ;
  RECT 353.423 0.000 353.743 0.600 ;
 END
 ANTENNAPARTIALMETALAREA                  1.058 LAYER ME2 ;
 ANTENNAGATEAREA                          0.072 LAYER ME2 ;
 ANTENNAGATEAREA                          0.072 LAYER ME3 ;
 ANTENNAGATEAREA                          0.072 LAYER ME4 ;
 ANTENNADIFFAREA                          0.160 LAYER ME2 ;
 ANTENNADIFFAREA                          0.160 LAYER ME3 ;
 ANTENNADIFFAREA                          0.160 LAYER ME4 ;
 ANTENNAMAXAREACAR                       21.782 LAYER ME2 ;
 ANTENNAMAXAREACAR                       24.449 LAYER ME3 ;
 ANTENNAMAXAREACAR                       27.116 LAYER ME4 ;
END DI78
PIN DO78
  DIRECTION OUTPUT ;
 PORT
  LAYER ME4 ;
  RECT 352.861 0.000 353.181 0.600 ;
  LAYER ME3 ;
  RECT 352.861 0.000 353.181 0.600 ;
  LAYER ME2 ;
  RECT 352.861 0.000 353.181 0.600 ;
  LAYER ME1 ;
  RECT 352.861 0.000 353.181 0.600 ;
 END
 ANTENNAPARTIALMETALAREA                  5.273 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME3 ;
 ANTENNADIFFAREA                          1.293 LAYER ME4 ;
END DO78
PIN DI77
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 349.419 0.000 349.739 0.600 ;
  LAYER ME3 ;
  RECT 349.419 0.000 349.739 0.600 ;
  LAYER ME2 ;
  RECT 349.419 0.000 349.739 0.600 ;
  LAYER ME1 ;
  RECT 349.419 0.000 349.739 0.600 ;
 END
 ANTENNAPARTIALMETALAREA                  1.058 LAYER ME2 ;
 ANTENNAGATEAREA                          0.072 LAYER ME2 ;
 ANTENNAGATEAREA                          0.072 LAYER ME3 ;
 ANTENNAGATEAREA                          0.072 LAYER ME4 ;
 ANTENNADIFFAREA                          0.160 LAYER ME2 ;
 ANTENNADIFFAREA                          0.160 LAYER ME3 ;
 ANTENNADIFFAREA                          0.160 LAYER ME4 ;
 ANTENNAMAXAREACAR                       21.782 LAYER ME2 ;
 ANTENNAMAXAREACAR                       24.449 LAYER ME3 ;
 ANTENNAMAXAREACAR                       27.116 LAYER ME4 ;
END DI77
PIN DO77
  DIRECTION OUTPUT ;
 PORT
  LAYER ME4 ;
  RECT 348.857 0.000 349.177 0.600 ;
  LAYER ME3 ;
  RECT 348.857 0.000 349.177 0.600 ;
  LAYER ME2 ;
  RECT 348.857 0.000 349.177 0.600 ;
  LAYER ME1 ;
  RECT 348.857 0.000 349.177 0.600 ;
 END
 ANTENNAPARTIALMETALAREA                  5.273 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME3 ;
 ANTENNADIFFAREA                          1.293 LAYER ME4 ;
END DO77
PIN DI76
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 345.415 0.000 345.735 0.600 ;
  LAYER ME3 ;
  RECT 345.415 0.000 345.735 0.600 ;
  LAYER ME2 ;
  RECT 345.415 0.000 345.735 0.600 ;
  LAYER ME1 ;
  RECT 345.415 0.000 345.735 0.600 ;
 END
 ANTENNAPARTIALMETALAREA                  1.058 LAYER ME2 ;
 ANTENNAGATEAREA                          0.072 LAYER ME2 ;
 ANTENNAGATEAREA                          0.072 LAYER ME3 ;
 ANTENNAGATEAREA                          0.072 LAYER ME4 ;
 ANTENNADIFFAREA                          0.160 LAYER ME2 ;
 ANTENNADIFFAREA                          0.160 LAYER ME3 ;
 ANTENNADIFFAREA                          0.160 LAYER ME4 ;
 ANTENNAMAXAREACAR                       21.782 LAYER ME2 ;
 ANTENNAMAXAREACAR                       24.449 LAYER ME3 ;
 ANTENNAMAXAREACAR                       27.116 LAYER ME4 ;
END DI76
PIN DO76
  DIRECTION OUTPUT ;
 PORT
  LAYER ME4 ;
  RECT 344.853 0.000 345.173 0.600 ;
  LAYER ME3 ;
  RECT 344.853 0.000 345.173 0.600 ;
  LAYER ME2 ;
  RECT 344.853 0.000 345.173 0.600 ;
  LAYER ME1 ;
  RECT 344.853 0.000 345.173 0.600 ;
 END
 ANTENNAPARTIALMETALAREA                  5.273 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME3 ;
 ANTENNADIFFAREA                          1.293 LAYER ME4 ;
END DO76
PIN DI75
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 341.411 0.000 341.731 0.600 ;
  LAYER ME3 ;
  RECT 341.411 0.000 341.731 0.600 ;
  LAYER ME2 ;
  RECT 341.411 0.000 341.731 0.600 ;
  LAYER ME1 ;
  RECT 341.411 0.000 341.731 0.600 ;
 END
 ANTENNAPARTIALMETALAREA                  1.058 LAYER ME2 ;
 ANTENNAGATEAREA                          0.072 LAYER ME2 ;
 ANTENNAGATEAREA                          0.072 LAYER ME3 ;
 ANTENNAGATEAREA                          0.072 LAYER ME4 ;
 ANTENNADIFFAREA                          0.160 LAYER ME2 ;
 ANTENNADIFFAREA                          0.160 LAYER ME3 ;
 ANTENNADIFFAREA                          0.160 LAYER ME4 ;
 ANTENNAMAXAREACAR                       21.782 LAYER ME2 ;
 ANTENNAMAXAREACAR                       24.449 LAYER ME3 ;
 ANTENNAMAXAREACAR                       27.116 LAYER ME4 ;
END DI75
PIN DO75
  DIRECTION OUTPUT ;
 PORT
  LAYER ME4 ;
  RECT 340.849 0.000 341.169 0.600 ;
  LAYER ME3 ;
  RECT 340.849 0.000 341.169 0.600 ;
  LAYER ME2 ;
  RECT 340.849 0.000 341.169 0.600 ;
  LAYER ME1 ;
  RECT 340.849 0.000 341.169 0.600 ;
 END
 ANTENNAPARTIALMETALAREA                  5.273 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME3 ;
 ANTENNADIFFAREA                          1.293 LAYER ME4 ;
END DO75
PIN DI74
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 337.407 0.000 337.727 0.600 ;
  LAYER ME3 ;
  RECT 337.407 0.000 337.727 0.600 ;
  LAYER ME2 ;
  RECT 337.407 0.000 337.727 0.600 ;
  LAYER ME1 ;
  RECT 337.407 0.000 337.727 0.600 ;
 END
 ANTENNAPARTIALMETALAREA                  1.058 LAYER ME2 ;
 ANTENNAGATEAREA                          0.072 LAYER ME2 ;
 ANTENNAGATEAREA                          0.072 LAYER ME3 ;
 ANTENNAGATEAREA                          0.072 LAYER ME4 ;
 ANTENNADIFFAREA                          0.160 LAYER ME2 ;
 ANTENNADIFFAREA                          0.160 LAYER ME3 ;
 ANTENNADIFFAREA                          0.160 LAYER ME4 ;
 ANTENNAMAXAREACAR                       21.782 LAYER ME2 ;
 ANTENNAMAXAREACAR                       24.449 LAYER ME3 ;
 ANTENNAMAXAREACAR                       27.116 LAYER ME4 ;
END DI74
PIN DO74
  DIRECTION OUTPUT ;
 PORT
  LAYER ME4 ;
  RECT 336.845 0.000 337.165 0.600 ;
  LAYER ME3 ;
  RECT 336.845 0.000 337.165 0.600 ;
  LAYER ME2 ;
  RECT 336.845 0.000 337.165 0.600 ;
  LAYER ME1 ;
  RECT 336.845 0.000 337.165 0.600 ;
 END
 ANTENNAPARTIALMETALAREA                  5.273 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME3 ;
 ANTENNADIFFAREA                          1.293 LAYER ME4 ;
END DO74
PIN DI73
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 333.403 0.000 333.723 0.600 ;
  LAYER ME3 ;
  RECT 333.403 0.000 333.723 0.600 ;
  LAYER ME2 ;
  RECT 333.403 0.000 333.723 0.600 ;
  LAYER ME1 ;
  RECT 333.403 0.000 333.723 0.600 ;
 END
 ANTENNAPARTIALMETALAREA                  1.058 LAYER ME2 ;
 ANTENNAGATEAREA                          0.072 LAYER ME2 ;
 ANTENNAGATEAREA                          0.072 LAYER ME3 ;
 ANTENNAGATEAREA                          0.072 LAYER ME4 ;
 ANTENNADIFFAREA                          0.160 LAYER ME2 ;
 ANTENNADIFFAREA                          0.160 LAYER ME3 ;
 ANTENNADIFFAREA                          0.160 LAYER ME4 ;
 ANTENNAMAXAREACAR                       21.782 LAYER ME2 ;
 ANTENNAMAXAREACAR                       24.449 LAYER ME3 ;
 ANTENNAMAXAREACAR                       27.116 LAYER ME4 ;
END DI73
PIN DO73
  DIRECTION OUTPUT ;
 PORT
  LAYER ME4 ;
  RECT 332.841 0.000 333.161 0.600 ;
  LAYER ME3 ;
  RECT 332.841 0.000 333.161 0.600 ;
  LAYER ME2 ;
  RECT 332.841 0.000 333.161 0.600 ;
  LAYER ME1 ;
  RECT 332.841 0.000 333.161 0.600 ;
 END
 ANTENNAPARTIALMETALAREA                  5.273 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME3 ;
 ANTENNADIFFAREA                          1.293 LAYER ME4 ;
END DO73
PIN DI72
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 328.837 0.000 329.157 0.600 ;
  LAYER ME3 ;
  RECT 328.837 0.000 329.157 0.600 ;
  LAYER ME2 ;
  RECT 328.837 0.000 329.157 0.600 ;
  LAYER ME1 ;
  RECT 328.837 0.000 329.157 0.600 ;
 END
 ANTENNAPARTIALMETALAREA                  0.346 LAYER ME1 ;
 ANTENNAPARTIALMETALAREA                  1.466 LAYER ME2 ;
 ANTENNAPARTIALMETALAREA                  0.508 LAYER ME3 ;
 ANTENNAGATEAREA                          0.072 LAYER ME3 ;
 ANTENNAGATEAREA                          0.072 LAYER ME4 ;
 ANTENNADIFFAREA                          0.218 LAYER ME1 ;
 ANTENNADIFFAREA                          0.218 LAYER ME2 ;
 ANTENNADIFFAREA                          0.218 LAYER ME3 ;
 ANTENNADIFFAREA                          0.218 LAYER ME4 ;
 ANTENNAMAXAREACAR                       17.267 LAYER ME3 ;
 ANTENNAMAXAREACAR                       19.933 LAYER ME4 ;
END DI72
PIN DO72
  DIRECTION OUTPUT ;
 PORT
  LAYER ME4 ;
  RECT 329.399 0.000 329.719 0.600 ;
  LAYER ME3 ;
  RECT 329.399 0.000 329.719 0.600 ;
  LAYER ME2 ;
  RECT 329.399 0.000 329.719 0.600 ;
  LAYER ME1 ;
  RECT 329.399 0.000 329.719 0.600 ;
 END
 ANTENNAPARTIALMETALAREA                  5.602 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME3 ;
 ANTENNADIFFAREA                          1.293 LAYER ME4 ;
END DO72
PIN WEB9
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 327.397 0.000 327.717 0.600 ;
  LAYER ME3 ;
  RECT 327.397 0.000 327.717 0.600 ;
  LAYER ME2 ;
  RECT 327.397 0.000 327.717 0.600 ;
  LAYER ME1 ;
  RECT 327.397 0.000 327.717 0.600 ;
 END
 ANTENNAPARTIALMETALAREA                  1.036 LAYER ME2 ;
 ANTENNAGATEAREA                          0.288 LAYER ME2 ;
 ANTENNAGATEAREA                          0.288 LAYER ME3 ;
 ANTENNAGATEAREA                          0.288 LAYER ME4 ;
 ANTENNADIFFAREA                          0.206 LAYER ME2 ;
 ANTENNADIFFAREA                          0.206 LAYER ME3 ;
 ANTENNADIFFAREA                          0.206 LAYER ME4 ;
 ANTENNAMAXAREACAR                        5.844 LAYER ME2 ;
 ANTENNAMAXAREACAR                        6.511 LAYER ME3 ;
 ANTENNAMAXAREACAR                        7.178 LAYER ME4 ;
END WEB9
PIN DI71
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 325.395 0.000 325.715 0.600 ;
  LAYER ME3 ;
  RECT 325.395 0.000 325.715 0.600 ;
  LAYER ME2 ;
  RECT 325.395 0.000 325.715 0.600 ;
  LAYER ME1 ;
  RECT 325.395 0.000 325.715 0.600 ;
 END
 ANTENNAPARTIALMETALAREA                  1.058 LAYER ME2 ;
 ANTENNAGATEAREA                          0.072 LAYER ME2 ;
 ANTENNAGATEAREA                          0.072 LAYER ME3 ;
 ANTENNAGATEAREA                          0.072 LAYER ME4 ;
 ANTENNADIFFAREA                          0.160 LAYER ME2 ;
 ANTENNADIFFAREA                          0.160 LAYER ME3 ;
 ANTENNADIFFAREA                          0.160 LAYER ME4 ;
 ANTENNAMAXAREACAR                       21.782 LAYER ME2 ;
 ANTENNAMAXAREACAR                       24.449 LAYER ME3 ;
 ANTENNAMAXAREACAR                       27.116 LAYER ME4 ;
END DI71
PIN DO71
  DIRECTION OUTPUT ;
 PORT
  LAYER ME4 ;
  RECT 324.833 0.000 325.153 0.600 ;
  LAYER ME3 ;
  RECT 324.833 0.000 325.153 0.600 ;
  LAYER ME2 ;
  RECT 324.833 0.000 325.153 0.600 ;
  LAYER ME1 ;
  RECT 324.833 0.000 325.153 0.600 ;
 END
 ANTENNAPARTIALMETALAREA                  5.273 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME3 ;
 ANTENNADIFFAREA                          1.293 LAYER ME4 ;
END DO71
PIN DI70
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 321.391 0.000 321.711 0.600 ;
  LAYER ME3 ;
  RECT 321.391 0.000 321.711 0.600 ;
  LAYER ME2 ;
  RECT 321.391 0.000 321.711 0.600 ;
  LAYER ME1 ;
  RECT 321.391 0.000 321.711 0.600 ;
 END
 ANTENNAPARTIALMETALAREA                  1.058 LAYER ME2 ;
 ANTENNAGATEAREA                          0.072 LAYER ME2 ;
 ANTENNAGATEAREA                          0.072 LAYER ME3 ;
 ANTENNAGATEAREA                          0.072 LAYER ME4 ;
 ANTENNADIFFAREA                          0.160 LAYER ME2 ;
 ANTENNADIFFAREA                          0.160 LAYER ME3 ;
 ANTENNADIFFAREA                          0.160 LAYER ME4 ;
 ANTENNAMAXAREACAR                       21.782 LAYER ME2 ;
 ANTENNAMAXAREACAR                       24.449 LAYER ME3 ;
 ANTENNAMAXAREACAR                       27.116 LAYER ME4 ;
END DI70
PIN DO70
  DIRECTION OUTPUT ;
 PORT
  LAYER ME4 ;
  RECT 320.829 0.000 321.149 0.600 ;
  LAYER ME3 ;
  RECT 320.829 0.000 321.149 0.600 ;
  LAYER ME2 ;
  RECT 320.829 0.000 321.149 0.600 ;
  LAYER ME1 ;
  RECT 320.829 0.000 321.149 0.600 ;
 END
 ANTENNAPARTIALMETALAREA                  5.273 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME3 ;
 ANTENNADIFFAREA                          1.293 LAYER ME4 ;
END DO70
PIN DI69
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 317.387 0.000 317.707 0.600 ;
  LAYER ME3 ;
  RECT 317.387 0.000 317.707 0.600 ;
  LAYER ME2 ;
  RECT 317.387 0.000 317.707 0.600 ;
  LAYER ME1 ;
  RECT 317.387 0.000 317.707 0.600 ;
 END
 ANTENNAPARTIALMETALAREA                  1.058 LAYER ME2 ;
 ANTENNAGATEAREA                          0.072 LAYER ME2 ;
 ANTENNAGATEAREA                          0.072 LAYER ME3 ;
 ANTENNAGATEAREA                          0.072 LAYER ME4 ;
 ANTENNADIFFAREA                          0.160 LAYER ME2 ;
 ANTENNADIFFAREA                          0.160 LAYER ME3 ;
 ANTENNADIFFAREA                          0.160 LAYER ME4 ;
 ANTENNAMAXAREACAR                       21.782 LAYER ME2 ;
 ANTENNAMAXAREACAR                       24.449 LAYER ME3 ;
 ANTENNAMAXAREACAR                       27.116 LAYER ME4 ;
END DI69
PIN DO69
  DIRECTION OUTPUT ;
 PORT
  LAYER ME4 ;
  RECT 316.825 0.000 317.145 0.600 ;
  LAYER ME3 ;
  RECT 316.825 0.000 317.145 0.600 ;
  LAYER ME2 ;
  RECT 316.825 0.000 317.145 0.600 ;
  LAYER ME1 ;
  RECT 316.825 0.000 317.145 0.600 ;
 END
 ANTENNAPARTIALMETALAREA                  5.273 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME3 ;
 ANTENNADIFFAREA                          1.293 LAYER ME4 ;
END DO69
PIN DI68
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 313.383 0.000 313.703 0.600 ;
  LAYER ME3 ;
  RECT 313.383 0.000 313.703 0.600 ;
  LAYER ME2 ;
  RECT 313.383 0.000 313.703 0.600 ;
  LAYER ME1 ;
  RECT 313.383 0.000 313.703 0.600 ;
 END
 ANTENNAPARTIALMETALAREA                  1.058 LAYER ME2 ;
 ANTENNAGATEAREA                          0.072 LAYER ME2 ;
 ANTENNAGATEAREA                          0.072 LAYER ME3 ;
 ANTENNAGATEAREA                          0.072 LAYER ME4 ;
 ANTENNADIFFAREA                          0.160 LAYER ME2 ;
 ANTENNADIFFAREA                          0.160 LAYER ME3 ;
 ANTENNADIFFAREA                          0.160 LAYER ME4 ;
 ANTENNAMAXAREACAR                       21.782 LAYER ME2 ;
 ANTENNAMAXAREACAR                       24.449 LAYER ME3 ;
 ANTENNAMAXAREACAR                       27.116 LAYER ME4 ;
END DI68
PIN DO68
  DIRECTION OUTPUT ;
 PORT
  LAYER ME4 ;
  RECT 312.821 0.000 313.141 0.600 ;
  LAYER ME3 ;
  RECT 312.821 0.000 313.141 0.600 ;
  LAYER ME2 ;
  RECT 312.821 0.000 313.141 0.600 ;
  LAYER ME1 ;
  RECT 312.821 0.000 313.141 0.600 ;
 END
 ANTENNAPARTIALMETALAREA                  5.273 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME3 ;
 ANTENNADIFFAREA                          1.293 LAYER ME4 ;
END DO68
PIN DI67
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 309.379 0.000 309.699 0.600 ;
  LAYER ME3 ;
  RECT 309.379 0.000 309.699 0.600 ;
  LAYER ME2 ;
  RECT 309.379 0.000 309.699 0.600 ;
  LAYER ME1 ;
  RECT 309.379 0.000 309.699 0.600 ;
 END
 ANTENNAPARTIALMETALAREA                  1.058 LAYER ME2 ;
 ANTENNAGATEAREA                          0.072 LAYER ME2 ;
 ANTENNAGATEAREA                          0.072 LAYER ME3 ;
 ANTENNAGATEAREA                          0.072 LAYER ME4 ;
 ANTENNADIFFAREA                          0.160 LAYER ME2 ;
 ANTENNADIFFAREA                          0.160 LAYER ME3 ;
 ANTENNADIFFAREA                          0.160 LAYER ME4 ;
 ANTENNAMAXAREACAR                       21.782 LAYER ME2 ;
 ANTENNAMAXAREACAR                       24.449 LAYER ME3 ;
 ANTENNAMAXAREACAR                       27.116 LAYER ME4 ;
END DI67
PIN DO67
  DIRECTION OUTPUT ;
 PORT
  LAYER ME4 ;
  RECT 308.817 0.000 309.137 0.600 ;
  LAYER ME3 ;
  RECT 308.817 0.000 309.137 0.600 ;
  LAYER ME2 ;
  RECT 308.817 0.000 309.137 0.600 ;
  LAYER ME1 ;
  RECT 308.817 0.000 309.137 0.600 ;
 END
 ANTENNAPARTIALMETALAREA                  5.273 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME3 ;
 ANTENNADIFFAREA                          1.293 LAYER ME4 ;
END DO67
PIN DI66
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 305.375 0.000 305.695 0.600 ;
  LAYER ME3 ;
  RECT 305.375 0.000 305.695 0.600 ;
  LAYER ME2 ;
  RECT 305.375 0.000 305.695 0.600 ;
  LAYER ME1 ;
  RECT 305.375 0.000 305.695 0.600 ;
 END
 ANTENNAPARTIALMETALAREA                  1.058 LAYER ME2 ;
 ANTENNAGATEAREA                          0.072 LAYER ME2 ;
 ANTENNAGATEAREA                          0.072 LAYER ME3 ;
 ANTENNAGATEAREA                          0.072 LAYER ME4 ;
 ANTENNADIFFAREA                          0.160 LAYER ME2 ;
 ANTENNADIFFAREA                          0.160 LAYER ME3 ;
 ANTENNADIFFAREA                          0.160 LAYER ME4 ;
 ANTENNAMAXAREACAR                       21.782 LAYER ME2 ;
 ANTENNAMAXAREACAR                       24.449 LAYER ME3 ;
 ANTENNAMAXAREACAR                       27.116 LAYER ME4 ;
END DI66
PIN DO66
  DIRECTION OUTPUT ;
 PORT
  LAYER ME4 ;
  RECT 304.813 0.000 305.133 0.600 ;
  LAYER ME3 ;
  RECT 304.813 0.000 305.133 0.600 ;
  LAYER ME2 ;
  RECT 304.813 0.000 305.133 0.600 ;
  LAYER ME1 ;
  RECT 304.813 0.000 305.133 0.600 ;
 END
 ANTENNAPARTIALMETALAREA                  5.273 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME3 ;
 ANTENNADIFFAREA                          1.293 LAYER ME4 ;
END DO66
PIN DI65
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 301.371 0.000 301.691 0.600 ;
  LAYER ME3 ;
  RECT 301.371 0.000 301.691 0.600 ;
  LAYER ME2 ;
  RECT 301.371 0.000 301.691 0.600 ;
  LAYER ME1 ;
  RECT 301.371 0.000 301.691 0.600 ;
 END
 ANTENNAPARTIALMETALAREA                  1.058 LAYER ME2 ;
 ANTENNAGATEAREA                          0.072 LAYER ME2 ;
 ANTENNAGATEAREA                          0.072 LAYER ME3 ;
 ANTENNAGATEAREA                          0.072 LAYER ME4 ;
 ANTENNADIFFAREA                          0.160 LAYER ME2 ;
 ANTENNADIFFAREA                          0.160 LAYER ME3 ;
 ANTENNADIFFAREA                          0.160 LAYER ME4 ;
 ANTENNAMAXAREACAR                       21.782 LAYER ME2 ;
 ANTENNAMAXAREACAR                       24.449 LAYER ME3 ;
 ANTENNAMAXAREACAR                       27.116 LAYER ME4 ;
END DI65
PIN DO65
  DIRECTION OUTPUT ;
 PORT
  LAYER ME4 ;
  RECT 300.809 0.000 301.129 0.600 ;
  LAYER ME3 ;
  RECT 300.809 0.000 301.129 0.600 ;
  LAYER ME2 ;
  RECT 300.809 0.000 301.129 0.600 ;
  LAYER ME1 ;
  RECT 300.809 0.000 301.129 0.600 ;
 END
 ANTENNAPARTIALMETALAREA                  5.273 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME3 ;
 ANTENNADIFFAREA                          1.293 LAYER ME4 ;
END DO65
PIN DI64
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 296.805 0.000 297.125 0.600 ;
  LAYER ME3 ;
  RECT 296.805 0.000 297.125 0.600 ;
  LAYER ME2 ;
  RECT 296.805 0.000 297.125 0.600 ;
  LAYER ME1 ;
  RECT 296.805 0.000 297.125 0.600 ;
 END
 ANTENNAPARTIALMETALAREA                  0.346 LAYER ME1 ;
 ANTENNAPARTIALMETALAREA                  1.466 LAYER ME2 ;
 ANTENNAPARTIALMETALAREA                  0.508 LAYER ME3 ;
 ANTENNAGATEAREA                          0.072 LAYER ME3 ;
 ANTENNAGATEAREA                          0.072 LAYER ME4 ;
 ANTENNADIFFAREA                          0.218 LAYER ME1 ;
 ANTENNADIFFAREA                          0.218 LAYER ME2 ;
 ANTENNADIFFAREA                          0.218 LAYER ME3 ;
 ANTENNADIFFAREA                          0.218 LAYER ME4 ;
 ANTENNAMAXAREACAR                       17.267 LAYER ME3 ;
 ANTENNAMAXAREACAR                       19.933 LAYER ME4 ;
END DI64
PIN DO64
  DIRECTION OUTPUT ;
 PORT
  LAYER ME4 ;
  RECT 297.367 0.000 297.687 0.600 ;
  LAYER ME3 ;
  RECT 297.367 0.000 297.687 0.600 ;
  LAYER ME2 ;
  RECT 297.367 0.000 297.687 0.600 ;
  LAYER ME1 ;
  RECT 297.367 0.000 297.687 0.600 ;
 END
 ANTENNAPARTIALMETALAREA                  5.602 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME3 ;
 ANTENNADIFFAREA                          1.293 LAYER ME4 ;
END DO64
PIN WEB8
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 295.365 0.000 295.685 0.600 ;
  LAYER ME3 ;
  RECT 295.365 0.000 295.685 0.600 ;
  LAYER ME2 ;
  RECT 295.365 0.000 295.685 0.600 ;
  LAYER ME1 ;
  RECT 295.365 0.000 295.685 0.600 ;
 END
 ANTENNAPARTIALMETALAREA                  1.036 LAYER ME2 ;
 ANTENNAGATEAREA                          0.288 LAYER ME2 ;
 ANTENNAGATEAREA                          0.288 LAYER ME3 ;
 ANTENNAGATEAREA                          0.288 LAYER ME4 ;
 ANTENNADIFFAREA                          0.206 LAYER ME2 ;
 ANTENNADIFFAREA                          0.206 LAYER ME3 ;
 ANTENNADIFFAREA                          0.206 LAYER ME4 ;
 ANTENNAMAXAREACAR                        5.844 LAYER ME2 ;
 ANTENNAMAXAREACAR                        6.511 LAYER ME3 ;
 ANTENNAMAXAREACAR                        7.178 LAYER ME4 ;
END WEB8
OBS
  LAYER ME3 SPACING 0.260 ;
  RECT 0.000 0.000 554.411 66.831 ;
  LAYER ME2 SPACING 0.260 ;
  RECT 0.000 0.000 554.411 66.831 ;
  LAYER ME1 SPACING 0.260 ;
  RECT 0.000 0.000 554.411 66.831 ;
  LAYER ME4 SPACING 0.260 ;
  RECT 0.000 0.000 270.398 66.831 ;
  LAYER ME4 SPACING 0.260 ;
  RECT 272.052 0.000 273.172 66.831 ;
  LAYER ME4 SPACING 0.260 ;
  RECT 274.767 0.000 275.487 66.831 ;
  LAYER ME4 SPACING 0.260 ;
  RECT 276.217 0.000 276.937 66.831 ;
  LAYER ME4 SPACING 0.260 ;
  RECT 278.997 0.000 279.597 66.831 ;
  LAYER ME4 SPACING 0.260 ;
  RECT 282.211 0.000 283.897 66.831 ;
  LAYER ME4 SPACING 0.260 ;
  RECT 285.287 0.000 286.407 66.831 ;
  LAYER ME4 SPACING 0.260 ;
  RECT 287.682 0.000 288.402 66.831 ;
  LAYER ME4 SPACING 0.260 ;
  RECT 289.397 0.000 290.117 66.831 ;
  LAYER ME4 SPACING 0.260 ;
  RECT 291.317 0.000 554.411 66.831 ;
END
END SYKB110_32X8X16CM2
END LIBRARY





