# ________________________________________________________________________________________________
# 
# 
#             Synchronous One-Port Register File Compiler
# 
#                 UMC 0.11um LL AE Logic Process
# 
# ________________________________________________________________________________________________
# 
#               
#         Copyright (C) 2024 Faraday Technology Corporation. All Rights Reserved.       
#                
#         This source code is an unpublished work belongs to Faraday Technology Corporation       
#         It is considered a trade secret and is not to be divulged or       
#         used by parties who have not received written authorization from       
#         Faraday Technology Corporation       
#                
#         Faraday's home page can be found at: http://www.faraday-tech.com/       
#                
# ________________________________________________________________________________________________
# 
#        IP Name            :  FSR0K_B_SY                
#        IP Version         :  1.4.0                     
#        IP Release Status  :  Active                    
#        Word               :  32                        
#        Bit                :  11                        
#        Byte               :  8                         
#        Mux                :  2                         
#        Output Loading     :  0.01                      
#        Clock Input Slew   :  0.016                     
#        Data Input Slew    :  0.016                     
#        Ring Type          :  Ringless Model            
#        Ring Width         :  0                         
#        Bus Format         :  0                         
#        Memaker Path       :  /home/mem/Desktop/memlib  
#        GUI Version        :  m20230904                 
#        Date               :  2024/09/06 20:28:37       
# ________________________________________________________________________________________________
# 

VERSION 5.5 ;
NAMESCASESENSITIVE ON ;
MACRO SYKB110_32X11X8CM2
CLASS BLOCK ;
FOREIGN SYKB110_32X11X8CM2 0.000 0.000 ;
ORIGIN 0.000 0.000 ;
SIZE 394.251 BY 66.831 ;
SYMMETRY x y r90 ;
SITE core ;
PIN GND
  DIRECTION INOUT ;
  USE GROUND ;
 PORT
  LAYER ME4 ;
  RECT 218.998 1.781 219.338 66.831 ;
 END
 PORT
  LAYER ME4 ;
  RECT 214.994 1.781 215.334 66.831 ;
 END
 PORT
  LAYER ME4 ;
  RECT 216.996 1.781 217.336 66.831 ;
 END
 PORT
  LAYER ME4 ;
  RECT 217.807 0.000 218.527 44.094 ;
 END
 PORT
  LAYER ME4 ;
  RECT 223.002 1.781 223.342 66.831 ;
 END
 PORT
  LAYER ME4 ;
  RECT 221.000 1.781 221.340 66.831 ;
 END
 PORT
  LAYER ME4 ;
  RECT 221.811 0.000 222.531 44.094 ;
 END
 PORT
  LAYER ME4 ;
  RECT 227.006 1.781 227.346 66.831 ;
 END
 PORT
  LAYER ME4 ;
  RECT 225.004 1.781 225.344 66.831 ;
 END
 PORT
  LAYER ME4 ;
  RECT 225.815 0.000 226.535 44.094 ;
 END
 PORT
  LAYER ME4 ;
  RECT 231.010 1.781 231.350 66.831 ;
 END
 PORT
  LAYER ME4 ;
  RECT 229.008 1.781 229.348 66.831 ;
 END
 PORT
  LAYER ME4 ;
  RECT 229.819 0.000 230.539 44.094 ;
 END
 PORT
  LAYER ME4 ;
  RECT 235.014 1.781 235.354 66.831 ;
 END
 PORT
  LAYER ME4 ;
  RECT 233.012 1.781 233.352 66.831 ;
 END
 PORT
  LAYER ME4 ;
  RECT 233.823 0.000 234.543 44.094 ;
 END
 PORT
  LAYER ME4 ;
  RECT 239.018 1.781 239.358 66.831 ;
 END
 PORT
  LAYER ME4 ;
  RECT 237.016 1.781 237.356 66.831 ;
 END
 PORT
  LAYER ME4 ;
  RECT 237.827 0.000 238.547 44.094 ;
 END
 PORT
  LAYER ME4 ;
  RECT 243.022 1.781 243.362 66.831 ;
 END
 PORT
  LAYER ME4 ;
  RECT 241.020 1.781 241.360 66.831 ;
 END
 PORT
  LAYER ME4 ;
  RECT 241.831 0.000 242.551 44.094 ;
 END
 PORT
  LAYER ME4 ;
  RECT 247.026 1.781 247.366 66.831 ;
 END
 PORT
  LAYER ME4 ;
  RECT 245.024 1.781 245.364 66.831 ;
 END
 PORT
  LAYER ME4 ;
  RECT 245.835 0.000 246.555 44.094 ;
 END
 PORT
  LAYER ME4 ;
  RECT 251.030 1.781 251.370 66.831 ;
 END
 PORT
  LAYER ME4 ;
  RECT 249.028 1.781 249.368 66.831 ;
 END
 PORT
  LAYER ME4 ;
  RECT 249.839 0.000 250.559 44.094 ;
 END
 PORT
  LAYER ME4 ;
  RECT 255.034 1.781 255.374 66.831 ;
 END
 PORT
  LAYER ME4 ;
  RECT 253.032 1.781 253.372 66.831 ;
 END
 PORT
  LAYER ME4 ;
  RECT 253.843 0.000 254.563 44.094 ;
 END
 PORT
  LAYER ME4 ;
  RECT 259.038 1.781 259.378 66.831 ;
 END
 PORT
  LAYER ME4 ;
  RECT 257.036 1.781 257.376 66.831 ;
 END
 PORT
  LAYER ME4 ;
  RECT 257.847 0.000 258.567 44.094 ;
 END
 PORT
  LAYER ME4 ;
  RECT 263.042 1.781 263.382 66.831 ;
 END
 PORT
  LAYER ME4 ;
  RECT 261.040 1.781 261.380 66.831 ;
 END
 PORT
  LAYER ME4 ;
  RECT 261.851 0.000 262.571 44.094 ;
 END
 PORT
  LAYER ME4 ;
  RECT 267.046 1.781 267.386 66.831 ;
 END
 PORT
  LAYER ME4 ;
  RECT 265.044 1.781 265.384 66.831 ;
 END
 PORT
  LAYER ME4 ;
  RECT 265.855 0.000 266.575 44.094 ;
 END
 PORT
  LAYER ME4 ;
  RECT 271.050 1.781 271.390 66.831 ;
 END
 PORT
  LAYER ME4 ;
  RECT 269.048 1.781 269.388 66.831 ;
 END
 PORT
  LAYER ME4 ;
  RECT 269.859 0.000 270.579 44.094 ;
 END
 PORT
  LAYER ME4 ;
  RECT 275.054 1.781 275.394 66.831 ;
 END
 PORT
  LAYER ME4 ;
  RECT 273.052 1.781 273.392 66.831 ;
 END
 PORT
  LAYER ME4 ;
  RECT 273.863 0.000 274.583 44.094 ;
 END
 PORT
  LAYER ME4 ;
  RECT 279.058 1.781 279.398 66.831 ;
 END
 PORT
  LAYER ME4 ;
  RECT 277.056 1.781 277.396 66.831 ;
 END
 PORT
  LAYER ME4 ;
  RECT 277.867 0.000 278.587 44.094 ;
 END
 PORT
  LAYER ME4 ;
  RECT 283.062 1.781 283.402 66.831 ;
 END
 PORT
  LAYER ME4 ;
  RECT 281.060 1.781 281.400 66.831 ;
 END
 PORT
  LAYER ME4 ;
  RECT 281.871 0.000 282.591 44.094 ;
 END
 PORT
  LAYER ME4 ;
  RECT 287.066 1.781 287.406 66.831 ;
 END
 PORT
  LAYER ME4 ;
  RECT 285.064 1.781 285.404 66.831 ;
 END
 PORT
  LAYER ME4 ;
  RECT 285.875 0.000 286.595 44.094 ;
 END
 PORT
  LAYER ME4 ;
  RECT 291.070 1.781 291.410 66.831 ;
 END
 PORT
  LAYER ME4 ;
  RECT 289.068 1.781 289.408 66.831 ;
 END
 PORT
  LAYER ME4 ;
  RECT 289.879 0.000 290.599 44.094 ;
 END
 PORT
  LAYER ME4 ;
  RECT 295.074 1.781 295.414 66.831 ;
 END
 PORT
  LAYER ME4 ;
  RECT 293.072 1.781 293.412 66.831 ;
 END
 PORT
  LAYER ME4 ;
  RECT 293.883 0.000 294.603 44.094 ;
 END
 PORT
  LAYER ME4 ;
  RECT 299.078 1.781 299.418 66.831 ;
 END
 PORT
  LAYER ME4 ;
  RECT 297.076 1.781 297.416 66.831 ;
 END
 PORT
  LAYER ME4 ;
  RECT 297.887 0.000 298.607 44.094 ;
 END
 PORT
  LAYER ME4 ;
  RECT 303.082 1.781 303.422 66.831 ;
 END
 PORT
  LAYER ME4 ;
  RECT 301.080 1.781 301.420 66.831 ;
 END
 PORT
  LAYER ME4 ;
  RECT 301.891 0.000 302.611 44.094 ;
 END
 PORT
  LAYER ME4 ;
  RECT 307.086 1.781 307.426 66.831 ;
 END
 PORT
  LAYER ME4 ;
  RECT 305.084 1.781 305.424 66.831 ;
 END
 PORT
  LAYER ME4 ;
  RECT 305.895 0.000 306.615 44.094 ;
 END
 PORT
  LAYER ME4 ;
  RECT 311.090 1.781 311.430 66.831 ;
 END
 PORT
  LAYER ME4 ;
  RECT 309.088 1.781 309.428 66.831 ;
 END
 PORT
  LAYER ME4 ;
  RECT 309.899 0.000 310.619 44.094 ;
 END
 PORT
  LAYER ME4 ;
  RECT 315.094 1.781 315.434 66.831 ;
 END
 PORT
  LAYER ME4 ;
  RECT 313.092 1.781 313.432 66.831 ;
 END
 PORT
  LAYER ME4 ;
  RECT 313.903 0.000 314.623 44.094 ;
 END
 PORT
  LAYER ME4 ;
  RECT 319.098 1.781 319.438 66.831 ;
 END
 PORT
  LAYER ME4 ;
  RECT 317.096 1.781 317.436 66.831 ;
 END
 PORT
  LAYER ME4 ;
  RECT 317.907 0.000 318.627 44.094 ;
 END
 PORT
  LAYER ME4 ;
  RECT 323.102 1.781 323.442 66.831 ;
 END
 PORT
  LAYER ME4 ;
  RECT 321.100 1.781 321.440 66.831 ;
 END
 PORT
  LAYER ME4 ;
  RECT 321.911 0.000 322.631 44.094 ;
 END
 PORT
  LAYER ME4 ;
  RECT 327.106 1.781 327.446 66.831 ;
 END
 PORT
  LAYER ME4 ;
  RECT 325.104 1.781 325.444 66.831 ;
 END
 PORT
  LAYER ME4 ;
  RECT 325.915 0.000 326.635 44.094 ;
 END
 PORT
  LAYER ME4 ;
  RECT 331.110 1.781 331.450 66.831 ;
 END
 PORT
  LAYER ME4 ;
  RECT 329.108 1.781 329.448 66.831 ;
 END
 PORT
  LAYER ME4 ;
  RECT 329.919 0.000 330.639 44.094 ;
 END
 PORT
  LAYER ME4 ;
  RECT 335.114 1.781 335.454 66.831 ;
 END
 PORT
  LAYER ME4 ;
  RECT 333.112 1.781 333.452 66.831 ;
 END
 PORT
  LAYER ME4 ;
  RECT 333.923 0.000 334.643 44.094 ;
 END
 PORT
  LAYER ME4 ;
  RECT 339.118 1.781 339.458 66.831 ;
 END
 PORT
  LAYER ME4 ;
  RECT 337.116 1.781 337.456 66.831 ;
 END
 PORT
  LAYER ME4 ;
  RECT 337.927 0.000 338.647 44.094 ;
 END
 PORT
  LAYER ME4 ;
  RECT 343.122 1.781 343.462 66.831 ;
 END
 PORT
  LAYER ME4 ;
  RECT 341.120 1.781 341.460 66.831 ;
 END
 PORT
  LAYER ME4 ;
  RECT 341.931 0.000 342.651 44.094 ;
 END
 PORT
  LAYER ME4 ;
  RECT 347.126 1.781 347.466 66.831 ;
 END
 PORT
  LAYER ME4 ;
  RECT 345.124 1.781 345.464 66.831 ;
 END
 PORT
  LAYER ME4 ;
  RECT 345.935 0.000 346.655 44.094 ;
 END
 PORT
  LAYER ME4 ;
  RECT 351.130 1.781 351.470 66.831 ;
 END
 PORT
  LAYER ME4 ;
  RECT 349.128 1.781 349.468 66.831 ;
 END
 PORT
  LAYER ME4 ;
  RECT 349.939 0.000 350.659 44.094 ;
 END
 PORT
  LAYER ME4 ;
  RECT 355.134 1.781 355.474 66.831 ;
 END
 PORT
  LAYER ME4 ;
  RECT 353.132 1.781 353.472 66.831 ;
 END
 PORT
  LAYER ME4 ;
  RECT 353.943 0.000 354.663 44.094 ;
 END
 PORT
  LAYER ME4 ;
  RECT 359.138 1.781 359.478 66.831 ;
 END
 PORT
  LAYER ME4 ;
  RECT 357.136 1.781 357.476 66.831 ;
 END
 PORT
  LAYER ME4 ;
  RECT 357.947 0.000 358.667 44.094 ;
 END
 PORT
  LAYER ME4 ;
  RECT 363.142 1.781 363.482 66.831 ;
 END
 PORT
  LAYER ME4 ;
  RECT 361.140 1.781 361.480 66.831 ;
 END
 PORT
  LAYER ME4 ;
  RECT 361.951 0.000 362.671 44.094 ;
 END
 PORT
  LAYER ME4 ;
  RECT 367.146 1.781 367.486 66.831 ;
 END
 PORT
  LAYER ME4 ;
  RECT 365.144 1.781 365.484 66.831 ;
 END
 PORT
  LAYER ME4 ;
  RECT 365.955 0.000 366.675 44.094 ;
 END
 PORT
  LAYER ME4 ;
  RECT 371.150 1.781 371.490 66.831 ;
 END
 PORT
  LAYER ME4 ;
  RECT 369.148 1.781 369.488 66.831 ;
 END
 PORT
  LAYER ME4 ;
  RECT 369.959 0.000 370.679 44.094 ;
 END
 PORT
  LAYER ME4 ;
  RECT 375.154 1.781 375.494 66.831 ;
 END
 PORT
  LAYER ME4 ;
  RECT 373.152 1.781 373.492 66.831 ;
 END
 PORT
  LAYER ME4 ;
  RECT 373.963 0.000 374.683 44.094 ;
 END
 PORT
  LAYER ME4 ;
  RECT 379.158 1.781 379.498 66.831 ;
 END
 PORT
  LAYER ME4 ;
  RECT 377.156 1.781 377.496 66.831 ;
 END
 PORT
  LAYER ME4 ;
  RECT 377.967 0.000 378.687 44.094 ;
 END
 PORT
  LAYER ME4 ;
  RECT 383.162 1.781 383.502 66.831 ;
 END
 PORT
  LAYER ME4 ;
  RECT 381.160 1.781 381.500 66.831 ;
 END
 PORT
  LAYER ME4 ;
  RECT 381.971 0.000 382.691 44.094 ;
 END
 PORT
  LAYER ME4 ;
  RECT 387.166 1.781 387.506 66.831 ;
 END
 PORT
  LAYER ME4 ;
  RECT 385.164 1.781 385.504 66.831 ;
 END
 PORT
  LAYER ME4 ;
  RECT 385.975 0.000 386.695 44.094 ;
 END
 PORT
  LAYER ME4 ;
  RECT 391.170 1.781 391.510 66.831 ;
 END
 PORT
  LAYER ME4 ;
  RECT 389.168 1.781 389.508 66.831 ;
 END
 PORT
  LAYER ME4 ;
  RECT 389.979 0.000 390.699 44.094 ;
 END
 PORT
  LAYER ME4 ;
  RECT 392.171 0.000 392.511 66.831 ;
 END
 PORT
  LAYER ME4 ;
  RECT 196.137 0.000 196.857 66.831 ;
 END
 PORT
  LAYER ME4 ;
  RECT 202.131 0.000 202.851 66.831 ;
 END
 PORT
  LAYER ME4 ;
  RECT 207.602 0.000 208.322 66.831 ;
 END
 PORT
  LAYER ME4 ;
  RECT 209.317 0.000 210.037 66.831 ;
 END
 PORT
  LAYER ME4 ;
  RECT 212.313 0.000 212.913 66.831 ;
 END
 PORT
  LAYER ME4 ;
  RECT 213.993 1.781 214.333 66.831 ;
 END
 PORT
  LAYER ME4 ;
  RECT 188.578 0.000 189.298 66.831 ;
 END
 PORT
  LAYER ME4 ;
  RECT 186.538 1.781 187.258 66.072 ;
 END
 PORT
  LAYER ME4 ;
  RECT 1.740 0.000 2.080 66.831 ;
 END
 PORT
  LAYER ME4 ;
  RECT 6.745 1.781 7.085 66.831 ;
 END
 PORT
  LAYER ME4 ;
  RECT 2.741 1.781 3.081 66.831 ;
 END
 PORT
  LAYER ME4 ;
  RECT 4.743 1.781 5.083 66.831 ;
 END
 PORT
  LAYER ME4 ;
  RECT 5.554 0.000 6.274 44.094 ;
 END
 PORT
  LAYER ME4 ;
  RECT 10.749 1.781 11.089 66.831 ;
 END
 PORT
  LAYER ME4 ;
  RECT 8.747 1.781 9.087 66.831 ;
 END
 PORT
  LAYER ME4 ;
  RECT 9.558 0.000 10.278 44.094 ;
 END
 PORT
  LAYER ME4 ;
  RECT 14.753 1.781 15.093 66.831 ;
 END
 PORT
  LAYER ME4 ;
  RECT 12.751 1.781 13.091 66.831 ;
 END
 PORT
  LAYER ME4 ;
  RECT 13.562 0.000 14.282 44.094 ;
 END
 PORT
  LAYER ME4 ;
  RECT 18.757 1.781 19.097 66.831 ;
 END
 PORT
  LAYER ME4 ;
  RECT 16.755 1.781 17.095 66.831 ;
 END
 PORT
  LAYER ME4 ;
  RECT 17.566 0.000 18.286 44.094 ;
 END
 PORT
  LAYER ME4 ;
  RECT 22.761 1.781 23.101 66.831 ;
 END
 PORT
  LAYER ME4 ;
  RECT 20.759 1.781 21.099 66.831 ;
 END
 PORT
  LAYER ME4 ;
  RECT 21.570 0.000 22.290 44.094 ;
 END
 PORT
  LAYER ME4 ;
  RECT 26.765 1.781 27.105 66.831 ;
 END
 PORT
  LAYER ME4 ;
  RECT 24.763 1.781 25.103 66.831 ;
 END
 PORT
  LAYER ME4 ;
  RECT 25.574 0.000 26.294 44.094 ;
 END
 PORT
  LAYER ME4 ;
  RECT 30.769 1.781 31.109 66.831 ;
 END
 PORT
  LAYER ME4 ;
  RECT 28.767 1.781 29.107 66.831 ;
 END
 PORT
  LAYER ME4 ;
  RECT 29.578 0.000 30.298 44.094 ;
 END
 PORT
  LAYER ME4 ;
  RECT 34.773 1.781 35.113 66.831 ;
 END
 PORT
  LAYER ME4 ;
  RECT 32.771 1.781 33.111 66.831 ;
 END
 PORT
  LAYER ME4 ;
  RECT 33.582 0.000 34.302 44.094 ;
 END
 PORT
  LAYER ME4 ;
  RECT 38.777 1.781 39.117 66.831 ;
 END
 PORT
  LAYER ME4 ;
  RECT 36.775 1.781 37.115 66.831 ;
 END
 PORT
  LAYER ME4 ;
  RECT 37.586 0.000 38.306 44.094 ;
 END
 PORT
  LAYER ME4 ;
  RECT 42.781 1.781 43.121 66.831 ;
 END
 PORT
  LAYER ME4 ;
  RECT 40.779 1.781 41.119 66.831 ;
 END
 PORT
  LAYER ME4 ;
  RECT 41.590 0.000 42.310 44.094 ;
 END
 PORT
  LAYER ME4 ;
  RECT 46.785 1.781 47.125 66.831 ;
 END
 PORT
  LAYER ME4 ;
  RECT 44.783 1.781 45.123 66.831 ;
 END
 PORT
  LAYER ME4 ;
  RECT 45.594 0.000 46.314 44.094 ;
 END
 PORT
  LAYER ME4 ;
  RECT 50.789 1.781 51.129 66.831 ;
 END
 PORT
  LAYER ME4 ;
  RECT 48.787 1.781 49.127 66.831 ;
 END
 PORT
  LAYER ME4 ;
  RECT 49.598 0.000 50.318 44.094 ;
 END
 PORT
  LAYER ME4 ;
  RECT 54.793 1.781 55.133 66.831 ;
 END
 PORT
  LAYER ME4 ;
  RECT 52.791 1.781 53.131 66.831 ;
 END
 PORT
  LAYER ME4 ;
  RECT 53.602 0.000 54.322 44.094 ;
 END
 PORT
  LAYER ME4 ;
  RECT 58.797 1.781 59.137 66.831 ;
 END
 PORT
  LAYER ME4 ;
  RECT 56.795 1.781 57.135 66.831 ;
 END
 PORT
  LAYER ME4 ;
  RECT 57.606 0.000 58.326 44.094 ;
 END
 PORT
  LAYER ME4 ;
  RECT 62.801 1.781 63.141 66.831 ;
 END
 PORT
  LAYER ME4 ;
  RECT 60.799 1.781 61.139 66.831 ;
 END
 PORT
  LAYER ME4 ;
  RECT 61.610 0.000 62.330 44.094 ;
 END
 PORT
  LAYER ME4 ;
  RECT 66.805 1.781 67.145 66.831 ;
 END
 PORT
  LAYER ME4 ;
  RECT 64.803 1.781 65.143 66.831 ;
 END
 PORT
  LAYER ME4 ;
  RECT 65.614 0.000 66.334 44.094 ;
 END
 PORT
  LAYER ME4 ;
  RECT 70.809 1.781 71.149 66.831 ;
 END
 PORT
  LAYER ME4 ;
  RECT 68.807 1.781 69.147 66.831 ;
 END
 PORT
  LAYER ME4 ;
  RECT 69.618 0.000 70.338 44.094 ;
 END
 PORT
  LAYER ME4 ;
  RECT 74.813 1.781 75.153 66.831 ;
 END
 PORT
  LAYER ME4 ;
  RECT 72.811 1.781 73.151 66.831 ;
 END
 PORT
  LAYER ME4 ;
  RECT 73.622 0.000 74.342 44.094 ;
 END
 PORT
  LAYER ME4 ;
  RECT 78.817 1.781 79.157 66.831 ;
 END
 PORT
  LAYER ME4 ;
  RECT 76.815 1.781 77.155 66.831 ;
 END
 PORT
  LAYER ME4 ;
  RECT 77.626 0.000 78.346 44.094 ;
 END
 PORT
  LAYER ME4 ;
  RECT 82.821 1.781 83.161 66.831 ;
 END
 PORT
  LAYER ME4 ;
  RECT 80.819 1.781 81.159 66.831 ;
 END
 PORT
  LAYER ME4 ;
  RECT 81.630 0.000 82.350 44.094 ;
 END
 PORT
  LAYER ME4 ;
  RECT 86.825 1.781 87.165 66.831 ;
 END
 PORT
  LAYER ME4 ;
  RECT 84.823 1.781 85.163 66.831 ;
 END
 PORT
  LAYER ME4 ;
  RECT 85.634 0.000 86.354 44.094 ;
 END
 PORT
  LAYER ME4 ;
  RECT 90.829 1.781 91.169 66.831 ;
 END
 PORT
  LAYER ME4 ;
  RECT 88.827 1.781 89.167 66.831 ;
 END
 PORT
  LAYER ME4 ;
  RECT 89.638 0.000 90.358 44.094 ;
 END
 PORT
  LAYER ME4 ;
  RECT 94.833 1.781 95.173 66.831 ;
 END
 PORT
  LAYER ME4 ;
  RECT 92.831 1.781 93.171 66.831 ;
 END
 PORT
  LAYER ME4 ;
  RECT 93.642 0.000 94.362 44.094 ;
 END
 PORT
  LAYER ME4 ;
  RECT 98.837 1.781 99.177 66.831 ;
 END
 PORT
  LAYER ME4 ;
  RECT 96.835 1.781 97.175 66.831 ;
 END
 PORT
  LAYER ME4 ;
  RECT 97.646 0.000 98.366 44.094 ;
 END
 PORT
  LAYER ME4 ;
  RECT 102.841 1.781 103.181 66.831 ;
 END
 PORT
  LAYER ME4 ;
  RECT 100.839 1.781 101.179 66.831 ;
 END
 PORT
  LAYER ME4 ;
  RECT 101.650 0.000 102.370 44.094 ;
 END
 PORT
  LAYER ME4 ;
  RECT 106.845 1.781 107.185 66.831 ;
 END
 PORT
  LAYER ME4 ;
  RECT 104.843 1.781 105.183 66.831 ;
 END
 PORT
  LAYER ME4 ;
  RECT 105.654 0.000 106.374 44.094 ;
 END
 PORT
  LAYER ME4 ;
  RECT 110.849 1.781 111.189 66.831 ;
 END
 PORT
  LAYER ME4 ;
  RECT 108.847 1.781 109.187 66.831 ;
 END
 PORT
  LAYER ME4 ;
  RECT 109.658 0.000 110.378 44.094 ;
 END
 PORT
  LAYER ME4 ;
  RECT 114.853 1.781 115.193 66.831 ;
 END
 PORT
  LAYER ME4 ;
  RECT 112.851 1.781 113.191 66.831 ;
 END
 PORT
  LAYER ME4 ;
  RECT 113.662 0.000 114.382 44.094 ;
 END
 PORT
  LAYER ME4 ;
  RECT 118.857 1.781 119.197 66.831 ;
 END
 PORT
  LAYER ME4 ;
  RECT 116.855 1.781 117.195 66.831 ;
 END
 PORT
  LAYER ME4 ;
  RECT 117.666 0.000 118.386 44.094 ;
 END
 PORT
  LAYER ME4 ;
  RECT 122.861 1.781 123.201 66.831 ;
 END
 PORT
  LAYER ME4 ;
  RECT 120.859 1.781 121.199 66.831 ;
 END
 PORT
  LAYER ME4 ;
  RECT 121.670 0.000 122.390 44.094 ;
 END
 PORT
  LAYER ME4 ;
  RECT 126.865 1.781 127.205 66.831 ;
 END
 PORT
  LAYER ME4 ;
  RECT 124.863 1.781 125.203 66.831 ;
 END
 PORT
  LAYER ME4 ;
  RECT 125.674 0.000 126.394 44.094 ;
 END
 PORT
  LAYER ME4 ;
  RECT 130.869 1.781 131.209 66.831 ;
 END
 PORT
  LAYER ME4 ;
  RECT 128.867 1.781 129.207 66.831 ;
 END
 PORT
  LAYER ME4 ;
  RECT 129.678 0.000 130.398 44.094 ;
 END
 PORT
  LAYER ME4 ;
  RECT 134.873 1.781 135.213 66.831 ;
 END
 PORT
  LAYER ME4 ;
  RECT 132.871 1.781 133.211 66.831 ;
 END
 PORT
  LAYER ME4 ;
  RECT 133.682 0.000 134.402 44.094 ;
 END
 PORT
  LAYER ME4 ;
  RECT 138.877 1.781 139.217 66.831 ;
 END
 PORT
  LAYER ME4 ;
  RECT 136.875 1.781 137.215 66.831 ;
 END
 PORT
  LAYER ME4 ;
  RECT 137.686 0.000 138.406 44.094 ;
 END
 PORT
  LAYER ME4 ;
  RECT 142.881 1.781 143.221 66.831 ;
 END
 PORT
  LAYER ME4 ;
  RECT 140.879 1.781 141.219 66.831 ;
 END
 PORT
  LAYER ME4 ;
  RECT 141.690 0.000 142.410 44.094 ;
 END
 PORT
  LAYER ME4 ;
  RECT 146.885 1.781 147.225 66.831 ;
 END
 PORT
  LAYER ME4 ;
  RECT 144.883 1.781 145.223 66.831 ;
 END
 PORT
  LAYER ME4 ;
  RECT 145.694 0.000 146.414 44.094 ;
 END
 PORT
  LAYER ME4 ;
  RECT 150.889 1.781 151.229 66.831 ;
 END
 PORT
  LAYER ME4 ;
  RECT 148.887 1.781 149.227 66.831 ;
 END
 PORT
  LAYER ME4 ;
  RECT 149.698 0.000 150.418 44.094 ;
 END
 PORT
  LAYER ME4 ;
  RECT 154.893 1.781 155.233 66.831 ;
 END
 PORT
  LAYER ME4 ;
  RECT 152.891 1.781 153.231 66.831 ;
 END
 PORT
  LAYER ME4 ;
  RECT 153.702 0.000 154.422 44.094 ;
 END
 PORT
  LAYER ME4 ;
  RECT 158.897 1.781 159.237 66.831 ;
 END
 PORT
  LAYER ME4 ;
  RECT 156.895 1.781 157.235 66.831 ;
 END
 PORT
  LAYER ME4 ;
  RECT 157.706 0.000 158.426 44.094 ;
 END
 PORT
  LAYER ME4 ;
  RECT 162.901 1.781 163.241 66.831 ;
 END
 PORT
  LAYER ME4 ;
  RECT 160.899 1.781 161.239 66.831 ;
 END
 PORT
  LAYER ME4 ;
  RECT 161.710 0.000 162.430 44.094 ;
 END
 PORT
  LAYER ME4 ;
  RECT 166.905 1.781 167.245 66.831 ;
 END
 PORT
  LAYER ME4 ;
  RECT 164.903 1.781 165.243 66.831 ;
 END
 PORT
  LAYER ME4 ;
  RECT 165.714 0.000 166.434 44.094 ;
 END
 PORT
  LAYER ME4 ;
  RECT 170.909 1.781 171.249 66.831 ;
 END
 PORT
  LAYER ME4 ;
  RECT 168.907 1.781 169.247 66.831 ;
 END
 PORT
  LAYER ME4 ;
  RECT 169.718 0.000 170.438 44.094 ;
 END
 PORT
  LAYER ME4 ;
  RECT 174.913 1.781 175.253 66.831 ;
 END
 PORT
  LAYER ME4 ;
  RECT 172.911 1.781 173.251 66.831 ;
 END
 PORT
  LAYER ME4 ;
  RECT 173.722 0.000 174.442 44.094 ;
 END
 PORT
  LAYER ME4 ;
  RECT 178.917 1.781 179.257 66.831 ;
 END
 PORT
  LAYER ME4 ;
  RECT 176.915 1.781 177.255 66.831 ;
 END
 PORT
  LAYER ME4 ;
  RECT 177.726 0.000 178.446 44.094 ;
 END
 PORT
  LAYER ME4 ;
  RECT 184.418 0.000 185.138 66.831 ;
 END
 PORT
  LAYER ME4 ;
  RECT 182.378 0.000 183.098 66.831 ;
 END
 PORT
  LAYER ME4 ;
  RECT 179.918 0.000 180.258 66.831 ;
 END
END GND
PIN VCC
  DIRECTION INOUT ;
  USE POWER ;
 PORT
  LAYER ME4 ;
  RECT 217.997 45.394 218.337 66.831 ;
 END
 PORT
  LAYER ME4 ;
  RECT 215.805 0.000 216.525 46.394 ;
 END
 PORT
  LAYER ME4 ;
  RECT 222.001 45.394 222.341 66.831 ;
 END
 PORT
  LAYER ME4 ;
  RECT 219.809 0.000 220.529 46.394 ;
 END
 PORT
  LAYER ME4 ;
  RECT 226.005 45.394 226.345 66.831 ;
 END
 PORT
  LAYER ME4 ;
  RECT 223.813 0.000 224.533 46.394 ;
 END
 PORT
  LAYER ME4 ;
  RECT 230.009 45.394 230.349 66.831 ;
 END
 PORT
  LAYER ME4 ;
  RECT 227.817 0.000 228.537 46.394 ;
 END
 PORT
  LAYER ME4 ;
  RECT 234.013 45.394 234.353 66.831 ;
 END
 PORT
  LAYER ME4 ;
  RECT 231.821 0.000 232.541 46.394 ;
 END
 PORT
  LAYER ME4 ;
  RECT 238.017 45.394 238.357 66.831 ;
 END
 PORT
  LAYER ME4 ;
  RECT 235.825 0.000 236.545 46.394 ;
 END
 PORT
  LAYER ME4 ;
  RECT 242.021 45.394 242.361 66.831 ;
 END
 PORT
  LAYER ME4 ;
  RECT 239.829 0.000 240.549 46.394 ;
 END
 PORT
  LAYER ME4 ;
  RECT 246.025 45.394 246.365 66.831 ;
 END
 PORT
  LAYER ME4 ;
  RECT 243.833 0.000 244.553 46.394 ;
 END
 PORT
  LAYER ME4 ;
  RECT 250.029 45.394 250.369 66.831 ;
 END
 PORT
  LAYER ME4 ;
  RECT 247.837 0.000 248.557 46.394 ;
 END
 PORT
  LAYER ME4 ;
  RECT 254.033 45.394 254.373 66.831 ;
 END
 PORT
  LAYER ME4 ;
  RECT 251.841 0.000 252.561 46.394 ;
 END
 PORT
  LAYER ME4 ;
  RECT 258.037 45.394 258.377 66.831 ;
 END
 PORT
  LAYER ME4 ;
  RECT 255.845 0.000 256.565 46.394 ;
 END
 PORT
  LAYER ME4 ;
  RECT 262.041 45.394 262.381 66.831 ;
 END
 PORT
  LAYER ME4 ;
  RECT 259.849 0.000 260.569 46.394 ;
 END
 PORT
  LAYER ME4 ;
  RECT 266.045 45.394 266.385 66.831 ;
 END
 PORT
  LAYER ME4 ;
  RECT 263.853 0.000 264.573 46.394 ;
 END
 PORT
  LAYER ME4 ;
  RECT 270.049 45.394 270.389 66.831 ;
 END
 PORT
  LAYER ME4 ;
  RECT 267.857 0.000 268.577 46.394 ;
 END
 PORT
  LAYER ME4 ;
  RECT 274.053 45.394 274.393 66.831 ;
 END
 PORT
  LAYER ME4 ;
  RECT 271.861 0.000 272.581 46.394 ;
 END
 PORT
  LAYER ME4 ;
  RECT 278.057 45.394 278.397 66.831 ;
 END
 PORT
  LAYER ME4 ;
  RECT 275.865 0.000 276.585 46.394 ;
 END
 PORT
  LAYER ME4 ;
  RECT 282.061 45.394 282.401 66.831 ;
 END
 PORT
  LAYER ME4 ;
  RECT 279.869 0.000 280.589 46.394 ;
 END
 PORT
  LAYER ME4 ;
  RECT 286.065 45.394 286.405 66.831 ;
 END
 PORT
  LAYER ME4 ;
  RECT 283.873 0.000 284.593 46.394 ;
 END
 PORT
  LAYER ME4 ;
  RECT 290.069 45.394 290.409 66.831 ;
 END
 PORT
  LAYER ME4 ;
  RECT 287.877 0.000 288.597 46.394 ;
 END
 PORT
  LAYER ME4 ;
  RECT 294.073 45.394 294.413 66.831 ;
 END
 PORT
  LAYER ME4 ;
  RECT 291.881 0.000 292.601 46.394 ;
 END
 PORT
  LAYER ME4 ;
  RECT 298.077 45.394 298.417 66.831 ;
 END
 PORT
  LAYER ME4 ;
  RECT 295.885 0.000 296.605 46.394 ;
 END
 PORT
  LAYER ME4 ;
  RECT 302.081 45.394 302.421 66.831 ;
 END
 PORT
  LAYER ME4 ;
  RECT 299.889 0.000 300.609 46.394 ;
 END
 PORT
  LAYER ME4 ;
  RECT 306.085 45.394 306.425 66.831 ;
 END
 PORT
  LAYER ME4 ;
  RECT 303.893 0.000 304.613 46.394 ;
 END
 PORT
  LAYER ME4 ;
  RECT 310.089 45.394 310.429 66.831 ;
 END
 PORT
  LAYER ME4 ;
  RECT 307.897 0.000 308.617 46.394 ;
 END
 PORT
  LAYER ME4 ;
  RECT 314.093 45.394 314.433 66.831 ;
 END
 PORT
  LAYER ME4 ;
  RECT 311.901 0.000 312.621 46.394 ;
 END
 PORT
  LAYER ME4 ;
  RECT 318.097 45.394 318.437 66.831 ;
 END
 PORT
  LAYER ME4 ;
  RECT 315.905 0.000 316.625 46.394 ;
 END
 PORT
  LAYER ME4 ;
  RECT 322.101 45.394 322.441 66.831 ;
 END
 PORT
  LAYER ME4 ;
  RECT 319.909 0.000 320.629 46.394 ;
 END
 PORT
  LAYER ME4 ;
  RECT 326.105 45.394 326.445 66.831 ;
 END
 PORT
  LAYER ME4 ;
  RECT 323.913 0.000 324.633 46.394 ;
 END
 PORT
  LAYER ME4 ;
  RECT 330.109 45.394 330.449 66.831 ;
 END
 PORT
  LAYER ME4 ;
  RECT 327.917 0.000 328.637 46.394 ;
 END
 PORT
  LAYER ME4 ;
  RECT 334.113 45.394 334.453 66.831 ;
 END
 PORT
  LAYER ME4 ;
  RECT 331.921 0.000 332.641 46.394 ;
 END
 PORT
  LAYER ME4 ;
  RECT 338.117 45.394 338.457 66.831 ;
 END
 PORT
  LAYER ME4 ;
  RECT 335.925 0.000 336.645 46.394 ;
 END
 PORT
  LAYER ME4 ;
  RECT 342.121 45.394 342.461 66.831 ;
 END
 PORT
  LAYER ME4 ;
  RECT 339.929 0.000 340.649 46.394 ;
 END
 PORT
  LAYER ME4 ;
  RECT 346.125 45.394 346.465 66.831 ;
 END
 PORT
  LAYER ME4 ;
  RECT 343.933 0.000 344.653 46.394 ;
 END
 PORT
  LAYER ME4 ;
  RECT 350.129 45.394 350.469 66.831 ;
 END
 PORT
  LAYER ME4 ;
  RECT 347.937 0.000 348.657 46.394 ;
 END
 PORT
  LAYER ME4 ;
  RECT 354.133 45.394 354.473 66.831 ;
 END
 PORT
  LAYER ME4 ;
  RECT 351.941 0.000 352.661 46.394 ;
 END
 PORT
  LAYER ME4 ;
  RECT 358.137 45.394 358.477 66.831 ;
 END
 PORT
  LAYER ME4 ;
  RECT 355.945 0.000 356.665 46.394 ;
 END
 PORT
  LAYER ME4 ;
  RECT 362.141 45.394 362.481 66.831 ;
 END
 PORT
  LAYER ME4 ;
  RECT 359.949 0.000 360.669 46.394 ;
 END
 PORT
  LAYER ME4 ;
  RECT 366.145 45.394 366.485 66.831 ;
 END
 PORT
  LAYER ME4 ;
  RECT 363.953 0.000 364.673 46.394 ;
 END
 PORT
  LAYER ME4 ;
  RECT 370.149 45.394 370.489 66.831 ;
 END
 PORT
  LAYER ME4 ;
  RECT 367.957 0.000 368.677 46.394 ;
 END
 PORT
  LAYER ME4 ;
  RECT 374.153 45.394 374.493 66.831 ;
 END
 PORT
  LAYER ME4 ;
  RECT 371.961 0.000 372.681 46.394 ;
 END
 PORT
  LAYER ME4 ;
  RECT 378.157 45.394 378.497 66.831 ;
 END
 PORT
  LAYER ME4 ;
  RECT 375.965 0.000 376.685 46.394 ;
 END
 PORT
  LAYER ME4 ;
  RECT 382.161 45.394 382.501 66.831 ;
 END
 PORT
  LAYER ME4 ;
  RECT 379.969 0.000 380.689 46.394 ;
 END
 PORT
  LAYER ME4 ;
  RECT 386.165 45.394 386.505 66.831 ;
 END
 PORT
  LAYER ME4 ;
  RECT 383.973 0.000 384.693 46.394 ;
 END
 PORT
  LAYER ME4 ;
  RECT 390.169 45.394 390.509 66.831 ;
 END
 PORT
  LAYER ME4 ;
  RECT 387.977 0.000 388.697 46.394 ;
 END
 PORT
  LAYER ME4 ;
  RECT 392.951 0.000 393.331 66.831 ;
 END
 PORT
  LAYER ME4 ;
  RECT 198.917 0.000 199.517 66.831 ;
 END
 PORT
  LAYER ME4 ;
  RECT 203.097 0.000 203.817 66.831 ;
 END
 PORT
  LAYER ME4 ;
  RECT 205.207 0.000 206.327 66.831 ;
 END
 PORT
  LAYER ME4 ;
  RECT 211.237 0.000 211.957 66.831 ;
 END
 PORT
  LAYER ME4 ;
  RECT 213.173 1.781 213.553 66.831 ;
 END
 PORT
  LAYER ME4 ;
  RECT 194.687 0.000 195.407 66.831 ;
 END
 PORT
  LAYER ME4 ;
  RECT 191.972 0.000 193.092 66.831 ;
 END
 PORT
  LAYER ME4 ;
  RECT 189.598 0.000 190.318 66.072 ;
 END
 PORT
  LAYER ME4 ;
  RECT 187.558 1.781 188.278 66.831 ;
 END
 PORT
  LAYER ME4 ;
  RECT 0.920 0.000 1.300 66.831 ;
 END
 PORT
  LAYER ME4 ;
  RECT 5.744 45.394 6.084 66.831 ;
 END
 PORT
  LAYER ME4 ;
  RECT 3.552 0.000 4.272 46.394 ;
 END
 PORT
  LAYER ME4 ;
  RECT 9.748 45.394 10.088 66.831 ;
 END
 PORT
  LAYER ME4 ;
  RECT 7.556 0.000 8.276 46.394 ;
 END
 PORT
  LAYER ME4 ;
  RECT 13.752 45.394 14.092 66.831 ;
 END
 PORT
  LAYER ME4 ;
  RECT 11.560 0.000 12.280 46.394 ;
 END
 PORT
  LAYER ME4 ;
  RECT 17.756 45.394 18.096 66.831 ;
 END
 PORT
  LAYER ME4 ;
  RECT 15.564 0.000 16.284 46.394 ;
 END
 PORT
  LAYER ME4 ;
  RECT 21.760 45.394 22.100 66.831 ;
 END
 PORT
  LAYER ME4 ;
  RECT 19.568 0.000 20.288 46.394 ;
 END
 PORT
  LAYER ME4 ;
  RECT 25.764 45.394 26.104 66.831 ;
 END
 PORT
  LAYER ME4 ;
  RECT 23.572 0.000 24.292 46.394 ;
 END
 PORT
  LAYER ME4 ;
  RECT 29.768 45.394 30.108 66.831 ;
 END
 PORT
  LAYER ME4 ;
  RECT 27.576 0.000 28.296 46.394 ;
 END
 PORT
  LAYER ME4 ;
  RECT 33.772 45.394 34.112 66.831 ;
 END
 PORT
  LAYER ME4 ;
  RECT 31.580 0.000 32.300 46.394 ;
 END
 PORT
  LAYER ME4 ;
  RECT 37.776 45.394 38.116 66.831 ;
 END
 PORT
  LAYER ME4 ;
  RECT 35.584 0.000 36.304 46.394 ;
 END
 PORT
  LAYER ME4 ;
  RECT 41.780 45.394 42.120 66.831 ;
 END
 PORT
  LAYER ME4 ;
  RECT 39.588 0.000 40.308 46.394 ;
 END
 PORT
  LAYER ME4 ;
  RECT 45.784 45.394 46.124 66.831 ;
 END
 PORT
  LAYER ME4 ;
  RECT 43.592 0.000 44.312 46.394 ;
 END
 PORT
  LAYER ME4 ;
  RECT 49.788 45.394 50.128 66.831 ;
 END
 PORT
  LAYER ME4 ;
  RECT 47.596 0.000 48.316 46.394 ;
 END
 PORT
  LAYER ME4 ;
  RECT 53.792 45.394 54.132 66.831 ;
 END
 PORT
  LAYER ME4 ;
  RECT 51.600 0.000 52.320 46.394 ;
 END
 PORT
  LAYER ME4 ;
  RECT 57.796 45.394 58.136 66.831 ;
 END
 PORT
  LAYER ME4 ;
  RECT 55.604 0.000 56.324 46.394 ;
 END
 PORT
  LAYER ME4 ;
  RECT 61.800 45.394 62.140 66.831 ;
 END
 PORT
  LAYER ME4 ;
  RECT 59.608 0.000 60.328 46.394 ;
 END
 PORT
  LAYER ME4 ;
  RECT 65.804 45.394 66.144 66.831 ;
 END
 PORT
  LAYER ME4 ;
  RECT 63.612 0.000 64.332 46.394 ;
 END
 PORT
  LAYER ME4 ;
  RECT 69.808 45.394 70.148 66.831 ;
 END
 PORT
  LAYER ME4 ;
  RECT 67.616 0.000 68.336 46.394 ;
 END
 PORT
  LAYER ME4 ;
  RECT 73.812 45.394 74.152 66.831 ;
 END
 PORT
  LAYER ME4 ;
  RECT 71.620 0.000 72.340 46.394 ;
 END
 PORT
  LAYER ME4 ;
  RECT 77.816 45.394 78.156 66.831 ;
 END
 PORT
  LAYER ME4 ;
  RECT 75.624 0.000 76.344 46.394 ;
 END
 PORT
  LAYER ME4 ;
  RECT 81.820 45.394 82.160 66.831 ;
 END
 PORT
  LAYER ME4 ;
  RECT 79.628 0.000 80.348 46.394 ;
 END
 PORT
  LAYER ME4 ;
  RECT 85.824 45.394 86.164 66.831 ;
 END
 PORT
  LAYER ME4 ;
  RECT 83.632 0.000 84.352 46.394 ;
 END
 PORT
  LAYER ME4 ;
  RECT 89.828 45.394 90.168 66.831 ;
 END
 PORT
  LAYER ME4 ;
  RECT 87.636 0.000 88.356 46.394 ;
 END
 PORT
  LAYER ME4 ;
  RECT 93.832 45.394 94.172 66.831 ;
 END
 PORT
  LAYER ME4 ;
  RECT 91.640 0.000 92.360 46.394 ;
 END
 PORT
  LAYER ME4 ;
  RECT 97.836 45.394 98.176 66.831 ;
 END
 PORT
  LAYER ME4 ;
  RECT 95.644 0.000 96.364 46.394 ;
 END
 PORT
  LAYER ME4 ;
  RECT 101.840 45.394 102.180 66.831 ;
 END
 PORT
  LAYER ME4 ;
  RECT 99.648 0.000 100.368 46.394 ;
 END
 PORT
  LAYER ME4 ;
  RECT 105.844 45.394 106.184 66.831 ;
 END
 PORT
  LAYER ME4 ;
  RECT 103.652 0.000 104.372 46.394 ;
 END
 PORT
  LAYER ME4 ;
  RECT 109.848 45.394 110.188 66.831 ;
 END
 PORT
  LAYER ME4 ;
  RECT 107.656 0.000 108.376 46.394 ;
 END
 PORT
  LAYER ME4 ;
  RECT 113.852 45.394 114.192 66.831 ;
 END
 PORT
  LAYER ME4 ;
  RECT 111.660 0.000 112.380 46.394 ;
 END
 PORT
  LAYER ME4 ;
  RECT 117.856 45.394 118.196 66.831 ;
 END
 PORT
  LAYER ME4 ;
  RECT 115.664 0.000 116.384 46.394 ;
 END
 PORT
  LAYER ME4 ;
  RECT 121.860 45.394 122.200 66.831 ;
 END
 PORT
  LAYER ME4 ;
  RECT 119.668 0.000 120.388 46.394 ;
 END
 PORT
  LAYER ME4 ;
  RECT 125.864 45.394 126.204 66.831 ;
 END
 PORT
  LAYER ME4 ;
  RECT 123.672 0.000 124.392 46.394 ;
 END
 PORT
  LAYER ME4 ;
  RECT 129.868 45.394 130.208 66.831 ;
 END
 PORT
  LAYER ME4 ;
  RECT 127.676 0.000 128.396 46.394 ;
 END
 PORT
  LAYER ME4 ;
  RECT 133.872 45.394 134.212 66.831 ;
 END
 PORT
  LAYER ME4 ;
  RECT 131.680 0.000 132.400 46.394 ;
 END
 PORT
  LAYER ME4 ;
  RECT 137.876 45.394 138.216 66.831 ;
 END
 PORT
  LAYER ME4 ;
  RECT 135.684 0.000 136.404 46.394 ;
 END
 PORT
  LAYER ME4 ;
  RECT 141.880 45.394 142.220 66.831 ;
 END
 PORT
  LAYER ME4 ;
  RECT 139.688 0.000 140.408 46.394 ;
 END
 PORT
  LAYER ME4 ;
  RECT 145.884 45.394 146.224 66.831 ;
 END
 PORT
  LAYER ME4 ;
  RECT 143.692 0.000 144.412 46.394 ;
 END
 PORT
  LAYER ME4 ;
  RECT 149.888 45.394 150.228 66.831 ;
 END
 PORT
  LAYER ME4 ;
  RECT 147.696 0.000 148.416 46.394 ;
 END
 PORT
  LAYER ME4 ;
  RECT 153.892 45.394 154.232 66.831 ;
 END
 PORT
  LAYER ME4 ;
  RECT 151.700 0.000 152.420 46.394 ;
 END
 PORT
  LAYER ME4 ;
  RECT 157.896 45.394 158.236 66.831 ;
 END
 PORT
  LAYER ME4 ;
  RECT 155.704 0.000 156.424 46.394 ;
 END
 PORT
  LAYER ME4 ;
  RECT 161.900 45.394 162.240 66.831 ;
 END
 PORT
  LAYER ME4 ;
  RECT 159.708 0.000 160.428 46.394 ;
 END
 PORT
  LAYER ME4 ;
  RECT 165.904 45.394 166.244 66.831 ;
 END
 PORT
  LAYER ME4 ;
  RECT 163.712 0.000 164.432 46.394 ;
 END
 PORT
  LAYER ME4 ;
  RECT 169.908 45.394 170.248 66.831 ;
 END
 PORT
  LAYER ME4 ;
  RECT 167.716 0.000 168.436 46.394 ;
 END
 PORT
  LAYER ME4 ;
  RECT 173.912 45.394 174.252 66.831 ;
 END
 PORT
  LAYER ME4 ;
  RECT 171.720 0.000 172.440 46.394 ;
 END
 PORT
  LAYER ME4 ;
  RECT 177.916 45.394 178.256 66.831 ;
 END
 PORT
  LAYER ME4 ;
  RECT 175.724 0.000 176.444 46.394 ;
 END
 PORT
  LAYER ME4 ;
  RECT 185.438 0.000 186.158 66.831 ;
 END
 PORT
  LAYER ME4 ;
  RECT 183.398 0.000 184.118 66.831 ;
 END
 PORT
  LAYER ME4 ;
  RECT 181.278 0.000 181.998 66.831 ;
 END
 PORT
  LAYER ME4 ;
  RECT 180.698 0.000 181.078 66.831 ;
 END
 PORT
  LAYER ME4 ;
  RECT 215.995 47.744 216.335 66.831 ;
 END
 PORT
  LAYER ME4 ;
  RECT 219.999 47.744 220.339 66.831 ;
 END
 PORT
  LAYER ME4 ;
  RECT 224.003 47.744 224.343 66.831 ;
 END
 PORT
  LAYER ME4 ;
  RECT 228.007 47.744 228.347 66.831 ;
 END
 PORT
  LAYER ME4 ;
  RECT 232.011 47.744 232.351 66.831 ;
 END
 PORT
  LAYER ME4 ;
  RECT 236.015 47.744 236.355 66.831 ;
 END
 PORT
  LAYER ME4 ;
  RECT 240.019 47.744 240.359 66.831 ;
 END
 PORT
  LAYER ME4 ;
  RECT 244.023 47.744 244.363 66.831 ;
 END
 PORT
  LAYER ME4 ;
  RECT 248.027 47.744 248.367 66.831 ;
 END
 PORT
  LAYER ME4 ;
  RECT 252.031 47.744 252.371 66.831 ;
 END
 PORT
  LAYER ME4 ;
  RECT 256.035 47.744 256.375 66.831 ;
 END
 PORT
  LAYER ME4 ;
  RECT 260.039 47.744 260.379 66.831 ;
 END
 PORT
  LAYER ME4 ;
  RECT 264.043 47.744 264.383 66.831 ;
 END
 PORT
  LAYER ME4 ;
  RECT 268.047 47.744 268.387 66.831 ;
 END
 PORT
  LAYER ME4 ;
  RECT 272.051 47.744 272.391 66.831 ;
 END
 PORT
  LAYER ME4 ;
  RECT 276.055 47.744 276.395 66.831 ;
 END
 PORT
  LAYER ME4 ;
  RECT 280.059 47.744 280.399 66.831 ;
 END
 PORT
  LAYER ME4 ;
  RECT 284.063 47.744 284.403 66.831 ;
 END
 PORT
  LAYER ME4 ;
  RECT 288.067 47.744 288.407 66.831 ;
 END
 PORT
  LAYER ME4 ;
  RECT 292.071 47.744 292.411 66.831 ;
 END
 PORT
  LAYER ME4 ;
  RECT 296.075 47.744 296.415 66.831 ;
 END
 PORT
  LAYER ME4 ;
  RECT 300.079 47.744 300.419 66.831 ;
 END
 PORT
  LAYER ME4 ;
  RECT 304.083 47.744 304.423 66.831 ;
 END
 PORT
  LAYER ME4 ;
  RECT 308.087 47.744 308.427 66.831 ;
 END
 PORT
  LAYER ME4 ;
  RECT 312.091 47.744 312.431 66.831 ;
 END
 PORT
  LAYER ME4 ;
  RECT 316.095 47.744 316.435 66.831 ;
 END
 PORT
  LAYER ME4 ;
  RECT 320.099 47.744 320.439 66.831 ;
 END
 PORT
  LAYER ME4 ;
  RECT 324.103 47.744 324.443 66.831 ;
 END
 PORT
  LAYER ME4 ;
  RECT 328.107 47.744 328.447 66.831 ;
 END
 PORT
  LAYER ME4 ;
  RECT 332.111 47.744 332.451 66.831 ;
 END
 PORT
  LAYER ME4 ;
  RECT 336.115 47.744 336.455 66.831 ;
 END
 PORT
  LAYER ME4 ;
  RECT 340.119 47.744 340.459 66.831 ;
 END
 PORT
  LAYER ME4 ;
  RECT 344.123 47.744 344.463 66.831 ;
 END
 PORT
  LAYER ME4 ;
  RECT 348.127 47.744 348.467 66.831 ;
 END
 PORT
  LAYER ME4 ;
  RECT 352.131 47.744 352.471 66.831 ;
 END
 PORT
  LAYER ME4 ;
  RECT 356.135 47.744 356.475 66.831 ;
 END
 PORT
  LAYER ME4 ;
  RECT 360.139 47.744 360.479 66.831 ;
 END
 PORT
  LAYER ME4 ;
  RECT 364.143 47.744 364.483 66.831 ;
 END
 PORT
  LAYER ME4 ;
  RECT 368.147 47.744 368.487 66.831 ;
 END
 PORT
  LAYER ME4 ;
  RECT 372.151 47.744 372.491 66.831 ;
 END
 PORT
  LAYER ME4 ;
  RECT 376.155 47.744 376.495 66.831 ;
 END
 PORT
  LAYER ME4 ;
  RECT 380.159 47.744 380.499 66.831 ;
 END
 PORT
  LAYER ME4 ;
  RECT 384.163 47.744 384.503 66.831 ;
 END
 PORT
  LAYER ME4 ;
  RECT 388.167 47.744 388.507 66.831 ;
 END
 PORT
  LAYER ME4 ;
  RECT 3.742 47.744 4.082 66.831 ;
 END
 PORT
  LAYER ME4 ;
  RECT 7.746 47.744 8.086 66.831 ;
 END
 PORT
  LAYER ME4 ;
  RECT 11.750 47.744 12.090 66.831 ;
 END
 PORT
  LAYER ME4 ;
  RECT 15.754 47.744 16.094 66.831 ;
 END
 PORT
  LAYER ME4 ;
  RECT 19.758 47.744 20.098 66.831 ;
 END
 PORT
  LAYER ME4 ;
  RECT 23.762 47.744 24.102 66.831 ;
 END
 PORT
  LAYER ME4 ;
  RECT 27.766 47.744 28.106 66.831 ;
 END
 PORT
  LAYER ME4 ;
  RECT 31.770 47.744 32.110 66.831 ;
 END
 PORT
  LAYER ME4 ;
  RECT 35.774 47.744 36.114 66.831 ;
 END
 PORT
  LAYER ME4 ;
  RECT 39.778 47.744 40.118 66.831 ;
 END
 PORT
  LAYER ME4 ;
  RECT 43.782 47.744 44.122 66.831 ;
 END
 PORT
  LAYER ME4 ;
  RECT 47.786 47.744 48.126 66.831 ;
 END
 PORT
  LAYER ME4 ;
  RECT 51.790 47.744 52.130 66.831 ;
 END
 PORT
  LAYER ME4 ;
  RECT 55.794 47.744 56.134 66.831 ;
 END
 PORT
  LAYER ME4 ;
  RECT 59.798 47.744 60.138 66.831 ;
 END
 PORT
  LAYER ME4 ;
  RECT 63.802 47.744 64.142 66.831 ;
 END
 PORT
  LAYER ME4 ;
  RECT 67.806 47.744 68.146 66.831 ;
 END
 PORT
  LAYER ME4 ;
  RECT 71.810 47.744 72.150 66.831 ;
 END
 PORT
  LAYER ME4 ;
  RECT 75.814 47.744 76.154 66.831 ;
 END
 PORT
  LAYER ME4 ;
  RECT 79.818 47.744 80.158 66.831 ;
 END
 PORT
  LAYER ME4 ;
  RECT 83.822 47.744 84.162 66.831 ;
 END
 PORT
  LAYER ME4 ;
  RECT 87.826 47.744 88.166 66.831 ;
 END
 PORT
  LAYER ME4 ;
  RECT 91.830 47.744 92.170 66.831 ;
 END
 PORT
  LAYER ME4 ;
  RECT 95.834 47.744 96.174 66.831 ;
 END
 PORT
  LAYER ME4 ;
  RECT 99.838 47.744 100.178 66.831 ;
 END
 PORT
  LAYER ME4 ;
  RECT 103.842 47.744 104.182 66.831 ;
 END
 PORT
  LAYER ME4 ;
  RECT 107.846 47.744 108.186 66.831 ;
 END
 PORT
  LAYER ME4 ;
  RECT 111.850 47.744 112.190 66.831 ;
 END
 PORT
  LAYER ME4 ;
  RECT 115.854 47.744 116.194 66.831 ;
 END
 PORT
  LAYER ME4 ;
  RECT 119.858 47.744 120.198 66.831 ;
 END
 PORT
  LAYER ME4 ;
  RECT 123.862 47.744 124.202 66.831 ;
 END
 PORT
  LAYER ME4 ;
  RECT 127.866 47.744 128.206 66.831 ;
 END
 PORT
  LAYER ME4 ;
  RECT 131.870 47.744 132.210 66.831 ;
 END
 PORT
  LAYER ME4 ;
  RECT 135.874 47.744 136.214 66.831 ;
 END
 PORT
  LAYER ME4 ;
  RECT 139.878 47.744 140.218 66.831 ;
 END
 PORT
  LAYER ME4 ;
  RECT 143.882 47.744 144.222 66.831 ;
 END
 PORT
  LAYER ME4 ;
  RECT 147.886 47.744 148.226 66.831 ;
 END
 PORT
  LAYER ME4 ;
  RECT 151.890 47.744 152.230 66.831 ;
 END
 PORT
  LAYER ME4 ;
  RECT 155.894 47.744 156.234 66.831 ;
 END
 PORT
  LAYER ME4 ;
  RECT 159.898 47.744 160.238 66.831 ;
 END
 PORT
  LAYER ME4 ;
  RECT 163.902 47.744 164.242 66.831 ;
 END
 PORT
  LAYER ME4 ;
  RECT 167.906 47.744 168.246 66.831 ;
 END
 PORT
  LAYER ME4 ;
  RECT 171.910 47.744 172.250 66.831 ;
 END
 PORT
  LAYER ME4 ;
  RECT 175.914 47.744 176.254 66.831 ;
 END
END VCC
PIN DI43
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 177.206 0.000 177.526 0.600 ;
  LAYER ME3 ;
  RECT 177.206 0.000 177.526 0.600 ;
  LAYER ME2 ;
  RECT 177.206 0.000 177.526 0.600 ;
  LAYER ME1 ;
  RECT 177.206 0.000 177.526 0.600 ;
 END
 ANTENNAPARTIALMETALAREA                  1.058 LAYER ME2 ;
 ANTENNAGATEAREA                          0.072 LAYER ME2 ;
 ANTENNAGATEAREA                          0.072 LAYER ME3 ;
 ANTENNAGATEAREA                          0.072 LAYER ME4 ;
 ANTENNADIFFAREA                          0.160 LAYER ME2 ;
 ANTENNADIFFAREA                          0.160 LAYER ME3 ;
 ANTENNADIFFAREA                          0.160 LAYER ME4 ;
 ANTENNAMAXAREACAR                       21.782 LAYER ME2 ;
 ANTENNAMAXAREACAR                       24.449 LAYER ME3 ;
 ANTENNAMAXAREACAR                       27.116 LAYER ME4 ;
END DI43
PIN DO43
  DIRECTION OUTPUT ;
 PORT
  LAYER ME4 ;
  RECT 176.644 0.000 176.964 0.600 ;
  LAYER ME3 ;
  RECT 176.644 0.000 176.964 0.600 ;
  LAYER ME2 ;
  RECT 176.644 0.000 176.964 0.600 ;
  LAYER ME1 ;
  RECT 176.644 0.000 176.964 0.600 ;
 END
 ANTENNAPARTIALMETALAREA                  5.273 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME3 ;
 ANTENNADIFFAREA                          1.293 LAYER ME4 ;
END DO43
PIN DI42
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 173.202 0.000 173.522 0.600 ;
  LAYER ME3 ;
  RECT 173.202 0.000 173.522 0.600 ;
  LAYER ME2 ;
  RECT 173.202 0.000 173.522 0.600 ;
  LAYER ME1 ;
  RECT 173.202 0.000 173.522 0.600 ;
 END
 ANTENNAPARTIALMETALAREA                  1.058 LAYER ME2 ;
 ANTENNAGATEAREA                          0.072 LAYER ME2 ;
 ANTENNAGATEAREA                          0.072 LAYER ME3 ;
 ANTENNAGATEAREA                          0.072 LAYER ME4 ;
 ANTENNADIFFAREA                          0.160 LAYER ME2 ;
 ANTENNADIFFAREA                          0.160 LAYER ME3 ;
 ANTENNADIFFAREA                          0.160 LAYER ME4 ;
 ANTENNAMAXAREACAR                       21.782 LAYER ME2 ;
 ANTENNAMAXAREACAR                       24.449 LAYER ME3 ;
 ANTENNAMAXAREACAR                       27.116 LAYER ME4 ;
END DI42
PIN DO42
  DIRECTION OUTPUT ;
 PORT
  LAYER ME4 ;
  RECT 172.640 0.000 172.960 0.600 ;
  LAYER ME3 ;
  RECT 172.640 0.000 172.960 0.600 ;
  LAYER ME2 ;
  RECT 172.640 0.000 172.960 0.600 ;
  LAYER ME1 ;
  RECT 172.640 0.000 172.960 0.600 ;
 END
 ANTENNAPARTIALMETALAREA                  5.273 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME3 ;
 ANTENNADIFFAREA                          1.293 LAYER ME4 ;
END DO42
PIN DI41
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 169.198 0.000 169.518 0.600 ;
  LAYER ME3 ;
  RECT 169.198 0.000 169.518 0.600 ;
  LAYER ME2 ;
  RECT 169.198 0.000 169.518 0.600 ;
  LAYER ME1 ;
  RECT 169.198 0.000 169.518 0.600 ;
 END
 ANTENNAPARTIALMETALAREA                  1.058 LAYER ME2 ;
 ANTENNAGATEAREA                          0.072 LAYER ME2 ;
 ANTENNAGATEAREA                          0.072 LAYER ME3 ;
 ANTENNAGATEAREA                          0.072 LAYER ME4 ;
 ANTENNADIFFAREA                          0.160 LAYER ME2 ;
 ANTENNADIFFAREA                          0.160 LAYER ME3 ;
 ANTENNADIFFAREA                          0.160 LAYER ME4 ;
 ANTENNAMAXAREACAR                       21.782 LAYER ME2 ;
 ANTENNAMAXAREACAR                       24.449 LAYER ME3 ;
 ANTENNAMAXAREACAR                       27.116 LAYER ME4 ;
END DI41
PIN DO41
  DIRECTION OUTPUT ;
 PORT
  LAYER ME4 ;
  RECT 168.636 0.000 168.956 0.600 ;
  LAYER ME3 ;
  RECT 168.636 0.000 168.956 0.600 ;
  LAYER ME2 ;
  RECT 168.636 0.000 168.956 0.600 ;
  LAYER ME1 ;
  RECT 168.636 0.000 168.956 0.600 ;
 END
 ANTENNAPARTIALMETALAREA                  5.273 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME3 ;
 ANTENNADIFFAREA                          1.293 LAYER ME4 ;
END DO41
PIN DI40
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 165.194 0.000 165.514 0.600 ;
  LAYER ME3 ;
  RECT 165.194 0.000 165.514 0.600 ;
  LAYER ME2 ;
  RECT 165.194 0.000 165.514 0.600 ;
  LAYER ME1 ;
  RECT 165.194 0.000 165.514 0.600 ;
 END
 ANTENNAPARTIALMETALAREA                  1.058 LAYER ME2 ;
 ANTENNAGATEAREA                          0.072 LAYER ME2 ;
 ANTENNAGATEAREA                          0.072 LAYER ME3 ;
 ANTENNAGATEAREA                          0.072 LAYER ME4 ;
 ANTENNADIFFAREA                          0.160 LAYER ME2 ;
 ANTENNADIFFAREA                          0.160 LAYER ME3 ;
 ANTENNADIFFAREA                          0.160 LAYER ME4 ;
 ANTENNAMAXAREACAR                       21.782 LAYER ME2 ;
 ANTENNAMAXAREACAR                       24.449 LAYER ME3 ;
 ANTENNAMAXAREACAR                       27.116 LAYER ME4 ;
END DI40
PIN DO40
  DIRECTION OUTPUT ;
 PORT
  LAYER ME4 ;
  RECT 164.632 0.000 164.952 0.600 ;
  LAYER ME3 ;
  RECT 164.632 0.000 164.952 0.600 ;
  LAYER ME2 ;
  RECT 164.632 0.000 164.952 0.600 ;
  LAYER ME1 ;
  RECT 164.632 0.000 164.952 0.600 ;
 END
 ANTENNAPARTIALMETALAREA                  5.273 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME3 ;
 ANTENNADIFFAREA                          1.293 LAYER ME4 ;
END DO40
PIN DI39
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 161.190 0.000 161.510 0.600 ;
  LAYER ME3 ;
  RECT 161.190 0.000 161.510 0.600 ;
  LAYER ME2 ;
  RECT 161.190 0.000 161.510 0.600 ;
  LAYER ME1 ;
  RECT 161.190 0.000 161.510 0.600 ;
 END
 ANTENNAPARTIALMETALAREA                  1.058 LAYER ME2 ;
 ANTENNAGATEAREA                          0.072 LAYER ME2 ;
 ANTENNAGATEAREA                          0.072 LAYER ME3 ;
 ANTENNAGATEAREA                          0.072 LAYER ME4 ;
 ANTENNADIFFAREA                          0.160 LAYER ME2 ;
 ANTENNADIFFAREA                          0.160 LAYER ME3 ;
 ANTENNADIFFAREA                          0.160 LAYER ME4 ;
 ANTENNAMAXAREACAR                       21.782 LAYER ME2 ;
 ANTENNAMAXAREACAR                       24.449 LAYER ME3 ;
 ANTENNAMAXAREACAR                       27.116 LAYER ME4 ;
END DI39
PIN DO39
  DIRECTION OUTPUT ;
 PORT
  LAYER ME4 ;
  RECT 160.628 0.000 160.948 0.600 ;
  LAYER ME3 ;
  RECT 160.628 0.000 160.948 0.600 ;
  LAYER ME2 ;
  RECT 160.628 0.000 160.948 0.600 ;
  LAYER ME1 ;
  RECT 160.628 0.000 160.948 0.600 ;
 END
 ANTENNAPARTIALMETALAREA                  5.273 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME3 ;
 ANTENNADIFFAREA                          1.293 LAYER ME4 ;
END DO39
PIN DI38
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 157.186 0.000 157.506 0.600 ;
  LAYER ME3 ;
  RECT 157.186 0.000 157.506 0.600 ;
  LAYER ME2 ;
  RECT 157.186 0.000 157.506 0.600 ;
  LAYER ME1 ;
  RECT 157.186 0.000 157.506 0.600 ;
 END
 ANTENNAPARTIALMETALAREA                  1.058 LAYER ME2 ;
 ANTENNAGATEAREA                          0.072 LAYER ME2 ;
 ANTENNAGATEAREA                          0.072 LAYER ME3 ;
 ANTENNAGATEAREA                          0.072 LAYER ME4 ;
 ANTENNADIFFAREA                          0.160 LAYER ME2 ;
 ANTENNADIFFAREA                          0.160 LAYER ME3 ;
 ANTENNADIFFAREA                          0.160 LAYER ME4 ;
 ANTENNAMAXAREACAR                       21.782 LAYER ME2 ;
 ANTENNAMAXAREACAR                       24.449 LAYER ME3 ;
 ANTENNAMAXAREACAR                       27.116 LAYER ME4 ;
END DI38
PIN DO38
  DIRECTION OUTPUT ;
 PORT
  LAYER ME4 ;
  RECT 156.624 0.000 156.944 0.600 ;
  LAYER ME3 ;
  RECT 156.624 0.000 156.944 0.600 ;
  LAYER ME2 ;
  RECT 156.624 0.000 156.944 0.600 ;
  LAYER ME1 ;
  RECT 156.624 0.000 156.944 0.600 ;
 END
 ANTENNAPARTIALMETALAREA                  5.273 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME3 ;
 ANTENNADIFFAREA                          1.293 LAYER ME4 ;
END DO38
PIN DI37
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 153.182 0.000 153.502 0.600 ;
  LAYER ME3 ;
  RECT 153.182 0.000 153.502 0.600 ;
  LAYER ME2 ;
  RECT 153.182 0.000 153.502 0.600 ;
  LAYER ME1 ;
  RECT 153.182 0.000 153.502 0.600 ;
 END
 ANTENNAPARTIALMETALAREA                  1.058 LAYER ME2 ;
 ANTENNAGATEAREA                          0.072 LAYER ME2 ;
 ANTENNAGATEAREA                          0.072 LAYER ME3 ;
 ANTENNAGATEAREA                          0.072 LAYER ME4 ;
 ANTENNADIFFAREA                          0.160 LAYER ME2 ;
 ANTENNADIFFAREA                          0.160 LAYER ME3 ;
 ANTENNADIFFAREA                          0.160 LAYER ME4 ;
 ANTENNAMAXAREACAR                       21.782 LAYER ME2 ;
 ANTENNAMAXAREACAR                       24.449 LAYER ME3 ;
 ANTENNAMAXAREACAR                       27.116 LAYER ME4 ;
END DI37
PIN DO37
  DIRECTION OUTPUT ;
 PORT
  LAYER ME4 ;
  RECT 152.620 0.000 152.940 0.600 ;
  LAYER ME3 ;
  RECT 152.620 0.000 152.940 0.600 ;
  LAYER ME2 ;
  RECT 152.620 0.000 152.940 0.600 ;
  LAYER ME1 ;
  RECT 152.620 0.000 152.940 0.600 ;
 END
 ANTENNAPARTIALMETALAREA                  5.273 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME3 ;
 ANTENNADIFFAREA                          1.293 LAYER ME4 ;
END DO37
PIN DI36
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 149.178 0.000 149.498 0.600 ;
  LAYER ME3 ;
  RECT 149.178 0.000 149.498 0.600 ;
  LAYER ME2 ;
  RECT 149.178 0.000 149.498 0.600 ;
  LAYER ME1 ;
  RECT 149.178 0.000 149.498 0.600 ;
 END
 ANTENNAPARTIALMETALAREA                  1.058 LAYER ME2 ;
 ANTENNAGATEAREA                          0.072 LAYER ME2 ;
 ANTENNAGATEAREA                          0.072 LAYER ME3 ;
 ANTENNAGATEAREA                          0.072 LAYER ME4 ;
 ANTENNADIFFAREA                          0.160 LAYER ME2 ;
 ANTENNADIFFAREA                          0.160 LAYER ME3 ;
 ANTENNADIFFAREA                          0.160 LAYER ME4 ;
 ANTENNAMAXAREACAR                       21.782 LAYER ME2 ;
 ANTENNAMAXAREACAR                       24.449 LAYER ME3 ;
 ANTENNAMAXAREACAR                       27.116 LAYER ME4 ;
END DI36
PIN DO36
  DIRECTION OUTPUT ;
 PORT
  LAYER ME4 ;
  RECT 148.616 0.000 148.936 0.600 ;
  LAYER ME3 ;
  RECT 148.616 0.000 148.936 0.600 ;
  LAYER ME2 ;
  RECT 148.616 0.000 148.936 0.600 ;
  LAYER ME1 ;
  RECT 148.616 0.000 148.936 0.600 ;
 END
 ANTENNAPARTIALMETALAREA                  5.273 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME3 ;
 ANTENNADIFFAREA                          1.293 LAYER ME4 ;
END DO36
PIN DI35
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 145.174 0.000 145.494 0.600 ;
  LAYER ME3 ;
  RECT 145.174 0.000 145.494 0.600 ;
  LAYER ME2 ;
  RECT 145.174 0.000 145.494 0.600 ;
  LAYER ME1 ;
  RECT 145.174 0.000 145.494 0.600 ;
 END
 ANTENNAPARTIALMETALAREA                  1.058 LAYER ME2 ;
 ANTENNAGATEAREA                          0.072 LAYER ME2 ;
 ANTENNAGATEAREA                          0.072 LAYER ME3 ;
 ANTENNAGATEAREA                          0.072 LAYER ME4 ;
 ANTENNADIFFAREA                          0.160 LAYER ME2 ;
 ANTENNADIFFAREA                          0.160 LAYER ME3 ;
 ANTENNADIFFAREA                          0.160 LAYER ME4 ;
 ANTENNAMAXAREACAR                       21.782 LAYER ME2 ;
 ANTENNAMAXAREACAR                       24.449 LAYER ME3 ;
 ANTENNAMAXAREACAR                       27.116 LAYER ME4 ;
END DI35
PIN DO35
  DIRECTION OUTPUT ;
 PORT
  LAYER ME4 ;
  RECT 144.612 0.000 144.932 0.600 ;
  LAYER ME3 ;
  RECT 144.612 0.000 144.932 0.600 ;
  LAYER ME2 ;
  RECT 144.612 0.000 144.932 0.600 ;
  LAYER ME1 ;
  RECT 144.612 0.000 144.932 0.600 ;
 END
 ANTENNAPARTIALMETALAREA                  5.273 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME3 ;
 ANTENNADIFFAREA                          1.293 LAYER ME4 ;
END DO35
PIN DI34
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 141.170 0.000 141.490 0.600 ;
  LAYER ME3 ;
  RECT 141.170 0.000 141.490 0.600 ;
  LAYER ME2 ;
  RECT 141.170 0.000 141.490 0.600 ;
  LAYER ME1 ;
  RECT 141.170 0.000 141.490 0.600 ;
 END
 ANTENNAPARTIALMETALAREA                  1.058 LAYER ME2 ;
 ANTENNAGATEAREA                          0.072 LAYER ME2 ;
 ANTENNAGATEAREA                          0.072 LAYER ME3 ;
 ANTENNAGATEAREA                          0.072 LAYER ME4 ;
 ANTENNADIFFAREA                          0.160 LAYER ME2 ;
 ANTENNADIFFAREA                          0.160 LAYER ME3 ;
 ANTENNADIFFAREA                          0.160 LAYER ME4 ;
 ANTENNAMAXAREACAR                       21.782 LAYER ME2 ;
 ANTENNAMAXAREACAR                       24.449 LAYER ME3 ;
 ANTENNAMAXAREACAR                       27.116 LAYER ME4 ;
END DI34
PIN DO34
  DIRECTION OUTPUT ;
 PORT
  LAYER ME4 ;
  RECT 140.608 0.000 140.928 0.600 ;
  LAYER ME3 ;
  RECT 140.608 0.000 140.928 0.600 ;
  LAYER ME2 ;
  RECT 140.608 0.000 140.928 0.600 ;
  LAYER ME1 ;
  RECT 140.608 0.000 140.928 0.600 ;
 END
 ANTENNAPARTIALMETALAREA                  5.273 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME3 ;
 ANTENNADIFFAREA                          1.293 LAYER ME4 ;
END DO34
PIN DI33
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 136.604 0.000 136.924 0.600 ;
  LAYER ME3 ;
  RECT 136.604 0.000 136.924 0.600 ;
  LAYER ME2 ;
  RECT 136.604 0.000 136.924 0.600 ;
  LAYER ME1 ;
  RECT 136.604 0.000 136.924 0.600 ;
 END
 ANTENNAPARTIALMETALAREA                  0.346 LAYER ME1 ;
 ANTENNAPARTIALMETALAREA                  1.466 LAYER ME2 ;
 ANTENNAPARTIALMETALAREA                  0.508 LAYER ME3 ;
 ANTENNAGATEAREA                          0.072 LAYER ME3 ;
 ANTENNAGATEAREA                          0.072 LAYER ME4 ;
 ANTENNADIFFAREA                          0.218 LAYER ME1 ;
 ANTENNADIFFAREA                          0.218 LAYER ME2 ;
 ANTENNADIFFAREA                          0.218 LAYER ME3 ;
 ANTENNADIFFAREA                          0.218 LAYER ME4 ;
 ANTENNAMAXAREACAR                       17.267 LAYER ME3 ;
 ANTENNAMAXAREACAR                       19.933 LAYER ME4 ;
END DI33
PIN DO33
  DIRECTION OUTPUT ;
 PORT
  LAYER ME4 ;
  RECT 137.166 0.000 137.486 0.600 ;
  LAYER ME3 ;
  RECT 137.166 0.000 137.486 0.600 ;
  LAYER ME2 ;
  RECT 137.166 0.000 137.486 0.600 ;
  LAYER ME1 ;
  RECT 137.166 0.000 137.486 0.600 ;
 END
 ANTENNAPARTIALMETALAREA                  5.602 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME3 ;
 ANTENNADIFFAREA                          1.293 LAYER ME4 ;
END DO33
PIN WEB3
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 135.164 0.000 135.484 0.600 ;
  LAYER ME3 ;
  RECT 135.164 0.000 135.484 0.600 ;
  LAYER ME2 ;
  RECT 135.164 0.000 135.484 0.600 ;
  LAYER ME1 ;
  RECT 135.164 0.000 135.484 0.600 ;
 END
 ANTENNAPARTIALMETALAREA                  1.036 LAYER ME2 ;
 ANTENNAGATEAREA                          0.288 LAYER ME2 ;
 ANTENNAGATEAREA                          0.288 LAYER ME3 ;
 ANTENNAGATEAREA                          0.288 LAYER ME4 ;
 ANTENNADIFFAREA                          0.206 LAYER ME2 ;
 ANTENNADIFFAREA                          0.206 LAYER ME3 ;
 ANTENNADIFFAREA                          0.206 LAYER ME4 ;
 ANTENNAMAXAREACAR                        5.844 LAYER ME2 ;
 ANTENNAMAXAREACAR                        6.511 LAYER ME3 ;
 ANTENNAMAXAREACAR                        7.178 LAYER ME4 ;
END WEB3
PIN DI32
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 133.162 0.000 133.482 0.600 ;
  LAYER ME3 ;
  RECT 133.162 0.000 133.482 0.600 ;
  LAYER ME2 ;
  RECT 133.162 0.000 133.482 0.600 ;
  LAYER ME1 ;
  RECT 133.162 0.000 133.482 0.600 ;
 END
 ANTENNAPARTIALMETALAREA                  1.058 LAYER ME2 ;
 ANTENNAGATEAREA                          0.072 LAYER ME2 ;
 ANTENNAGATEAREA                          0.072 LAYER ME3 ;
 ANTENNAGATEAREA                          0.072 LAYER ME4 ;
 ANTENNADIFFAREA                          0.160 LAYER ME2 ;
 ANTENNADIFFAREA                          0.160 LAYER ME3 ;
 ANTENNADIFFAREA                          0.160 LAYER ME4 ;
 ANTENNAMAXAREACAR                       21.782 LAYER ME2 ;
 ANTENNAMAXAREACAR                       24.449 LAYER ME3 ;
 ANTENNAMAXAREACAR                       27.116 LAYER ME4 ;
END DI32
PIN DO32
  DIRECTION OUTPUT ;
 PORT
  LAYER ME4 ;
  RECT 132.600 0.000 132.920 0.600 ;
  LAYER ME3 ;
  RECT 132.600 0.000 132.920 0.600 ;
  LAYER ME2 ;
  RECT 132.600 0.000 132.920 0.600 ;
  LAYER ME1 ;
  RECT 132.600 0.000 132.920 0.600 ;
 END
 ANTENNAPARTIALMETALAREA                  5.273 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME3 ;
 ANTENNADIFFAREA                          1.293 LAYER ME4 ;
END DO32
PIN DI31
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 129.158 0.000 129.478 0.600 ;
  LAYER ME3 ;
  RECT 129.158 0.000 129.478 0.600 ;
  LAYER ME2 ;
  RECT 129.158 0.000 129.478 0.600 ;
  LAYER ME1 ;
  RECT 129.158 0.000 129.478 0.600 ;
 END
 ANTENNAPARTIALMETALAREA                  1.058 LAYER ME2 ;
 ANTENNAGATEAREA                          0.072 LAYER ME2 ;
 ANTENNAGATEAREA                          0.072 LAYER ME3 ;
 ANTENNAGATEAREA                          0.072 LAYER ME4 ;
 ANTENNADIFFAREA                          0.160 LAYER ME2 ;
 ANTENNADIFFAREA                          0.160 LAYER ME3 ;
 ANTENNADIFFAREA                          0.160 LAYER ME4 ;
 ANTENNAMAXAREACAR                       21.782 LAYER ME2 ;
 ANTENNAMAXAREACAR                       24.449 LAYER ME3 ;
 ANTENNAMAXAREACAR                       27.116 LAYER ME4 ;
END DI31
PIN DO31
  DIRECTION OUTPUT ;
 PORT
  LAYER ME4 ;
  RECT 128.596 0.000 128.916 0.600 ;
  LAYER ME3 ;
  RECT 128.596 0.000 128.916 0.600 ;
  LAYER ME2 ;
  RECT 128.596 0.000 128.916 0.600 ;
  LAYER ME1 ;
  RECT 128.596 0.000 128.916 0.600 ;
 END
 ANTENNAPARTIALMETALAREA                  5.273 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME3 ;
 ANTENNADIFFAREA                          1.293 LAYER ME4 ;
END DO31
PIN DI30
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 125.154 0.000 125.474 0.600 ;
  LAYER ME3 ;
  RECT 125.154 0.000 125.474 0.600 ;
  LAYER ME2 ;
  RECT 125.154 0.000 125.474 0.600 ;
  LAYER ME1 ;
  RECT 125.154 0.000 125.474 0.600 ;
 END
 ANTENNAPARTIALMETALAREA                  1.058 LAYER ME2 ;
 ANTENNAGATEAREA                          0.072 LAYER ME2 ;
 ANTENNAGATEAREA                          0.072 LAYER ME3 ;
 ANTENNAGATEAREA                          0.072 LAYER ME4 ;
 ANTENNADIFFAREA                          0.160 LAYER ME2 ;
 ANTENNADIFFAREA                          0.160 LAYER ME3 ;
 ANTENNADIFFAREA                          0.160 LAYER ME4 ;
 ANTENNAMAXAREACAR                       21.782 LAYER ME2 ;
 ANTENNAMAXAREACAR                       24.449 LAYER ME3 ;
 ANTENNAMAXAREACAR                       27.116 LAYER ME4 ;
END DI30
PIN DO30
  DIRECTION OUTPUT ;
 PORT
  LAYER ME4 ;
  RECT 124.592 0.000 124.912 0.600 ;
  LAYER ME3 ;
  RECT 124.592 0.000 124.912 0.600 ;
  LAYER ME2 ;
  RECT 124.592 0.000 124.912 0.600 ;
  LAYER ME1 ;
  RECT 124.592 0.000 124.912 0.600 ;
 END
 ANTENNAPARTIALMETALAREA                  5.273 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME3 ;
 ANTENNADIFFAREA                          1.293 LAYER ME4 ;
END DO30
PIN DI29
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 121.150 0.000 121.470 0.600 ;
  LAYER ME3 ;
  RECT 121.150 0.000 121.470 0.600 ;
  LAYER ME2 ;
  RECT 121.150 0.000 121.470 0.600 ;
  LAYER ME1 ;
  RECT 121.150 0.000 121.470 0.600 ;
 END
 ANTENNAPARTIALMETALAREA                  1.058 LAYER ME2 ;
 ANTENNAGATEAREA                          0.072 LAYER ME2 ;
 ANTENNAGATEAREA                          0.072 LAYER ME3 ;
 ANTENNAGATEAREA                          0.072 LAYER ME4 ;
 ANTENNADIFFAREA                          0.160 LAYER ME2 ;
 ANTENNADIFFAREA                          0.160 LAYER ME3 ;
 ANTENNADIFFAREA                          0.160 LAYER ME4 ;
 ANTENNAMAXAREACAR                       21.782 LAYER ME2 ;
 ANTENNAMAXAREACAR                       24.449 LAYER ME3 ;
 ANTENNAMAXAREACAR                       27.116 LAYER ME4 ;
END DI29
PIN DO29
  DIRECTION OUTPUT ;
 PORT
  LAYER ME4 ;
  RECT 120.588 0.000 120.908 0.600 ;
  LAYER ME3 ;
  RECT 120.588 0.000 120.908 0.600 ;
  LAYER ME2 ;
  RECT 120.588 0.000 120.908 0.600 ;
  LAYER ME1 ;
  RECT 120.588 0.000 120.908 0.600 ;
 END
 ANTENNAPARTIALMETALAREA                  5.273 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME3 ;
 ANTENNADIFFAREA                          1.293 LAYER ME4 ;
END DO29
PIN DI28
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 117.146 0.000 117.466 0.600 ;
  LAYER ME3 ;
  RECT 117.146 0.000 117.466 0.600 ;
  LAYER ME2 ;
  RECT 117.146 0.000 117.466 0.600 ;
  LAYER ME1 ;
  RECT 117.146 0.000 117.466 0.600 ;
 END
 ANTENNAPARTIALMETALAREA                  1.058 LAYER ME2 ;
 ANTENNAGATEAREA                          0.072 LAYER ME2 ;
 ANTENNAGATEAREA                          0.072 LAYER ME3 ;
 ANTENNAGATEAREA                          0.072 LAYER ME4 ;
 ANTENNADIFFAREA                          0.160 LAYER ME2 ;
 ANTENNADIFFAREA                          0.160 LAYER ME3 ;
 ANTENNADIFFAREA                          0.160 LAYER ME4 ;
 ANTENNAMAXAREACAR                       21.782 LAYER ME2 ;
 ANTENNAMAXAREACAR                       24.449 LAYER ME3 ;
 ANTENNAMAXAREACAR                       27.116 LAYER ME4 ;
END DI28
PIN DO28
  DIRECTION OUTPUT ;
 PORT
  LAYER ME4 ;
  RECT 116.584 0.000 116.904 0.600 ;
  LAYER ME3 ;
  RECT 116.584 0.000 116.904 0.600 ;
  LAYER ME2 ;
  RECT 116.584 0.000 116.904 0.600 ;
  LAYER ME1 ;
  RECT 116.584 0.000 116.904 0.600 ;
 END
 ANTENNAPARTIALMETALAREA                  5.273 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME3 ;
 ANTENNADIFFAREA                          1.293 LAYER ME4 ;
END DO28
PIN DI27
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 113.142 0.000 113.462 0.600 ;
  LAYER ME3 ;
  RECT 113.142 0.000 113.462 0.600 ;
  LAYER ME2 ;
  RECT 113.142 0.000 113.462 0.600 ;
  LAYER ME1 ;
  RECT 113.142 0.000 113.462 0.600 ;
 END
 ANTENNAPARTIALMETALAREA                  1.058 LAYER ME2 ;
 ANTENNAGATEAREA                          0.072 LAYER ME2 ;
 ANTENNAGATEAREA                          0.072 LAYER ME3 ;
 ANTENNAGATEAREA                          0.072 LAYER ME4 ;
 ANTENNADIFFAREA                          0.160 LAYER ME2 ;
 ANTENNADIFFAREA                          0.160 LAYER ME3 ;
 ANTENNADIFFAREA                          0.160 LAYER ME4 ;
 ANTENNAMAXAREACAR                       21.782 LAYER ME2 ;
 ANTENNAMAXAREACAR                       24.449 LAYER ME3 ;
 ANTENNAMAXAREACAR                       27.116 LAYER ME4 ;
END DI27
PIN DO27
  DIRECTION OUTPUT ;
 PORT
  LAYER ME4 ;
  RECT 112.580 0.000 112.900 0.600 ;
  LAYER ME3 ;
  RECT 112.580 0.000 112.900 0.600 ;
  LAYER ME2 ;
  RECT 112.580 0.000 112.900 0.600 ;
  LAYER ME1 ;
  RECT 112.580 0.000 112.900 0.600 ;
 END
 ANTENNAPARTIALMETALAREA                  5.273 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME3 ;
 ANTENNADIFFAREA                          1.293 LAYER ME4 ;
END DO27
PIN DI26
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 109.138 0.000 109.458 0.600 ;
  LAYER ME3 ;
  RECT 109.138 0.000 109.458 0.600 ;
  LAYER ME2 ;
  RECT 109.138 0.000 109.458 0.600 ;
  LAYER ME1 ;
  RECT 109.138 0.000 109.458 0.600 ;
 END
 ANTENNAPARTIALMETALAREA                  1.058 LAYER ME2 ;
 ANTENNAGATEAREA                          0.072 LAYER ME2 ;
 ANTENNAGATEAREA                          0.072 LAYER ME3 ;
 ANTENNAGATEAREA                          0.072 LAYER ME4 ;
 ANTENNADIFFAREA                          0.160 LAYER ME2 ;
 ANTENNADIFFAREA                          0.160 LAYER ME3 ;
 ANTENNADIFFAREA                          0.160 LAYER ME4 ;
 ANTENNAMAXAREACAR                       21.782 LAYER ME2 ;
 ANTENNAMAXAREACAR                       24.449 LAYER ME3 ;
 ANTENNAMAXAREACAR                       27.116 LAYER ME4 ;
END DI26
PIN DO26
  DIRECTION OUTPUT ;
 PORT
  LAYER ME4 ;
  RECT 108.576 0.000 108.896 0.600 ;
  LAYER ME3 ;
  RECT 108.576 0.000 108.896 0.600 ;
  LAYER ME2 ;
  RECT 108.576 0.000 108.896 0.600 ;
  LAYER ME1 ;
  RECT 108.576 0.000 108.896 0.600 ;
 END
 ANTENNAPARTIALMETALAREA                  5.273 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME3 ;
 ANTENNADIFFAREA                          1.293 LAYER ME4 ;
END DO26
PIN DI25
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 105.134 0.000 105.454 0.600 ;
  LAYER ME3 ;
  RECT 105.134 0.000 105.454 0.600 ;
  LAYER ME2 ;
  RECT 105.134 0.000 105.454 0.600 ;
  LAYER ME1 ;
  RECT 105.134 0.000 105.454 0.600 ;
 END
 ANTENNAPARTIALMETALAREA                  1.058 LAYER ME2 ;
 ANTENNAGATEAREA                          0.072 LAYER ME2 ;
 ANTENNAGATEAREA                          0.072 LAYER ME3 ;
 ANTENNAGATEAREA                          0.072 LAYER ME4 ;
 ANTENNADIFFAREA                          0.160 LAYER ME2 ;
 ANTENNADIFFAREA                          0.160 LAYER ME3 ;
 ANTENNADIFFAREA                          0.160 LAYER ME4 ;
 ANTENNAMAXAREACAR                       21.782 LAYER ME2 ;
 ANTENNAMAXAREACAR                       24.449 LAYER ME3 ;
 ANTENNAMAXAREACAR                       27.116 LAYER ME4 ;
END DI25
PIN DO25
  DIRECTION OUTPUT ;
 PORT
  LAYER ME4 ;
  RECT 104.572 0.000 104.892 0.600 ;
  LAYER ME3 ;
  RECT 104.572 0.000 104.892 0.600 ;
  LAYER ME2 ;
  RECT 104.572 0.000 104.892 0.600 ;
  LAYER ME1 ;
  RECT 104.572 0.000 104.892 0.600 ;
 END
 ANTENNAPARTIALMETALAREA                  5.273 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME3 ;
 ANTENNADIFFAREA                          1.293 LAYER ME4 ;
END DO25
PIN DI24
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 101.130 0.000 101.450 0.600 ;
  LAYER ME3 ;
  RECT 101.130 0.000 101.450 0.600 ;
  LAYER ME2 ;
  RECT 101.130 0.000 101.450 0.600 ;
  LAYER ME1 ;
  RECT 101.130 0.000 101.450 0.600 ;
 END
 ANTENNAPARTIALMETALAREA                  1.058 LAYER ME2 ;
 ANTENNAGATEAREA                          0.072 LAYER ME2 ;
 ANTENNAGATEAREA                          0.072 LAYER ME3 ;
 ANTENNAGATEAREA                          0.072 LAYER ME4 ;
 ANTENNADIFFAREA                          0.160 LAYER ME2 ;
 ANTENNADIFFAREA                          0.160 LAYER ME3 ;
 ANTENNADIFFAREA                          0.160 LAYER ME4 ;
 ANTENNAMAXAREACAR                       21.782 LAYER ME2 ;
 ANTENNAMAXAREACAR                       24.449 LAYER ME3 ;
 ANTENNAMAXAREACAR                       27.116 LAYER ME4 ;
END DI24
PIN DO24
  DIRECTION OUTPUT ;
 PORT
  LAYER ME4 ;
  RECT 100.568 0.000 100.888 0.600 ;
  LAYER ME3 ;
  RECT 100.568 0.000 100.888 0.600 ;
  LAYER ME2 ;
  RECT 100.568 0.000 100.888 0.600 ;
  LAYER ME1 ;
  RECT 100.568 0.000 100.888 0.600 ;
 END
 ANTENNAPARTIALMETALAREA                  5.273 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME3 ;
 ANTENNADIFFAREA                          1.293 LAYER ME4 ;
END DO24
PIN DI23
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 97.126 0.000 97.446 0.600 ;
  LAYER ME3 ;
  RECT 97.126 0.000 97.446 0.600 ;
  LAYER ME2 ;
  RECT 97.126 0.000 97.446 0.600 ;
  LAYER ME1 ;
  RECT 97.126 0.000 97.446 0.600 ;
 END
 ANTENNAPARTIALMETALAREA                  1.058 LAYER ME2 ;
 ANTENNAGATEAREA                          0.072 LAYER ME2 ;
 ANTENNAGATEAREA                          0.072 LAYER ME3 ;
 ANTENNAGATEAREA                          0.072 LAYER ME4 ;
 ANTENNADIFFAREA                          0.160 LAYER ME2 ;
 ANTENNADIFFAREA                          0.160 LAYER ME3 ;
 ANTENNADIFFAREA                          0.160 LAYER ME4 ;
 ANTENNAMAXAREACAR                       21.782 LAYER ME2 ;
 ANTENNAMAXAREACAR                       24.449 LAYER ME3 ;
 ANTENNAMAXAREACAR                       27.116 LAYER ME4 ;
END DI23
PIN DO23
  DIRECTION OUTPUT ;
 PORT
  LAYER ME4 ;
  RECT 96.564 0.000 96.884 0.600 ;
  LAYER ME3 ;
  RECT 96.564 0.000 96.884 0.600 ;
  LAYER ME2 ;
  RECT 96.564 0.000 96.884 0.600 ;
  LAYER ME1 ;
  RECT 96.564 0.000 96.884 0.600 ;
 END
 ANTENNAPARTIALMETALAREA                  5.273 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME3 ;
 ANTENNADIFFAREA                          1.293 LAYER ME4 ;
END DO23
PIN DI22
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 92.560 0.000 92.880 0.600 ;
  LAYER ME3 ;
  RECT 92.560 0.000 92.880 0.600 ;
  LAYER ME2 ;
  RECT 92.560 0.000 92.880 0.600 ;
  LAYER ME1 ;
  RECT 92.560 0.000 92.880 0.600 ;
 END
 ANTENNAPARTIALMETALAREA                  0.346 LAYER ME1 ;
 ANTENNAPARTIALMETALAREA                  1.466 LAYER ME2 ;
 ANTENNAPARTIALMETALAREA                  0.508 LAYER ME3 ;
 ANTENNAGATEAREA                          0.072 LAYER ME3 ;
 ANTENNAGATEAREA                          0.072 LAYER ME4 ;
 ANTENNADIFFAREA                          0.218 LAYER ME1 ;
 ANTENNADIFFAREA                          0.218 LAYER ME2 ;
 ANTENNADIFFAREA                          0.218 LAYER ME3 ;
 ANTENNADIFFAREA                          0.218 LAYER ME4 ;
 ANTENNAMAXAREACAR                       17.267 LAYER ME3 ;
 ANTENNAMAXAREACAR                       19.933 LAYER ME4 ;
END DI22
PIN DO22
  DIRECTION OUTPUT ;
 PORT
  LAYER ME4 ;
  RECT 93.122 0.000 93.442 0.600 ;
  LAYER ME3 ;
  RECT 93.122 0.000 93.442 0.600 ;
  LAYER ME2 ;
  RECT 93.122 0.000 93.442 0.600 ;
  LAYER ME1 ;
  RECT 93.122 0.000 93.442 0.600 ;
 END
 ANTENNAPARTIALMETALAREA                  5.602 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME3 ;
 ANTENNADIFFAREA                          1.293 LAYER ME4 ;
END DO22
PIN WEB2
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 91.120 0.000 91.440 0.600 ;
  LAYER ME3 ;
  RECT 91.120 0.000 91.440 0.600 ;
  LAYER ME2 ;
  RECT 91.120 0.000 91.440 0.600 ;
  LAYER ME1 ;
  RECT 91.120 0.000 91.440 0.600 ;
 END
 ANTENNAPARTIALMETALAREA                  1.036 LAYER ME2 ;
 ANTENNAGATEAREA                          0.288 LAYER ME2 ;
 ANTENNAGATEAREA                          0.288 LAYER ME3 ;
 ANTENNAGATEAREA                          0.288 LAYER ME4 ;
 ANTENNADIFFAREA                          0.206 LAYER ME2 ;
 ANTENNADIFFAREA                          0.206 LAYER ME3 ;
 ANTENNADIFFAREA                          0.206 LAYER ME4 ;
 ANTENNAMAXAREACAR                        5.844 LAYER ME2 ;
 ANTENNAMAXAREACAR                        6.511 LAYER ME3 ;
 ANTENNAMAXAREACAR                        7.178 LAYER ME4 ;
END WEB2
PIN DI21
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 89.118 0.000 89.438 0.600 ;
  LAYER ME3 ;
  RECT 89.118 0.000 89.438 0.600 ;
  LAYER ME2 ;
  RECT 89.118 0.000 89.438 0.600 ;
  LAYER ME1 ;
  RECT 89.118 0.000 89.438 0.600 ;
 END
 ANTENNAPARTIALMETALAREA                  1.058 LAYER ME2 ;
 ANTENNAGATEAREA                          0.072 LAYER ME2 ;
 ANTENNAGATEAREA                          0.072 LAYER ME3 ;
 ANTENNAGATEAREA                          0.072 LAYER ME4 ;
 ANTENNADIFFAREA                          0.160 LAYER ME2 ;
 ANTENNADIFFAREA                          0.160 LAYER ME3 ;
 ANTENNADIFFAREA                          0.160 LAYER ME4 ;
 ANTENNAMAXAREACAR                       21.782 LAYER ME2 ;
 ANTENNAMAXAREACAR                       24.449 LAYER ME3 ;
 ANTENNAMAXAREACAR                       27.116 LAYER ME4 ;
END DI21
PIN DO21
  DIRECTION OUTPUT ;
 PORT
  LAYER ME4 ;
  RECT 88.556 0.000 88.876 0.600 ;
  LAYER ME3 ;
  RECT 88.556 0.000 88.876 0.600 ;
  LAYER ME2 ;
  RECT 88.556 0.000 88.876 0.600 ;
  LAYER ME1 ;
  RECT 88.556 0.000 88.876 0.600 ;
 END
 ANTENNAPARTIALMETALAREA                  5.273 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME3 ;
 ANTENNADIFFAREA                          1.293 LAYER ME4 ;
END DO21
PIN DI20
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 85.114 0.000 85.434 0.600 ;
  LAYER ME3 ;
  RECT 85.114 0.000 85.434 0.600 ;
  LAYER ME2 ;
  RECT 85.114 0.000 85.434 0.600 ;
  LAYER ME1 ;
  RECT 85.114 0.000 85.434 0.600 ;
 END
 ANTENNAPARTIALMETALAREA                  1.058 LAYER ME2 ;
 ANTENNAGATEAREA                          0.072 LAYER ME2 ;
 ANTENNAGATEAREA                          0.072 LAYER ME3 ;
 ANTENNAGATEAREA                          0.072 LAYER ME4 ;
 ANTENNADIFFAREA                          0.160 LAYER ME2 ;
 ANTENNADIFFAREA                          0.160 LAYER ME3 ;
 ANTENNADIFFAREA                          0.160 LAYER ME4 ;
 ANTENNAMAXAREACAR                       21.782 LAYER ME2 ;
 ANTENNAMAXAREACAR                       24.449 LAYER ME3 ;
 ANTENNAMAXAREACAR                       27.116 LAYER ME4 ;
END DI20
PIN DO20
  DIRECTION OUTPUT ;
 PORT
  LAYER ME4 ;
  RECT 84.552 0.000 84.872 0.600 ;
  LAYER ME3 ;
  RECT 84.552 0.000 84.872 0.600 ;
  LAYER ME2 ;
  RECT 84.552 0.000 84.872 0.600 ;
  LAYER ME1 ;
  RECT 84.552 0.000 84.872 0.600 ;
 END
 ANTENNAPARTIALMETALAREA                  5.273 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME3 ;
 ANTENNADIFFAREA                          1.293 LAYER ME4 ;
END DO20
PIN DI19
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 81.110 0.000 81.430 0.600 ;
  LAYER ME3 ;
  RECT 81.110 0.000 81.430 0.600 ;
  LAYER ME2 ;
  RECT 81.110 0.000 81.430 0.600 ;
  LAYER ME1 ;
  RECT 81.110 0.000 81.430 0.600 ;
 END
 ANTENNAPARTIALMETALAREA                  1.058 LAYER ME2 ;
 ANTENNAGATEAREA                          0.072 LAYER ME2 ;
 ANTENNAGATEAREA                          0.072 LAYER ME3 ;
 ANTENNAGATEAREA                          0.072 LAYER ME4 ;
 ANTENNADIFFAREA                          0.160 LAYER ME2 ;
 ANTENNADIFFAREA                          0.160 LAYER ME3 ;
 ANTENNADIFFAREA                          0.160 LAYER ME4 ;
 ANTENNAMAXAREACAR                       21.782 LAYER ME2 ;
 ANTENNAMAXAREACAR                       24.449 LAYER ME3 ;
 ANTENNAMAXAREACAR                       27.116 LAYER ME4 ;
END DI19
PIN DO19
  DIRECTION OUTPUT ;
 PORT
  LAYER ME4 ;
  RECT 80.548 0.000 80.868 0.600 ;
  LAYER ME3 ;
  RECT 80.548 0.000 80.868 0.600 ;
  LAYER ME2 ;
  RECT 80.548 0.000 80.868 0.600 ;
  LAYER ME1 ;
  RECT 80.548 0.000 80.868 0.600 ;
 END
 ANTENNAPARTIALMETALAREA                  5.273 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME3 ;
 ANTENNADIFFAREA                          1.293 LAYER ME4 ;
END DO19
PIN DI18
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 77.106 0.000 77.426 0.600 ;
  LAYER ME3 ;
  RECT 77.106 0.000 77.426 0.600 ;
  LAYER ME2 ;
  RECT 77.106 0.000 77.426 0.600 ;
  LAYER ME1 ;
  RECT 77.106 0.000 77.426 0.600 ;
 END
 ANTENNAPARTIALMETALAREA                  1.058 LAYER ME2 ;
 ANTENNAGATEAREA                          0.072 LAYER ME2 ;
 ANTENNAGATEAREA                          0.072 LAYER ME3 ;
 ANTENNAGATEAREA                          0.072 LAYER ME4 ;
 ANTENNADIFFAREA                          0.160 LAYER ME2 ;
 ANTENNADIFFAREA                          0.160 LAYER ME3 ;
 ANTENNADIFFAREA                          0.160 LAYER ME4 ;
 ANTENNAMAXAREACAR                       21.782 LAYER ME2 ;
 ANTENNAMAXAREACAR                       24.449 LAYER ME3 ;
 ANTENNAMAXAREACAR                       27.116 LAYER ME4 ;
END DI18
PIN DO18
  DIRECTION OUTPUT ;
 PORT
  LAYER ME4 ;
  RECT 76.544 0.000 76.864 0.600 ;
  LAYER ME3 ;
  RECT 76.544 0.000 76.864 0.600 ;
  LAYER ME2 ;
  RECT 76.544 0.000 76.864 0.600 ;
  LAYER ME1 ;
  RECT 76.544 0.000 76.864 0.600 ;
 END
 ANTENNAPARTIALMETALAREA                  5.273 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME3 ;
 ANTENNADIFFAREA                          1.293 LAYER ME4 ;
END DO18
PIN DI17
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 73.102 0.000 73.422 0.600 ;
  LAYER ME3 ;
  RECT 73.102 0.000 73.422 0.600 ;
  LAYER ME2 ;
  RECT 73.102 0.000 73.422 0.600 ;
  LAYER ME1 ;
  RECT 73.102 0.000 73.422 0.600 ;
 END
 ANTENNAPARTIALMETALAREA                  1.058 LAYER ME2 ;
 ANTENNAGATEAREA                          0.072 LAYER ME2 ;
 ANTENNAGATEAREA                          0.072 LAYER ME3 ;
 ANTENNAGATEAREA                          0.072 LAYER ME4 ;
 ANTENNADIFFAREA                          0.160 LAYER ME2 ;
 ANTENNADIFFAREA                          0.160 LAYER ME3 ;
 ANTENNADIFFAREA                          0.160 LAYER ME4 ;
 ANTENNAMAXAREACAR                       21.782 LAYER ME2 ;
 ANTENNAMAXAREACAR                       24.449 LAYER ME3 ;
 ANTENNAMAXAREACAR                       27.116 LAYER ME4 ;
END DI17
PIN DO17
  DIRECTION OUTPUT ;
 PORT
  LAYER ME4 ;
  RECT 72.540 0.000 72.860 0.600 ;
  LAYER ME3 ;
  RECT 72.540 0.000 72.860 0.600 ;
  LAYER ME2 ;
  RECT 72.540 0.000 72.860 0.600 ;
  LAYER ME1 ;
  RECT 72.540 0.000 72.860 0.600 ;
 END
 ANTENNAPARTIALMETALAREA                  5.273 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME3 ;
 ANTENNADIFFAREA                          1.293 LAYER ME4 ;
END DO17
PIN DI16
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 69.098 0.000 69.418 0.600 ;
  LAYER ME3 ;
  RECT 69.098 0.000 69.418 0.600 ;
  LAYER ME2 ;
  RECT 69.098 0.000 69.418 0.600 ;
  LAYER ME1 ;
  RECT 69.098 0.000 69.418 0.600 ;
 END
 ANTENNAPARTIALMETALAREA                  1.058 LAYER ME2 ;
 ANTENNAGATEAREA                          0.072 LAYER ME2 ;
 ANTENNAGATEAREA                          0.072 LAYER ME3 ;
 ANTENNAGATEAREA                          0.072 LAYER ME4 ;
 ANTENNADIFFAREA                          0.160 LAYER ME2 ;
 ANTENNADIFFAREA                          0.160 LAYER ME3 ;
 ANTENNADIFFAREA                          0.160 LAYER ME4 ;
 ANTENNAMAXAREACAR                       21.782 LAYER ME2 ;
 ANTENNAMAXAREACAR                       24.449 LAYER ME3 ;
 ANTENNAMAXAREACAR                       27.116 LAYER ME4 ;
END DI16
PIN DO16
  DIRECTION OUTPUT ;
 PORT
  LAYER ME4 ;
  RECT 68.536 0.000 68.856 0.600 ;
  LAYER ME3 ;
  RECT 68.536 0.000 68.856 0.600 ;
  LAYER ME2 ;
  RECT 68.536 0.000 68.856 0.600 ;
  LAYER ME1 ;
  RECT 68.536 0.000 68.856 0.600 ;
 END
 ANTENNAPARTIALMETALAREA                  5.273 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME3 ;
 ANTENNADIFFAREA                          1.293 LAYER ME4 ;
END DO16
PIN DI15
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 65.094 0.000 65.414 0.600 ;
  LAYER ME3 ;
  RECT 65.094 0.000 65.414 0.600 ;
  LAYER ME2 ;
  RECT 65.094 0.000 65.414 0.600 ;
  LAYER ME1 ;
  RECT 65.094 0.000 65.414 0.600 ;
 END
 ANTENNAPARTIALMETALAREA                  1.058 LAYER ME2 ;
 ANTENNAGATEAREA                          0.072 LAYER ME2 ;
 ANTENNAGATEAREA                          0.072 LAYER ME3 ;
 ANTENNAGATEAREA                          0.072 LAYER ME4 ;
 ANTENNADIFFAREA                          0.160 LAYER ME2 ;
 ANTENNADIFFAREA                          0.160 LAYER ME3 ;
 ANTENNADIFFAREA                          0.160 LAYER ME4 ;
 ANTENNAMAXAREACAR                       21.782 LAYER ME2 ;
 ANTENNAMAXAREACAR                       24.449 LAYER ME3 ;
 ANTENNAMAXAREACAR                       27.116 LAYER ME4 ;
END DI15
PIN DO15
  DIRECTION OUTPUT ;
 PORT
  LAYER ME4 ;
  RECT 64.532 0.000 64.852 0.600 ;
  LAYER ME3 ;
  RECT 64.532 0.000 64.852 0.600 ;
  LAYER ME2 ;
  RECT 64.532 0.000 64.852 0.600 ;
  LAYER ME1 ;
  RECT 64.532 0.000 64.852 0.600 ;
 END
 ANTENNAPARTIALMETALAREA                  5.273 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME3 ;
 ANTENNADIFFAREA                          1.293 LAYER ME4 ;
END DO15
PIN DI14
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 61.090 0.000 61.410 0.600 ;
  LAYER ME3 ;
  RECT 61.090 0.000 61.410 0.600 ;
  LAYER ME2 ;
  RECT 61.090 0.000 61.410 0.600 ;
  LAYER ME1 ;
  RECT 61.090 0.000 61.410 0.600 ;
 END
 ANTENNAPARTIALMETALAREA                  1.058 LAYER ME2 ;
 ANTENNAGATEAREA                          0.072 LAYER ME2 ;
 ANTENNAGATEAREA                          0.072 LAYER ME3 ;
 ANTENNAGATEAREA                          0.072 LAYER ME4 ;
 ANTENNADIFFAREA                          0.160 LAYER ME2 ;
 ANTENNADIFFAREA                          0.160 LAYER ME3 ;
 ANTENNADIFFAREA                          0.160 LAYER ME4 ;
 ANTENNAMAXAREACAR                       21.782 LAYER ME2 ;
 ANTENNAMAXAREACAR                       24.449 LAYER ME3 ;
 ANTENNAMAXAREACAR                       27.116 LAYER ME4 ;
END DI14
PIN DO14
  DIRECTION OUTPUT ;
 PORT
  LAYER ME4 ;
  RECT 60.528 0.000 60.848 0.600 ;
  LAYER ME3 ;
  RECT 60.528 0.000 60.848 0.600 ;
  LAYER ME2 ;
  RECT 60.528 0.000 60.848 0.600 ;
  LAYER ME1 ;
  RECT 60.528 0.000 60.848 0.600 ;
 END
 ANTENNAPARTIALMETALAREA                  5.273 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME3 ;
 ANTENNADIFFAREA                          1.293 LAYER ME4 ;
END DO14
PIN DI13
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 57.086 0.000 57.406 0.600 ;
  LAYER ME3 ;
  RECT 57.086 0.000 57.406 0.600 ;
  LAYER ME2 ;
  RECT 57.086 0.000 57.406 0.600 ;
  LAYER ME1 ;
  RECT 57.086 0.000 57.406 0.600 ;
 END
 ANTENNAPARTIALMETALAREA                  1.058 LAYER ME2 ;
 ANTENNAGATEAREA                          0.072 LAYER ME2 ;
 ANTENNAGATEAREA                          0.072 LAYER ME3 ;
 ANTENNAGATEAREA                          0.072 LAYER ME4 ;
 ANTENNADIFFAREA                          0.160 LAYER ME2 ;
 ANTENNADIFFAREA                          0.160 LAYER ME3 ;
 ANTENNADIFFAREA                          0.160 LAYER ME4 ;
 ANTENNAMAXAREACAR                       21.782 LAYER ME2 ;
 ANTENNAMAXAREACAR                       24.449 LAYER ME3 ;
 ANTENNAMAXAREACAR                       27.116 LAYER ME4 ;
END DI13
PIN DO13
  DIRECTION OUTPUT ;
 PORT
  LAYER ME4 ;
  RECT 56.524 0.000 56.844 0.600 ;
  LAYER ME3 ;
  RECT 56.524 0.000 56.844 0.600 ;
  LAYER ME2 ;
  RECT 56.524 0.000 56.844 0.600 ;
  LAYER ME1 ;
  RECT 56.524 0.000 56.844 0.600 ;
 END
 ANTENNAPARTIALMETALAREA                  5.273 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME3 ;
 ANTENNADIFFAREA                          1.293 LAYER ME4 ;
END DO13
PIN DI12
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 53.082 0.000 53.402 0.600 ;
  LAYER ME3 ;
  RECT 53.082 0.000 53.402 0.600 ;
  LAYER ME2 ;
  RECT 53.082 0.000 53.402 0.600 ;
  LAYER ME1 ;
  RECT 53.082 0.000 53.402 0.600 ;
 END
 ANTENNAPARTIALMETALAREA                  1.058 LAYER ME2 ;
 ANTENNAGATEAREA                          0.072 LAYER ME2 ;
 ANTENNAGATEAREA                          0.072 LAYER ME3 ;
 ANTENNAGATEAREA                          0.072 LAYER ME4 ;
 ANTENNADIFFAREA                          0.160 LAYER ME2 ;
 ANTENNADIFFAREA                          0.160 LAYER ME3 ;
 ANTENNADIFFAREA                          0.160 LAYER ME4 ;
 ANTENNAMAXAREACAR                       21.782 LAYER ME2 ;
 ANTENNAMAXAREACAR                       24.449 LAYER ME3 ;
 ANTENNAMAXAREACAR                       27.116 LAYER ME4 ;
END DI12
PIN DO12
  DIRECTION OUTPUT ;
 PORT
  LAYER ME4 ;
  RECT 52.520 0.000 52.840 0.600 ;
  LAYER ME3 ;
  RECT 52.520 0.000 52.840 0.600 ;
  LAYER ME2 ;
  RECT 52.520 0.000 52.840 0.600 ;
  LAYER ME1 ;
  RECT 52.520 0.000 52.840 0.600 ;
 END
 ANTENNAPARTIALMETALAREA                  5.273 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME3 ;
 ANTENNADIFFAREA                          1.293 LAYER ME4 ;
END DO12
PIN DI11
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 48.516 0.000 48.836 0.600 ;
  LAYER ME3 ;
  RECT 48.516 0.000 48.836 0.600 ;
  LAYER ME2 ;
  RECT 48.516 0.000 48.836 0.600 ;
  LAYER ME1 ;
  RECT 48.516 0.000 48.836 0.600 ;
 END
 ANTENNAPARTIALMETALAREA                  0.346 LAYER ME1 ;
 ANTENNAPARTIALMETALAREA                  1.466 LAYER ME2 ;
 ANTENNAPARTIALMETALAREA                  0.508 LAYER ME3 ;
 ANTENNAGATEAREA                          0.072 LAYER ME3 ;
 ANTENNAGATEAREA                          0.072 LAYER ME4 ;
 ANTENNADIFFAREA                          0.218 LAYER ME1 ;
 ANTENNADIFFAREA                          0.218 LAYER ME2 ;
 ANTENNADIFFAREA                          0.218 LAYER ME3 ;
 ANTENNADIFFAREA                          0.218 LAYER ME4 ;
 ANTENNAMAXAREACAR                       17.267 LAYER ME3 ;
 ANTENNAMAXAREACAR                       19.933 LAYER ME4 ;
END DI11
PIN DO11
  DIRECTION OUTPUT ;
 PORT
  LAYER ME4 ;
  RECT 49.078 0.000 49.398 0.600 ;
  LAYER ME3 ;
  RECT 49.078 0.000 49.398 0.600 ;
  LAYER ME2 ;
  RECT 49.078 0.000 49.398 0.600 ;
  LAYER ME1 ;
  RECT 49.078 0.000 49.398 0.600 ;
 END
 ANTENNAPARTIALMETALAREA                  5.602 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME3 ;
 ANTENNADIFFAREA                          1.293 LAYER ME4 ;
END DO11
PIN WEB1
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 47.076 0.000 47.396 0.600 ;
  LAYER ME3 ;
  RECT 47.076 0.000 47.396 0.600 ;
  LAYER ME2 ;
  RECT 47.076 0.000 47.396 0.600 ;
  LAYER ME1 ;
  RECT 47.076 0.000 47.396 0.600 ;
 END
 ANTENNAPARTIALMETALAREA                  1.036 LAYER ME2 ;
 ANTENNAGATEAREA                          0.288 LAYER ME2 ;
 ANTENNAGATEAREA                          0.288 LAYER ME3 ;
 ANTENNAGATEAREA                          0.288 LAYER ME4 ;
 ANTENNADIFFAREA                          0.206 LAYER ME2 ;
 ANTENNADIFFAREA                          0.206 LAYER ME3 ;
 ANTENNADIFFAREA                          0.206 LAYER ME4 ;
 ANTENNAMAXAREACAR                        5.844 LAYER ME2 ;
 ANTENNAMAXAREACAR                        6.511 LAYER ME3 ;
 ANTENNAMAXAREACAR                        7.178 LAYER ME4 ;
END WEB1
PIN DI10
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 45.074 0.000 45.394 0.600 ;
  LAYER ME3 ;
  RECT 45.074 0.000 45.394 0.600 ;
  LAYER ME2 ;
  RECT 45.074 0.000 45.394 0.600 ;
  LAYER ME1 ;
  RECT 45.074 0.000 45.394 0.600 ;
 END
 ANTENNAPARTIALMETALAREA                  1.058 LAYER ME2 ;
 ANTENNAGATEAREA                          0.072 LAYER ME2 ;
 ANTENNAGATEAREA                          0.072 LAYER ME3 ;
 ANTENNAGATEAREA                          0.072 LAYER ME4 ;
 ANTENNADIFFAREA                          0.160 LAYER ME2 ;
 ANTENNADIFFAREA                          0.160 LAYER ME3 ;
 ANTENNADIFFAREA                          0.160 LAYER ME4 ;
 ANTENNAMAXAREACAR                       21.782 LAYER ME2 ;
 ANTENNAMAXAREACAR                       24.449 LAYER ME3 ;
 ANTENNAMAXAREACAR                       27.116 LAYER ME4 ;
END DI10
PIN DO10
  DIRECTION OUTPUT ;
 PORT
  LAYER ME4 ;
  RECT 44.512 0.000 44.832 0.600 ;
  LAYER ME3 ;
  RECT 44.512 0.000 44.832 0.600 ;
  LAYER ME2 ;
  RECT 44.512 0.000 44.832 0.600 ;
  LAYER ME1 ;
  RECT 44.512 0.000 44.832 0.600 ;
 END
 ANTENNAPARTIALMETALAREA                  5.273 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME3 ;
 ANTENNADIFFAREA                          1.293 LAYER ME4 ;
END DO10
PIN DI9
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 41.070 0.000 41.390 0.600 ;
  LAYER ME3 ;
  RECT 41.070 0.000 41.390 0.600 ;
  LAYER ME2 ;
  RECT 41.070 0.000 41.390 0.600 ;
  LAYER ME1 ;
  RECT 41.070 0.000 41.390 0.600 ;
 END
 ANTENNAPARTIALMETALAREA                  1.058 LAYER ME2 ;
 ANTENNAGATEAREA                          0.072 LAYER ME2 ;
 ANTENNAGATEAREA                          0.072 LAYER ME3 ;
 ANTENNAGATEAREA                          0.072 LAYER ME4 ;
 ANTENNADIFFAREA                          0.160 LAYER ME2 ;
 ANTENNADIFFAREA                          0.160 LAYER ME3 ;
 ANTENNADIFFAREA                          0.160 LAYER ME4 ;
 ANTENNAMAXAREACAR                       21.782 LAYER ME2 ;
 ANTENNAMAXAREACAR                       24.449 LAYER ME3 ;
 ANTENNAMAXAREACAR                       27.116 LAYER ME4 ;
END DI9
PIN DO9
  DIRECTION OUTPUT ;
 PORT
  LAYER ME4 ;
  RECT 40.508 0.000 40.828 0.600 ;
  LAYER ME3 ;
  RECT 40.508 0.000 40.828 0.600 ;
  LAYER ME2 ;
  RECT 40.508 0.000 40.828 0.600 ;
  LAYER ME1 ;
  RECT 40.508 0.000 40.828 0.600 ;
 END
 ANTENNAPARTIALMETALAREA                  5.273 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME3 ;
 ANTENNADIFFAREA                          1.293 LAYER ME4 ;
END DO9
PIN DI8
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 37.066 0.000 37.386 0.600 ;
  LAYER ME3 ;
  RECT 37.066 0.000 37.386 0.600 ;
  LAYER ME2 ;
  RECT 37.066 0.000 37.386 0.600 ;
  LAYER ME1 ;
  RECT 37.066 0.000 37.386 0.600 ;
 END
 ANTENNAPARTIALMETALAREA                  1.058 LAYER ME2 ;
 ANTENNAGATEAREA                          0.072 LAYER ME2 ;
 ANTENNAGATEAREA                          0.072 LAYER ME3 ;
 ANTENNAGATEAREA                          0.072 LAYER ME4 ;
 ANTENNADIFFAREA                          0.160 LAYER ME2 ;
 ANTENNADIFFAREA                          0.160 LAYER ME3 ;
 ANTENNADIFFAREA                          0.160 LAYER ME4 ;
 ANTENNAMAXAREACAR                       21.782 LAYER ME2 ;
 ANTENNAMAXAREACAR                       24.449 LAYER ME3 ;
 ANTENNAMAXAREACAR                       27.116 LAYER ME4 ;
END DI8
PIN DO8
  DIRECTION OUTPUT ;
 PORT
  LAYER ME4 ;
  RECT 36.504 0.000 36.824 0.600 ;
  LAYER ME3 ;
  RECT 36.504 0.000 36.824 0.600 ;
  LAYER ME2 ;
  RECT 36.504 0.000 36.824 0.600 ;
  LAYER ME1 ;
  RECT 36.504 0.000 36.824 0.600 ;
 END
 ANTENNAPARTIALMETALAREA                  5.273 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME3 ;
 ANTENNADIFFAREA                          1.293 LAYER ME4 ;
END DO8
PIN DI7
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 33.062 0.000 33.382 0.600 ;
  LAYER ME3 ;
  RECT 33.062 0.000 33.382 0.600 ;
  LAYER ME2 ;
  RECT 33.062 0.000 33.382 0.600 ;
  LAYER ME1 ;
  RECT 33.062 0.000 33.382 0.600 ;
 END
 ANTENNAPARTIALMETALAREA                  1.058 LAYER ME2 ;
 ANTENNAGATEAREA                          0.072 LAYER ME2 ;
 ANTENNAGATEAREA                          0.072 LAYER ME3 ;
 ANTENNAGATEAREA                          0.072 LAYER ME4 ;
 ANTENNADIFFAREA                          0.160 LAYER ME2 ;
 ANTENNADIFFAREA                          0.160 LAYER ME3 ;
 ANTENNADIFFAREA                          0.160 LAYER ME4 ;
 ANTENNAMAXAREACAR                       21.782 LAYER ME2 ;
 ANTENNAMAXAREACAR                       24.449 LAYER ME3 ;
 ANTENNAMAXAREACAR                       27.116 LAYER ME4 ;
END DI7
PIN DO7
  DIRECTION OUTPUT ;
 PORT
  LAYER ME4 ;
  RECT 32.500 0.000 32.820 0.600 ;
  LAYER ME3 ;
  RECT 32.500 0.000 32.820 0.600 ;
  LAYER ME2 ;
  RECT 32.500 0.000 32.820 0.600 ;
  LAYER ME1 ;
  RECT 32.500 0.000 32.820 0.600 ;
 END
 ANTENNAPARTIALMETALAREA                  5.273 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME3 ;
 ANTENNADIFFAREA                          1.293 LAYER ME4 ;
END DO7
PIN DI6
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 29.058 0.000 29.378 0.600 ;
  LAYER ME3 ;
  RECT 29.058 0.000 29.378 0.600 ;
  LAYER ME2 ;
  RECT 29.058 0.000 29.378 0.600 ;
  LAYER ME1 ;
  RECT 29.058 0.000 29.378 0.600 ;
 END
 ANTENNAPARTIALMETALAREA                  1.058 LAYER ME2 ;
 ANTENNAGATEAREA                          0.072 LAYER ME2 ;
 ANTENNAGATEAREA                          0.072 LAYER ME3 ;
 ANTENNAGATEAREA                          0.072 LAYER ME4 ;
 ANTENNADIFFAREA                          0.160 LAYER ME2 ;
 ANTENNADIFFAREA                          0.160 LAYER ME3 ;
 ANTENNADIFFAREA                          0.160 LAYER ME4 ;
 ANTENNAMAXAREACAR                       21.782 LAYER ME2 ;
 ANTENNAMAXAREACAR                       24.449 LAYER ME3 ;
 ANTENNAMAXAREACAR                       27.116 LAYER ME4 ;
END DI6
PIN DO6
  DIRECTION OUTPUT ;
 PORT
  LAYER ME4 ;
  RECT 28.496 0.000 28.816 0.600 ;
  LAYER ME3 ;
  RECT 28.496 0.000 28.816 0.600 ;
  LAYER ME2 ;
  RECT 28.496 0.000 28.816 0.600 ;
  LAYER ME1 ;
  RECT 28.496 0.000 28.816 0.600 ;
 END
 ANTENNAPARTIALMETALAREA                  5.273 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME3 ;
 ANTENNADIFFAREA                          1.293 LAYER ME4 ;
END DO6
PIN DI5
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 25.054 0.000 25.374 0.600 ;
  LAYER ME3 ;
  RECT 25.054 0.000 25.374 0.600 ;
  LAYER ME2 ;
  RECT 25.054 0.000 25.374 0.600 ;
  LAYER ME1 ;
  RECT 25.054 0.000 25.374 0.600 ;
 END
 ANTENNAPARTIALMETALAREA                  1.058 LAYER ME2 ;
 ANTENNAGATEAREA                          0.072 LAYER ME2 ;
 ANTENNAGATEAREA                          0.072 LAYER ME3 ;
 ANTENNAGATEAREA                          0.072 LAYER ME4 ;
 ANTENNADIFFAREA                          0.160 LAYER ME2 ;
 ANTENNADIFFAREA                          0.160 LAYER ME3 ;
 ANTENNADIFFAREA                          0.160 LAYER ME4 ;
 ANTENNAMAXAREACAR                       21.782 LAYER ME2 ;
 ANTENNAMAXAREACAR                       24.449 LAYER ME3 ;
 ANTENNAMAXAREACAR                       27.116 LAYER ME4 ;
END DI5
PIN DO5
  DIRECTION OUTPUT ;
 PORT
  LAYER ME4 ;
  RECT 24.492 0.000 24.812 0.600 ;
  LAYER ME3 ;
  RECT 24.492 0.000 24.812 0.600 ;
  LAYER ME2 ;
  RECT 24.492 0.000 24.812 0.600 ;
  LAYER ME1 ;
  RECT 24.492 0.000 24.812 0.600 ;
 END
 ANTENNAPARTIALMETALAREA                  5.273 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME3 ;
 ANTENNADIFFAREA                          1.293 LAYER ME4 ;
END DO5
PIN DI4
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 21.050 0.000 21.370 0.600 ;
  LAYER ME3 ;
  RECT 21.050 0.000 21.370 0.600 ;
  LAYER ME2 ;
  RECT 21.050 0.000 21.370 0.600 ;
  LAYER ME1 ;
  RECT 21.050 0.000 21.370 0.600 ;
 END
 ANTENNAPARTIALMETALAREA                  1.058 LAYER ME2 ;
 ANTENNAGATEAREA                          0.072 LAYER ME2 ;
 ANTENNAGATEAREA                          0.072 LAYER ME3 ;
 ANTENNAGATEAREA                          0.072 LAYER ME4 ;
 ANTENNADIFFAREA                          0.160 LAYER ME2 ;
 ANTENNADIFFAREA                          0.160 LAYER ME3 ;
 ANTENNADIFFAREA                          0.160 LAYER ME4 ;
 ANTENNAMAXAREACAR                       21.782 LAYER ME2 ;
 ANTENNAMAXAREACAR                       24.449 LAYER ME3 ;
 ANTENNAMAXAREACAR                       27.116 LAYER ME4 ;
END DI4
PIN DO4
  DIRECTION OUTPUT ;
 PORT
  LAYER ME4 ;
  RECT 20.488 0.000 20.808 0.600 ;
  LAYER ME3 ;
  RECT 20.488 0.000 20.808 0.600 ;
  LAYER ME2 ;
  RECT 20.488 0.000 20.808 0.600 ;
  LAYER ME1 ;
  RECT 20.488 0.000 20.808 0.600 ;
 END
 ANTENNAPARTIALMETALAREA                  5.273 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME3 ;
 ANTENNADIFFAREA                          1.293 LAYER ME4 ;
END DO4
PIN DI3
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 17.046 0.000 17.366 0.600 ;
  LAYER ME3 ;
  RECT 17.046 0.000 17.366 0.600 ;
  LAYER ME2 ;
  RECT 17.046 0.000 17.366 0.600 ;
  LAYER ME1 ;
  RECT 17.046 0.000 17.366 0.600 ;
 END
 ANTENNAPARTIALMETALAREA                  1.058 LAYER ME2 ;
 ANTENNAGATEAREA                          0.072 LAYER ME2 ;
 ANTENNAGATEAREA                          0.072 LAYER ME3 ;
 ANTENNAGATEAREA                          0.072 LAYER ME4 ;
 ANTENNADIFFAREA                          0.160 LAYER ME2 ;
 ANTENNADIFFAREA                          0.160 LAYER ME3 ;
 ANTENNADIFFAREA                          0.160 LAYER ME4 ;
 ANTENNAMAXAREACAR                       21.782 LAYER ME2 ;
 ANTENNAMAXAREACAR                       24.449 LAYER ME3 ;
 ANTENNAMAXAREACAR                       27.116 LAYER ME4 ;
END DI3
PIN DO3
  DIRECTION OUTPUT ;
 PORT
  LAYER ME4 ;
  RECT 16.484 0.000 16.804 0.600 ;
  LAYER ME3 ;
  RECT 16.484 0.000 16.804 0.600 ;
  LAYER ME2 ;
  RECT 16.484 0.000 16.804 0.600 ;
  LAYER ME1 ;
  RECT 16.484 0.000 16.804 0.600 ;
 END
 ANTENNAPARTIALMETALAREA                  5.273 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME3 ;
 ANTENNADIFFAREA                          1.293 LAYER ME4 ;
END DO3
PIN DI2
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 13.042 0.000 13.362 0.600 ;
  LAYER ME3 ;
  RECT 13.042 0.000 13.362 0.600 ;
  LAYER ME2 ;
  RECT 13.042 0.000 13.362 0.600 ;
  LAYER ME1 ;
  RECT 13.042 0.000 13.362 0.600 ;
 END
 ANTENNAPARTIALMETALAREA                  1.058 LAYER ME2 ;
 ANTENNAGATEAREA                          0.072 LAYER ME2 ;
 ANTENNAGATEAREA                          0.072 LAYER ME3 ;
 ANTENNAGATEAREA                          0.072 LAYER ME4 ;
 ANTENNADIFFAREA                          0.160 LAYER ME2 ;
 ANTENNADIFFAREA                          0.160 LAYER ME3 ;
 ANTENNADIFFAREA                          0.160 LAYER ME4 ;
 ANTENNAMAXAREACAR                       21.782 LAYER ME2 ;
 ANTENNAMAXAREACAR                       24.449 LAYER ME3 ;
 ANTENNAMAXAREACAR                       27.116 LAYER ME4 ;
END DI2
PIN DO2
  DIRECTION OUTPUT ;
 PORT
  LAYER ME4 ;
  RECT 12.480 0.000 12.800 0.600 ;
  LAYER ME3 ;
  RECT 12.480 0.000 12.800 0.600 ;
  LAYER ME2 ;
  RECT 12.480 0.000 12.800 0.600 ;
  LAYER ME1 ;
  RECT 12.480 0.000 12.800 0.600 ;
 END
 ANTENNAPARTIALMETALAREA                  5.273 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME3 ;
 ANTENNADIFFAREA                          1.293 LAYER ME4 ;
END DO2
PIN DI1
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 9.038 0.000 9.358 0.600 ;
  LAYER ME3 ;
  RECT 9.038 0.000 9.358 0.600 ;
  LAYER ME2 ;
  RECT 9.038 0.000 9.358 0.600 ;
  LAYER ME1 ;
  RECT 9.038 0.000 9.358 0.600 ;
 END
 ANTENNAPARTIALMETALAREA                  1.058 LAYER ME2 ;
 ANTENNAGATEAREA                          0.072 LAYER ME2 ;
 ANTENNAGATEAREA                          0.072 LAYER ME3 ;
 ANTENNAGATEAREA                          0.072 LAYER ME4 ;
 ANTENNADIFFAREA                          0.160 LAYER ME2 ;
 ANTENNADIFFAREA                          0.160 LAYER ME3 ;
 ANTENNADIFFAREA                          0.160 LAYER ME4 ;
 ANTENNAMAXAREACAR                       21.782 LAYER ME2 ;
 ANTENNAMAXAREACAR                       24.449 LAYER ME3 ;
 ANTENNAMAXAREACAR                       27.116 LAYER ME4 ;
END DI1
PIN DO1
  DIRECTION OUTPUT ;
 PORT
  LAYER ME4 ;
  RECT 8.476 0.000 8.796 0.600 ;
  LAYER ME3 ;
  RECT 8.476 0.000 8.796 0.600 ;
  LAYER ME2 ;
  RECT 8.476 0.000 8.796 0.600 ;
  LAYER ME1 ;
  RECT 8.476 0.000 8.796 0.600 ;
 END
 ANTENNAPARTIALMETALAREA                  5.273 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME3 ;
 ANTENNADIFFAREA                          1.293 LAYER ME4 ;
END DO1
PIN DI0
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 4.472 0.000 4.792 0.600 ;
  LAYER ME3 ;
  RECT 4.472 0.000 4.792 0.600 ;
  LAYER ME2 ;
  RECT 4.472 0.000 4.792 0.600 ;
  LAYER ME1 ;
  RECT 4.472 0.000 4.792 0.600 ;
 END
 ANTENNAPARTIALMETALAREA                  0.346 LAYER ME1 ;
 ANTENNAPARTIALMETALAREA                  1.466 LAYER ME2 ;
 ANTENNAPARTIALMETALAREA                  0.508 LAYER ME3 ;
 ANTENNAGATEAREA                          0.072 LAYER ME3 ;
 ANTENNAGATEAREA                          0.072 LAYER ME4 ;
 ANTENNADIFFAREA                          0.218 LAYER ME1 ;
 ANTENNADIFFAREA                          0.218 LAYER ME2 ;
 ANTENNADIFFAREA                          0.218 LAYER ME3 ;
 ANTENNADIFFAREA                          0.218 LAYER ME4 ;
 ANTENNAMAXAREACAR                       17.267 LAYER ME3 ;
 ANTENNAMAXAREACAR                       19.933 LAYER ME4 ;
END DI0
PIN DO0
  DIRECTION OUTPUT ;
 PORT
  LAYER ME4 ;
  RECT 5.034 0.000 5.354 0.600 ;
  LAYER ME3 ;
  RECT 5.034 0.000 5.354 0.600 ;
  LAYER ME2 ;
  RECT 5.034 0.000 5.354 0.600 ;
  LAYER ME1 ;
  RECT 5.034 0.000 5.354 0.600 ;
 END
 ANTENNAPARTIALMETALAREA                  5.602 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME3 ;
 ANTENNADIFFAREA                          1.293 LAYER ME4 ;
END DO0
PIN WEB0
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 3.032 0.000 3.352 0.600 ;
  LAYER ME3 ;
  RECT 3.032 0.000 3.352 0.600 ;
  LAYER ME2 ;
  RECT 3.032 0.000 3.352 0.600 ;
  LAYER ME1 ;
  RECT 3.032 0.000 3.352 0.600 ;
 END
 ANTENNAPARTIALMETALAREA                  1.036 LAYER ME2 ;
 ANTENNAGATEAREA                          0.288 LAYER ME2 ;
 ANTENNAGATEAREA                          0.288 LAYER ME3 ;
 ANTENNAGATEAREA                          0.288 LAYER ME4 ;
 ANTENNADIFFAREA                          0.206 LAYER ME2 ;
 ANTENNADIFFAREA                          0.206 LAYER ME3 ;
 ANTENNADIFFAREA                          0.206 LAYER ME4 ;
 ANTENNAMAXAREACAR                        5.844 LAYER ME2 ;
 ANTENNAMAXAREACAR                        6.511 LAYER ME3 ;
 ANTENNAMAXAREACAR                        7.178 LAYER ME4 ;
END WEB0
PIN A1
  DIRECTION INPUT ;
 PORT
  LAYER ME3 ;
  RECT 193.456 0.000 193.776 0.720 ;
  LAYER ME2 ;
  RECT 193.456 0.000 193.776 0.720 ;
  LAYER ME1 ;
  RECT 193.456 0.000 193.776 0.720 ;
 END
 ANTENNAPARTIALMETALAREA                  3.547 LAYER ME2 ;
 ANTENNAGATEAREA                          0.144 LAYER ME2 ;
 ANTENNAGATEAREA                          0.144 LAYER ME3 ;
 ANTENNADIFFAREA                          0.218 LAYER ME2 ;
 ANTENNADIFFAREA                          0.218 LAYER ME3 ;
 ANTENNAMAXAREACAR                       27.235 LAYER ME2 ;
 ANTENNAMAXAREACAR                       28.835 LAYER ME3 ;
END A1
PIN A2
  DIRECTION INPUT ;
 PORT
  LAYER ME3 ;
  RECT 194.026 0.000 194.346 0.720 ;
  LAYER ME2 ;
  RECT 194.026 0.000 194.346 0.720 ;
  LAYER ME1 ;
  RECT 194.026 0.000 194.346 0.720 ;
 END
 ANTENNAPARTIALMETALAREA                  3.688 LAYER ME2 ;
 ANTENNAGATEAREA                          0.144 LAYER ME2 ;
 ANTENNAGATEAREA                          0.144 LAYER ME3 ;
 ANTENNADIFFAREA                          0.218 LAYER ME2 ;
 ANTENNADIFFAREA                          0.218 LAYER ME3 ;
 ANTENNAMAXAREACAR                       28.214 LAYER ME2 ;
 ANTENNAMAXAREACAR                       29.814 LAYER ME3 ;
END A2
PIN A3
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 187.208 0.000 187.528 0.720 ;
  LAYER ME3 ;
  RECT 187.208 0.000 187.528 0.720 ;
  LAYER ME2 ;
  RECT 187.208 0.000 187.528 0.720 ;
  LAYER ME1 ;
  RECT 187.208 0.000 187.528 0.720 ;
 END
 ANTENNAPARTIALMETALAREA                  4.391 LAYER ME2 ;
 ANTENNAGATEAREA                          0.180 LAYER ME2 ;
 ANTENNAGATEAREA                          0.180 LAYER ME3 ;
 ANTENNAGATEAREA                          0.180 LAYER ME4 ;
 ANTENNADIFFAREA                          0.218 LAYER ME2 ;
 ANTENNADIFFAREA                          0.218 LAYER ME3 ;
 ANTENNADIFFAREA                          0.218 LAYER ME4 ;
 ANTENNAMAXAREACAR                       27.451 LAYER ME2 ;
 ANTENNAMAXAREACAR                       28.731 LAYER ME3 ;
 ANTENNAMAXAREACAR                       30.011 LAYER ME4 ;
END A3
PIN A4
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 186.528 0.000 186.848 0.720 ;
  LAYER ME3 ;
  RECT 186.528 0.000 186.848 0.720 ;
  LAYER ME2 ;
  RECT 186.528 0.000 186.848 0.720 ;
  LAYER ME1 ;
  RECT 186.528 0.000 186.848 0.720 ;
 END
 ANTENNAPARTIALMETALAREA                  3.928 LAYER ME2 ;
 ANTENNAGATEAREA                          0.180 LAYER ME2 ;
 ANTENNAGATEAREA                          0.180 LAYER ME3 ;
 ANTENNAGATEAREA                          0.180 LAYER ME4 ;
 ANTENNADIFFAREA                          0.218 LAYER ME2 ;
 ANTENNADIFFAREA                          0.218 LAYER ME3 ;
 ANTENNADIFFAREA                          0.218 LAYER ME4 ;
 ANTENNAMAXAREACAR                       26.813 LAYER ME2 ;
 ANTENNAMAXAREACAR                       28.093 LAYER ME3 ;
 ANTENNAMAXAREACAR                       29.373 LAYER ME4 ;
END A4
PIN A0
  DIRECTION INPUT ;
 PORT
  LAYER ME3 ;
  RECT 204.042 0.000 204.362 0.662 ;
  LAYER ME2 ;
  RECT 204.042 0.000 204.362 0.662 ;
  LAYER ME1 ;
  RECT 204.042 0.000 204.362 0.662 ;
 END
 ANTENNAPARTIALMETALAREA                  5.907 LAYER ME2 ;
 ANTENNAGATEAREA                          0.108 LAYER ME2 ;
 ANTENNAGATEAREA                          0.108 LAYER ME3 ;
 ANTENNADIFFAREA                          0.218 LAYER ME2 ;
 ANTENNADIFFAREA                          0.218 LAYER ME3 ;
 ANTENNAMAXAREACAR                       58.521 LAYER ME2 ;
 ANTENNAMAXAREACAR                       60.482 LAYER ME3 ;
END A0
PIN DVSE
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 213.633 0.000 213.953 0.720 ;
  LAYER ME3 ;
  RECT 213.633 0.000 213.953 0.720 ;
  LAYER ME3 ;
  RECT 213.633 0.000 213.953 0.720 ;
  LAYER ME2 ;
  RECT 213.633 0.000 213.953 0.720 ;
  LAYER ME2 ;
  RECT 213.633 0.000 213.953 0.720 ;
  LAYER ME1 ;
  RECT 213.633 0.000 213.953 0.720 ;
  LAYER ME1 ;
  RECT 213.633 0.000 213.953 0.720 ;
 END
 ANTENNAPARTIALMETALAREA                  7.809 LAYER ME2 ;
 ANTENNAGATEAREA                          0.612 LAYER ME2 ;
 ANTENNAGATEAREA                          0.612 LAYER ME3 ;
 ANTENNAGATEAREA                          0.612 LAYER ME4 ;
 ANTENNADIFFAREA                          0.218 LAYER ME2 ;
 ANTENNADIFFAREA                          0.218 LAYER ME3 ;
 ANTENNADIFFAREA                          0.218 LAYER ME4 ;
 ANTENNAMAXAREACAR                       76.330 LAYER ME2 ;
 ANTENNAMAXAREACAR                       78.463 LAYER ME3 ;
 ANTENNAMAXAREACAR                       80.596 LAYER ME4 ;
END DVSE
PIN DVS3
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 213.113 0.000 213.433 0.720 ;
  LAYER ME3 ;
  RECT 213.113 0.000 213.433 0.720 ;
  LAYER ME3 ;
  RECT 213.113 0.000 213.433 0.720 ;
  LAYER ME2 ;
  RECT 213.113 0.000 213.433 0.720 ;
  LAYER ME2 ;
  RECT 213.113 0.000 213.433 0.720 ;
  LAYER ME1 ;
  RECT 213.113 0.000 213.433 0.720 ;
  LAYER ME1 ;
  RECT 213.113 0.000 213.433 0.720 ;
 END
 ANTENNAPARTIALMETALAREA                  6.179 LAYER ME2 ;
 ANTENNAGATEAREA                          0.108 LAYER ME2 ;
 ANTENNAGATEAREA                          0.108 LAYER ME3 ;
 ANTENNAGATEAREA                          0.108 LAYER ME4 ;
 ANTENNADIFFAREA                          0.218 LAYER ME2 ;
 ANTENNADIFFAREA                          0.218 LAYER ME3 ;
 ANTENNADIFFAREA                          0.218 LAYER ME4 ;
 ANTENNAMAXAREACAR                       68.823 LAYER ME2 ;
 ANTENNAMAXAREACAR                       70.956 LAYER ME3 ;
 ANTENNAMAXAREACAR                       73.089 LAYER ME4 ;
END DVS3
PIN DVS2
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 214.153 0.000 214.473 0.720 ;
  LAYER ME3 ;
  RECT 214.153 0.000 214.473 0.720 ;
  LAYER ME3 ;
  RECT 214.153 0.000 214.473 0.720 ;
  LAYER ME2 ;
  RECT 214.153 0.000 214.473 0.720 ;
  LAYER ME2 ;
  RECT 214.153 0.000 214.473 0.720 ;
  LAYER ME1 ;
  RECT 214.153 0.000 214.473 0.720 ;
  LAYER ME1 ;
  RECT 214.153 0.000 214.473 0.720 ;
 END
 ANTENNAPARTIALMETALAREA                  7.876 LAYER ME2 ;
 ANTENNAGATEAREA                          0.108 LAYER ME2 ;
 ANTENNAGATEAREA                          0.108 LAYER ME3 ;
 ANTENNAGATEAREA                          0.108 LAYER ME4 ;
 ANTENNADIFFAREA                          0.218 LAYER ME2 ;
 ANTENNADIFFAREA                          0.218 LAYER ME3 ;
 ANTENNADIFFAREA                          0.218 LAYER ME4 ;
 ANTENNAMAXAREACAR                       83.257 LAYER ME2 ;
 ANTENNAMAXAREACAR                       85.391 LAYER ME3 ;
 ANTENNAMAXAREACAR                       87.524 LAYER ME4 ;
END DVS2
PIN DVS1
  DIRECTION INPUT ;
 PORT
  LAYER ME3 ;
  RECT 210.497 0.000 210.817 0.720 ;
  LAYER ME2 ;
  RECT 210.497 0.000 210.817 0.720 ;
  LAYER ME1 ;
  RECT 210.497 0.000 210.817 0.720 ;
 END
 ANTENNAPARTIALMETALAREA                  6.247 LAYER ME2 ;
 ANTENNAGATEAREA                          0.108 LAYER ME2 ;
 ANTENNAGATEAREA                          0.108 LAYER ME3 ;
 ANTENNADIFFAREA                          0.218 LAYER ME2 ;
 ANTENNADIFFAREA                          0.218 LAYER ME3 ;
 ANTENNAMAXAREACAR                       69.294 LAYER ME2 ;
 ANTENNAMAXAREACAR                       71.427 LAYER ME3 ;
END DVS1
PIN DVS0
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 214.673 0.000 214.993 0.720 ;
  LAYER ME3 ;
  RECT 214.673 0.000 214.993 0.720 ;
  LAYER ME3 ;
  RECT 214.673 0.000 214.993 0.720 ;
  LAYER ME2 ;
  RECT 214.673 0.000 214.993 0.720 ;
  LAYER ME2 ;
  RECT 214.673 0.000 214.993 0.720 ;
  LAYER ME1 ;
  RECT 214.673 0.000 214.993 0.720 ;
  LAYER ME1 ;
  RECT 214.673 0.000 214.993 0.720 ;
 END
 ANTENNAPARTIALMETALAREA                  7.119 LAYER ME2 ;
 ANTENNAGATEAREA                          0.108 LAYER ME2 ;
 ANTENNAGATEAREA                          0.108 LAYER ME3 ;
 ANTENNAGATEAREA                          0.108 LAYER ME4 ;
 ANTENNADIFFAREA                          0.218 LAYER ME2 ;
 ANTENNADIFFAREA                          0.218 LAYER ME3 ;
 ANTENNADIFFAREA                          0.218 LAYER ME4 ;
 ANTENNAMAXAREACAR                       77.987 LAYER ME2 ;
 ANTENNAMAXAREACAR                       80.120 LAYER ME3 ;
 ANTENNAMAXAREACAR                       82.254 LAYER ME4 ;
END DVS0
PIN CK
  DIRECTION INPUT ;
 PORT
  LAYER ME3 ;
  RECT 206.581 0.000 206.901 0.720 ;
  LAYER ME2 ;
  RECT 206.581 0.000 206.901 0.720 ;
  LAYER ME1 ;
  RECT 206.581 0.000 206.901 0.720 ;
 END
 ANTENNAPARTIALMETALAREA                  5.257 LAYER ME2 ;
 ANTENNAPARTIALMETALAREA                  6.084 LAYER ME3 ;
 ANTENNAGATEAREA                          0.072 LAYER ME2 ;
 ANTENNAGATEAREA                          0.792 LAYER ME3 ;
 ANTENNADIFFAREA                          0.218 LAYER ME2 ;
 ANTENNADIFFAREA                          0.218 LAYER ME3 ;
 ANTENNAMAXAREACAR                       86.308 LAYER ME2 ;
 ANTENNAMAXAREACAR                      174.014 LAYER ME3 ;
END CK
PIN CSB
  DIRECTION INPUT ;
 PORT
  LAYER ME3 ;
  RECT 197.967 0.000 198.287 0.720 ;
  LAYER ME2 ;
  RECT 197.967 0.000 198.287 0.720 ;
  LAYER ME1 ;
  RECT 197.967 0.000 198.287 0.720 ;
 END
 ANTENNAPARTIALMETALAREA                  5.788 LAYER ME2 ;
 ANTENNAPARTIALMETALAREA                  6.164 LAYER ME3 ;
 ANTENNAGATEAREA                          2.508 LAYER ME2 ;
 ANTENNAGATEAREA                          3.228 LAYER ME3 ;
 ANTENNADIFFAREA                          0.218 LAYER ME2 ;
 ANTENNADIFFAREA                          0.218 LAYER ME3 ;
 ANTENNAMAXAREACAR                        3.046 LAYER ME2 ;
 ANTENNAMAXAREACAR                       32.772 LAYER ME3 ;
END CSB
PIN DI87
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 389.459 0.000 389.779 0.600 ;
  LAYER ME3 ;
  RECT 389.459 0.000 389.779 0.600 ;
  LAYER ME2 ;
  RECT 389.459 0.000 389.779 0.600 ;
  LAYER ME1 ;
  RECT 389.459 0.000 389.779 0.600 ;
 END
 ANTENNAPARTIALMETALAREA                  1.058 LAYER ME2 ;
 ANTENNAGATEAREA                          0.072 LAYER ME2 ;
 ANTENNAGATEAREA                          0.072 LAYER ME3 ;
 ANTENNAGATEAREA                          0.072 LAYER ME4 ;
 ANTENNADIFFAREA                          0.160 LAYER ME2 ;
 ANTENNADIFFAREA                          0.160 LAYER ME3 ;
 ANTENNADIFFAREA                          0.160 LAYER ME4 ;
 ANTENNAMAXAREACAR                       21.782 LAYER ME2 ;
 ANTENNAMAXAREACAR                       24.449 LAYER ME3 ;
 ANTENNAMAXAREACAR                       27.116 LAYER ME4 ;
END DI87
PIN DO87
  DIRECTION OUTPUT ;
 PORT
  LAYER ME4 ;
  RECT 388.897 0.000 389.217 0.600 ;
  LAYER ME3 ;
  RECT 388.897 0.000 389.217 0.600 ;
  LAYER ME2 ;
  RECT 388.897 0.000 389.217 0.600 ;
  LAYER ME1 ;
  RECT 388.897 0.000 389.217 0.600 ;
 END
 ANTENNAPARTIALMETALAREA                  5.273 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME3 ;
 ANTENNADIFFAREA                          1.293 LAYER ME4 ;
END DO87
PIN DI86
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 385.455 0.000 385.775 0.600 ;
  LAYER ME3 ;
  RECT 385.455 0.000 385.775 0.600 ;
  LAYER ME2 ;
  RECT 385.455 0.000 385.775 0.600 ;
  LAYER ME1 ;
  RECT 385.455 0.000 385.775 0.600 ;
 END
 ANTENNAPARTIALMETALAREA                  1.058 LAYER ME2 ;
 ANTENNAGATEAREA                          0.072 LAYER ME2 ;
 ANTENNAGATEAREA                          0.072 LAYER ME3 ;
 ANTENNAGATEAREA                          0.072 LAYER ME4 ;
 ANTENNADIFFAREA                          0.160 LAYER ME2 ;
 ANTENNADIFFAREA                          0.160 LAYER ME3 ;
 ANTENNADIFFAREA                          0.160 LAYER ME4 ;
 ANTENNAMAXAREACAR                       21.782 LAYER ME2 ;
 ANTENNAMAXAREACAR                       24.449 LAYER ME3 ;
 ANTENNAMAXAREACAR                       27.116 LAYER ME4 ;
END DI86
PIN DO86
  DIRECTION OUTPUT ;
 PORT
  LAYER ME4 ;
  RECT 384.893 0.000 385.213 0.600 ;
  LAYER ME3 ;
  RECT 384.893 0.000 385.213 0.600 ;
  LAYER ME2 ;
  RECT 384.893 0.000 385.213 0.600 ;
  LAYER ME1 ;
  RECT 384.893 0.000 385.213 0.600 ;
 END
 ANTENNAPARTIALMETALAREA                  5.273 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME3 ;
 ANTENNADIFFAREA                          1.293 LAYER ME4 ;
END DO86
PIN DI85
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 381.451 0.000 381.771 0.600 ;
  LAYER ME3 ;
  RECT 381.451 0.000 381.771 0.600 ;
  LAYER ME2 ;
  RECT 381.451 0.000 381.771 0.600 ;
  LAYER ME1 ;
  RECT 381.451 0.000 381.771 0.600 ;
 END
 ANTENNAPARTIALMETALAREA                  1.058 LAYER ME2 ;
 ANTENNAGATEAREA                          0.072 LAYER ME2 ;
 ANTENNAGATEAREA                          0.072 LAYER ME3 ;
 ANTENNAGATEAREA                          0.072 LAYER ME4 ;
 ANTENNADIFFAREA                          0.160 LAYER ME2 ;
 ANTENNADIFFAREA                          0.160 LAYER ME3 ;
 ANTENNADIFFAREA                          0.160 LAYER ME4 ;
 ANTENNAMAXAREACAR                       21.782 LAYER ME2 ;
 ANTENNAMAXAREACAR                       24.449 LAYER ME3 ;
 ANTENNAMAXAREACAR                       27.116 LAYER ME4 ;
END DI85
PIN DO85
  DIRECTION OUTPUT ;
 PORT
  LAYER ME4 ;
  RECT 380.889 0.000 381.209 0.600 ;
  LAYER ME3 ;
  RECT 380.889 0.000 381.209 0.600 ;
  LAYER ME2 ;
  RECT 380.889 0.000 381.209 0.600 ;
  LAYER ME1 ;
  RECT 380.889 0.000 381.209 0.600 ;
 END
 ANTENNAPARTIALMETALAREA                  5.273 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME3 ;
 ANTENNADIFFAREA                          1.293 LAYER ME4 ;
END DO85
PIN DI84
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 377.447 0.000 377.767 0.600 ;
  LAYER ME3 ;
  RECT 377.447 0.000 377.767 0.600 ;
  LAYER ME2 ;
  RECT 377.447 0.000 377.767 0.600 ;
  LAYER ME1 ;
  RECT 377.447 0.000 377.767 0.600 ;
 END
 ANTENNAPARTIALMETALAREA                  1.058 LAYER ME2 ;
 ANTENNAGATEAREA                          0.072 LAYER ME2 ;
 ANTENNAGATEAREA                          0.072 LAYER ME3 ;
 ANTENNAGATEAREA                          0.072 LAYER ME4 ;
 ANTENNADIFFAREA                          0.160 LAYER ME2 ;
 ANTENNADIFFAREA                          0.160 LAYER ME3 ;
 ANTENNADIFFAREA                          0.160 LAYER ME4 ;
 ANTENNAMAXAREACAR                       21.782 LAYER ME2 ;
 ANTENNAMAXAREACAR                       24.449 LAYER ME3 ;
 ANTENNAMAXAREACAR                       27.116 LAYER ME4 ;
END DI84
PIN DO84
  DIRECTION OUTPUT ;
 PORT
  LAYER ME4 ;
  RECT 376.885 0.000 377.205 0.600 ;
  LAYER ME3 ;
  RECT 376.885 0.000 377.205 0.600 ;
  LAYER ME2 ;
  RECT 376.885 0.000 377.205 0.600 ;
  LAYER ME1 ;
  RECT 376.885 0.000 377.205 0.600 ;
 END
 ANTENNAPARTIALMETALAREA                  5.273 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME3 ;
 ANTENNADIFFAREA                          1.293 LAYER ME4 ;
END DO84
PIN DI83
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 373.443 0.000 373.763 0.600 ;
  LAYER ME3 ;
  RECT 373.443 0.000 373.763 0.600 ;
  LAYER ME2 ;
  RECT 373.443 0.000 373.763 0.600 ;
  LAYER ME1 ;
  RECT 373.443 0.000 373.763 0.600 ;
 END
 ANTENNAPARTIALMETALAREA                  1.058 LAYER ME2 ;
 ANTENNAGATEAREA                          0.072 LAYER ME2 ;
 ANTENNAGATEAREA                          0.072 LAYER ME3 ;
 ANTENNAGATEAREA                          0.072 LAYER ME4 ;
 ANTENNADIFFAREA                          0.160 LAYER ME2 ;
 ANTENNADIFFAREA                          0.160 LAYER ME3 ;
 ANTENNADIFFAREA                          0.160 LAYER ME4 ;
 ANTENNAMAXAREACAR                       21.782 LAYER ME2 ;
 ANTENNAMAXAREACAR                       24.449 LAYER ME3 ;
 ANTENNAMAXAREACAR                       27.116 LAYER ME4 ;
END DI83
PIN DO83
  DIRECTION OUTPUT ;
 PORT
  LAYER ME4 ;
  RECT 372.881 0.000 373.201 0.600 ;
  LAYER ME3 ;
  RECT 372.881 0.000 373.201 0.600 ;
  LAYER ME2 ;
  RECT 372.881 0.000 373.201 0.600 ;
  LAYER ME1 ;
  RECT 372.881 0.000 373.201 0.600 ;
 END
 ANTENNAPARTIALMETALAREA                  5.273 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME3 ;
 ANTENNADIFFAREA                          1.293 LAYER ME4 ;
END DO83
PIN DI82
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 369.439 0.000 369.759 0.600 ;
  LAYER ME3 ;
  RECT 369.439 0.000 369.759 0.600 ;
  LAYER ME2 ;
  RECT 369.439 0.000 369.759 0.600 ;
  LAYER ME1 ;
  RECT 369.439 0.000 369.759 0.600 ;
 END
 ANTENNAPARTIALMETALAREA                  1.058 LAYER ME2 ;
 ANTENNAGATEAREA                          0.072 LAYER ME2 ;
 ANTENNAGATEAREA                          0.072 LAYER ME3 ;
 ANTENNAGATEAREA                          0.072 LAYER ME4 ;
 ANTENNADIFFAREA                          0.160 LAYER ME2 ;
 ANTENNADIFFAREA                          0.160 LAYER ME3 ;
 ANTENNADIFFAREA                          0.160 LAYER ME4 ;
 ANTENNAMAXAREACAR                       21.782 LAYER ME2 ;
 ANTENNAMAXAREACAR                       24.449 LAYER ME3 ;
 ANTENNAMAXAREACAR                       27.116 LAYER ME4 ;
END DI82
PIN DO82
  DIRECTION OUTPUT ;
 PORT
  LAYER ME4 ;
  RECT 368.877 0.000 369.197 0.600 ;
  LAYER ME3 ;
  RECT 368.877 0.000 369.197 0.600 ;
  LAYER ME2 ;
  RECT 368.877 0.000 369.197 0.600 ;
  LAYER ME1 ;
  RECT 368.877 0.000 369.197 0.600 ;
 END
 ANTENNAPARTIALMETALAREA                  5.273 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME3 ;
 ANTENNADIFFAREA                          1.293 LAYER ME4 ;
END DO82
PIN DI81
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 365.435 0.000 365.755 0.600 ;
  LAYER ME3 ;
  RECT 365.435 0.000 365.755 0.600 ;
  LAYER ME2 ;
  RECT 365.435 0.000 365.755 0.600 ;
  LAYER ME1 ;
  RECT 365.435 0.000 365.755 0.600 ;
 END
 ANTENNAPARTIALMETALAREA                  1.058 LAYER ME2 ;
 ANTENNAGATEAREA                          0.072 LAYER ME2 ;
 ANTENNAGATEAREA                          0.072 LAYER ME3 ;
 ANTENNAGATEAREA                          0.072 LAYER ME4 ;
 ANTENNADIFFAREA                          0.160 LAYER ME2 ;
 ANTENNADIFFAREA                          0.160 LAYER ME3 ;
 ANTENNADIFFAREA                          0.160 LAYER ME4 ;
 ANTENNAMAXAREACAR                       21.782 LAYER ME2 ;
 ANTENNAMAXAREACAR                       24.449 LAYER ME3 ;
 ANTENNAMAXAREACAR                       27.116 LAYER ME4 ;
END DI81
PIN DO81
  DIRECTION OUTPUT ;
 PORT
  LAYER ME4 ;
  RECT 364.873 0.000 365.193 0.600 ;
  LAYER ME3 ;
  RECT 364.873 0.000 365.193 0.600 ;
  LAYER ME2 ;
  RECT 364.873 0.000 365.193 0.600 ;
  LAYER ME1 ;
  RECT 364.873 0.000 365.193 0.600 ;
 END
 ANTENNAPARTIALMETALAREA                  5.273 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME3 ;
 ANTENNADIFFAREA                          1.293 LAYER ME4 ;
END DO81
PIN DI80
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 361.431 0.000 361.751 0.600 ;
  LAYER ME3 ;
  RECT 361.431 0.000 361.751 0.600 ;
  LAYER ME2 ;
  RECT 361.431 0.000 361.751 0.600 ;
  LAYER ME1 ;
  RECT 361.431 0.000 361.751 0.600 ;
 END
 ANTENNAPARTIALMETALAREA                  1.058 LAYER ME2 ;
 ANTENNAGATEAREA                          0.072 LAYER ME2 ;
 ANTENNAGATEAREA                          0.072 LAYER ME3 ;
 ANTENNAGATEAREA                          0.072 LAYER ME4 ;
 ANTENNADIFFAREA                          0.160 LAYER ME2 ;
 ANTENNADIFFAREA                          0.160 LAYER ME3 ;
 ANTENNADIFFAREA                          0.160 LAYER ME4 ;
 ANTENNAMAXAREACAR                       21.782 LAYER ME2 ;
 ANTENNAMAXAREACAR                       24.449 LAYER ME3 ;
 ANTENNAMAXAREACAR                       27.116 LAYER ME4 ;
END DI80
PIN DO80
  DIRECTION OUTPUT ;
 PORT
  LAYER ME4 ;
  RECT 360.869 0.000 361.189 0.600 ;
  LAYER ME3 ;
  RECT 360.869 0.000 361.189 0.600 ;
  LAYER ME2 ;
  RECT 360.869 0.000 361.189 0.600 ;
  LAYER ME1 ;
  RECT 360.869 0.000 361.189 0.600 ;
 END
 ANTENNAPARTIALMETALAREA                  5.273 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME3 ;
 ANTENNADIFFAREA                          1.293 LAYER ME4 ;
END DO80
PIN DI79
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 357.427 0.000 357.747 0.600 ;
  LAYER ME3 ;
  RECT 357.427 0.000 357.747 0.600 ;
  LAYER ME2 ;
  RECT 357.427 0.000 357.747 0.600 ;
  LAYER ME1 ;
  RECT 357.427 0.000 357.747 0.600 ;
 END
 ANTENNAPARTIALMETALAREA                  1.058 LAYER ME2 ;
 ANTENNAGATEAREA                          0.072 LAYER ME2 ;
 ANTENNAGATEAREA                          0.072 LAYER ME3 ;
 ANTENNAGATEAREA                          0.072 LAYER ME4 ;
 ANTENNADIFFAREA                          0.160 LAYER ME2 ;
 ANTENNADIFFAREA                          0.160 LAYER ME3 ;
 ANTENNADIFFAREA                          0.160 LAYER ME4 ;
 ANTENNAMAXAREACAR                       21.782 LAYER ME2 ;
 ANTENNAMAXAREACAR                       24.449 LAYER ME3 ;
 ANTENNAMAXAREACAR                       27.116 LAYER ME4 ;
END DI79
PIN DO79
  DIRECTION OUTPUT ;
 PORT
  LAYER ME4 ;
  RECT 356.865 0.000 357.185 0.600 ;
  LAYER ME3 ;
  RECT 356.865 0.000 357.185 0.600 ;
  LAYER ME2 ;
  RECT 356.865 0.000 357.185 0.600 ;
  LAYER ME1 ;
  RECT 356.865 0.000 357.185 0.600 ;
 END
 ANTENNAPARTIALMETALAREA                  5.273 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME3 ;
 ANTENNADIFFAREA                          1.293 LAYER ME4 ;
END DO79
PIN DI78
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 353.423 0.000 353.743 0.600 ;
  LAYER ME3 ;
  RECT 353.423 0.000 353.743 0.600 ;
  LAYER ME2 ;
  RECT 353.423 0.000 353.743 0.600 ;
  LAYER ME1 ;
  RECT 353.423 0.000 353.743 0.600 ;
 END
 ANTENNAPARTIALMETALAREA                  1.058 LAYER ME2 ;
 ANTENNAGATEAREA                          0.072 LAYER ME2 ;
 ANTENNAGATEAREA                          0.072 LAYER ME3 ;
 ANTENNAGATEAREA                          0.072 LAYER ME4 ;
 ANTENNADIFFAREA                          0.160 LAYER ME2 ;
 ANTENNADIFFAREA                          0.160 LAYER ME3 ;
 ANTENNADIFFAREA                          0.160 LAYER ME4 ;
 ANTENNAMAXAREACAR                       21.782 LAYER ME2 ;
 ANTENNAMAXAREACAR                       24.449 LAYER ME3 ;
 ANTENNAMAXAREACAR                       27.116 LAYER ME4 ;
END DI78
PIN DO78
  DIRECTION OUTPUT ;
 PORT
  LAYER ME4 ;
  RECT 352.861 0.000 353.181 0.600 ;
  LAYER ME3 ;
  RECT 352.861 0.000 353.181 0.600 ;
  LAYER ME2 ;
  RECT 352.861 0.000 353.181 0.600 ;
  LAYER ME1 ;
  RECT 352.861 0.000 353.181 0.600 ;
 END
 ANTENNAPARTIALMETALAREA                  5.273 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME3 ;
 ANTENNADIFFAREA                          1.293 LAYER ME4 ;
END DO78
PIN DI77
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 348.857 0.000 349.177 0.600 ;
  LAYER ME3 ;
  RECT 348.857 0.000 349.177 0.600 ;
  LAYER ME2 ;
  RECT 348.857 0.000 349.177 0.600 ;
  LAYER ME1 ;
  RECT 348.857 0.000 349.177 0.600 ;
 END
 ANTENNAPARTIALMETALAREA                  0.346 LAYER ME1 ;
 ANTENNAPARTIALMETALAREA                  1.466 LAYER ME2 ;
 ANTENNAPARTIALMETALAREA                  0.508 LAYER ME3 ;
 ANTENNAGATEAREA                          0.072 LAYER ME3 ;
 ANTENNAGATEAREA                          0.072 LAYER ME4 ;
 ANTENNADIFFAREA                          0.218 LAYER ME1 ;
 ANTENNADIFFAREA                          0.218 LAYER ME2 ;
 ANTENNADIFFAREA                          0.218 LAYER ME3 ;
 ANTENNADIFFAREA                          0.218 LAYER ME4 ;
 ANTENNAMAXAREACAR                       17.267 LAYER ME3 ;
 ANTENNAMAXAREACAR                       19.933 LAYER ME4 ;
END DI77
PIN DO77
  DIRECTION OUTPUT ;
 PORT
  LAYER ME4 ;
  RECT 349.419 0.000 349.739 0.600 ;
  LAYER ME3 ;
  RECT 349.419 0.000 349.739 0.600 ;
  LAYER ME2 ;
  RECT 349.419 0.000 349.739 0.600 ;
  LAYER ME1 ;
  RECT 349.419 0.000 349.739 0.600 ;
 END
 ANTENNAPARTIALMETALAREA                  5.602 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME3 ;
 ANTENNADIFFAREA                          1.293 LAYER ME4 ;
END DO77
PIN WEB7
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 347.417 0.000 347.737 0.600 ;
  LAYER ME3 ;
  RECT 347.417 0.000 347.737 0.600 ;
  LAYER ME2 ;
  RECT 347.417 0.000 347.737 0.600 ;
  LAYER ME1 ;
  RECT 347.417 0.000 347.737 0.600 ;
 END
 ANTENNAPARTIALMETALAREA                  1.036 LAYER ME2 ;
 ANTENNAGATEAREA                          0.288 LAYER ME2 ;
 ANTENNAGATEAREA                          0.288 LAYER ME3 ;
 ANTENNAGATEAREA                          0.288 LAYER ME4 ;
 ANTENNADIFFAREA                          0.206 LAYER ME2 ;
 ANTENNADIFFAREA                          0.206 LAYER ME3 ;
 ANTENNADIFFAREA                          0.206 LAYER ME4 ;
 ANTENNAMAXAREACAR                        5.844 LAYER ME2 ;
 ANTENNAMAXAREACAR                        6.511 LAYER ME3 ;
 ANTENNAMAXAREACAR                        7.178 LAYER ME4 ;
END WEB7
PIN DI76
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 345.415 0.000 345.735 0.600 ;
  LAYER ME3 ;
  RECT 345.415 0.000 345.735 0.600 ;
  LAYER ME2 ;
  RECT 345.415 0.000 345.735 0.600 ;
  LAYER ME1 ;
  RECT 345.415 0.000 345.735 0.600 ;
 END
 ANTENNAPARTIALMETALAREA                  1.058 LAYER ME2 ;
 ANTENNAGATEAREA                          0.072 LAYER ME2 ;
 ANTENNAGATEAREA                          0.072 LAYER ME3 ;
 ANTENNAGATEAREA                          0.072 LAYER ME4 ;
 ANTENNADIFFAREA                          0.160 LAYER ME2 ;
 ANTENNADIFFAREA                          0.160 LAYER ME3 ;
 ANTENNADIFFAREA                          0.160 LAYER ME4 ;
 ANTENNAMAXAREACAR                       21.782 LAYER ME2 ;
 ANTENNAMAXAREACAR                       24.449 LAYER ME3 ;
 ANTENNAMAXAREACAR                       27.116 LAYER ME4 ;
END DI76
PIN DO76
  DIRECTION OUTPUT ;
 PORT
  LAYER ME4 ;
  RECT 344.853 0.000 345.173 0.600 ;
  LAYER ME3 ;
  RECT 344.853 0.000 345.173 0.600 ;
  LAYER ME2 ;
  RECT 344.853 0.000 345.173 0.600 ;
  LAYER ME1 ;
  RECT 344.853 0.000 345.173 0.600 ;
 END
 ANTENNAPARTIALMETALAREA                  5.273 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME3 ;
 ANTENNADIFFAREA                          1.293 LAYER ME4 ;
END DO76
PIN DI75
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 341.411 0.000 341.731 0.600 ;
  LAYER ME3 ;
  RECT 341.411 0.000 341.731 0.600 ;
  LAYER ME2 ;
  RECT 341.411 0.000 341.731 0.600 ;
  LAYER ME1 ;
  RECT 341.411 0.000 341.731 0.600 ;
 END
 ANTENNAPARTIALMETALAREA                  1.058 LAYER ME2 ;
 ANTENNAGATEAREA                          0.072 LAYER ME2 ;
 ANTENNAGATEAREA                          0.072 LAYER ME3 ;
 ANTENNAGATEAREA                          0.072 LAYER ME4 ;
 ANTENNADIFFAREA                          0.160 LAYER ME2 ;
 ANTENNADIFFAREA                          0.160 LAYER ME3 ;
 ANTENNADIFFAREA                          0.160 LAYER ME4 ;
 ANTENNAMAXAREACAR                       21.782 LAYER ME2 ;
 ANTENNAMAXAREACAR                       24.449 LAYER ME3 ;
 ANTENNAMAXAREACAR                       27.116 LAYER ME4 ;
END DI75
PIN DO75
  DIRECTION OUTPUT ;
 PORT
  LAYER ME4 ;
  RECT 340.849 0.000 341.169 0.600 ;
  LAYER ME3 ;
  RECT 340.849 0.000 341.169 0.600 ;
  LAYER ME2 ;
  RECT 340.849 0.000 341.169 0.600 ;
  LAYER ME1 ;
  RECT 340.849 0.000 341.169 0.600 ;
 END
 ANTENNAPARTIALMETALAREA                  5.273 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME3 ;
 ANTENNADIFFAREA                          1.293 LAYER ME4 ;
END DO75
PIN DI74
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 337.407 0.000 337.727 0.600 ;
  LAYER ME3 ;
  RECT 337.407 0.000 337.727 0.600 ;
  LAYER ME2 ;
  RECT 337.407 0.000 337.727 0.600 ;
  LAYER ME1 ;
  RECT 337.407 0.000 337.727 0.600 ;
 END
 ANTENNAPARTIALMETALAREA                  1.058 LAYER ME2 ;
 ANTENNAGATEAREA                          0.072 LAYER ME2 ;
 ANTENNAGATEAREA                          0.072 LAYER ME3 ;
 ANTENNAGATEAREA                          0.072 LAYER ME4 ;
 ANTENNADIFFAREA                          0.160 LAYER ME2 ;
 ANTENNADIFFAREA                          0.160 LAYER ME3 ;
 ANTENNADIFFAREA                          0.160 LAYER ME4 ;
 ANTENNAMAXAREACAR                       21.782 LAYER ME2 ;
 ANTENNAMAXAREACAR                       24.449 LAYER ME3 ;
 ANTENNAMAXAREACAR                       27.116 LAYER ME4 ;
END DI74
PIN DO74
  DIRECTION OUTPUT ;
 PORT
  LAYER ME4 ;
  RECT 336.845 0.000 337.165 0.600 ;
  LAYER ME3 ;
  RECT 336.845 0.000 337.165 0.600 ;
  LAYER ME2 ;
  RECT 336.845 0.000 337.165 0.600 ;
  LAYER ME1 ;
  RECT 336.845 0.000 337.165 0.600 ;
 END
 ANTENNAPARTIALMETALAREA                  5.273 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME3 ;
 ANTENNADIFFAREA                          1.293 LAYER ME4 ;
END DO74
PIN DI73
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 333.403 0.000 333.723 0.600 ;
  LAYER ME3 ;
  RECT 333.403 0.000 333.723 0.600 ;
  LAYER ME2 ;
  RECT 333.403 0.000 333.723 0.600 ;
  LAYER ME1 ;
  RECT 333.403 0.000 333.723 0.600 ;
 END
 ANTENNAPARTIALMETALAREA                  1.058 LAYER ME2 ;
 ANTENNAGATEAREA                          0.072 LAYER ME2 ;
 ANTENNAGATEAREA                          0.072 LAYER ME3 ;
 ANTENNAGATEAREA                          0.072 LAYER ME4 ;
 ANTENNADIFFAREA                          0.160 LAYER ME2 ;
 ANTENNADIFFAREA                          0.160 LAYER ME3 ;
 ANTENNADIFFAREA                          0.160 LAYER ME4 ;
 ANTENNAMAXAREACAR                       21.782 LAYER ME2 ;
 ANTENNAMAXAREACAR                       24.449 LAYER ME3 ;
 ANTENNAMAXAREACAR                       27.116 LAYER ME4 ;
END DI73
PIN DO73
  DIRECTION OUTPUT ;
 PORT
  LAYER ME4 ;
  RECT 332.841 0.000 333.161 0.600 ;
  LAYER ME3 ;
  RECT 332.841 0.000 333.161 0.600 ;
  LAYER ME2 ;
  RECT 332.841 0.000 333.161 0.600 ;
  LAYER ME1 ;
  RECT 332.841 0.000 333.161 0.600 ;
 END
 ANTENNAPARTIALMETALAREA                  5.273 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME3 ;
 ANTENNADIFFAREA                          1.293 LAYER ME4 ;
END DO73
PIN DI72
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 329.399 0.000 329.719 0.600 ;
  LAYER ME3 ;
  RECT 329.399 0.000 329.719 0.600 ;
  LAYER ME2 ;
  RECT 329.399 0.000 329.719 0.600 ;
  LAYER ME1 ;
  RECT 329.399 0.000 329.719 0.600 ;
 END
 ANTENNAPARTIALMETALAREA                  1.058 LAYER ME2 ;
 ANTENNAGATEAREA                          0.072 LAYER ME2 ;
 ANTENNAGATEAREA                          0.072 LAYER ME3 ;
 ANTENNAGATEAREA                          0.072 LAYER ME4 ;
 ANTENNADIFFAREA                          0.160 LAYER ME2 ;
 ANTENNADIFFAREA                          0.160 LAYER ME3 ;
 ANTENNADIFFAREA                          0.160 LAYER ME4 ;
 ANTENNAMAXAREACAR                       21.782 LAYER ME2 ;
 ANTENNAMAXAREACAR                       24.449 LAYER ME3 ;
 ANTENNAMAXAREACAR                       27.116 LAYER ME4 ;
END DI72
PIN DO72
  DIRECTION OUTPUT ;
 PORT
  LAYER ME4 ;
  RECT 328.837 0.000 329.157 0.600 ;
  LAYER ME3 ;
  RECT 328.837 0.000 329.157 0.600 ;
  LAYER ME2 ;
  RECT 328.837 0.000 329.157 0.600 ;
  LAYER ME1 ;
  RECT 328.837 0.000 329.157 0.600 ;
 END
 ANTENNAPARTIALMETALAREA                  5.273 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME3 ;
 ANTENNADIFFAREA                          1.293 LAYER ME4 ;
END DO72
PIN DI71
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 325.395 0.000 325.715 0.600 ;
  LAYER ME3 ;
  RECT 325.395 0.000 325.715 0.600 ;
  LAYER ME2 ;
  RECT 325.395 0.000 325.715 0.600 ;
  LAYER ME1 ;
  RECT 325.395 0.000 325.715 0.600 ;
 END
 ANTENNAPARTIALMETALAREA                  1.058 LAYER ME2 ;
 ANTENNAGATEAREA                          0.072 LAYER ME2 ;
 ANTENNAGATEAREA                          0.072 LAYER ME3 ;
 ANTENNAGATEAREA                          0.072 LAYER ME4 ;
 ANTENNADIFFAREA                          0.160 LAYER ME2 ;
 ANTENNADIFFAREA                          0.160 LAYER ME3 ;
 ANTENNADIFFAREA                          0.160 LAYER ME4 ;
 ANTENNAMAXAREACAR                       21.782 LAYER ME2 ;
 ANTENNAMAXAREACAR                       24.449 LAYER ME3 ;
 ANTENNAMAXAREACAR                       27.116 LAYER ME4 ;
END DI71
PIN DO71
  DIRECTION OUTPUT ;
 PORT
  LAYER ME4 ;
  RECT 324.833 0.000 325.153 0.600 ;
  LAYER ME3 ;
  RECT 324.833 0.000 325.153 0.600 ;
  LAYER ME2 ;
  RECT 324.833 0.000 325.153 0.600 ;
  LAYER ME1 ;
  RECT 324.833 0.000 325.153 0.600 ;
 END
 ANTENNAPARTIALMETALAREA                  5.273 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME3 ;
 ANTENNADIFFAREA                          1.293 LAYER ME4 ;
END DO71
PIN DI70
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 321.391 0.000 321.711 0.600 ;
  LAYER ME3 ;
  RECT 321.391 0.000 321.711 0.600 ;
  LAYER ME2 ;
  RECT 321.391 0.000 321.711 0.600 ;
  LAYER ME1 ;
  RECT 321.391 0.000 321.711 0.600 ;
 END
 ANTENNAPARTIALMETALAREA                  1.058 LAYER ME2 ;
 ANTENNAGATEAREA                          0.072 LAYER ME2 ;
 ANTENNAGATEAREA                          0.072 LAYER ME3 ;
 ANTENNAGATEAREA                          0.072 LAYER ME4 ;
 ANTENNADIFFAREA                          0.160 LAYER ME2 ;
 ANTENNADIFFAREA                          0.160 LAYER ME3 ;
 ANTENNADIFFAREA                          0.160 LAYER ME4 ;
 ANTENNAMAXAREACAR                       21.782 LAYER ME2 ;
 ANTENNAMAXAREACAR                       24.449 LAYER ME3 ;
 ANTENNAMAXAREACAR                       27.116 LAYER ME4 ;
END DI70
PIN DO70
  DIRECTION OUTPUT ;
 PORT
  LAYER ME4 ;
  RECT 320.829 0.000 321.149 0.600 ;
  LAYER ME3 ;
  RECT 320.829 0.000 321.149 0.600 ;
  LAYER ME2 ;
  RECT 320.829 0.000 321.149 0.600 ;
  LAYER ME1 ;
  RECT 320.829 0.000 321.149 0.600 ;
 END
 ANTENNAPARTIALMETALAREA                  5.273 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME3 ;
 ANTENNADIFFAREA                          1.293 LAYER ME4 ;
END DO70
PIN DI69
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 317.387 0.000 317.707 0.600 ;
  LAYER ME3 ;
  RECT 317.387 0.000 317.707 0.600 ;
  LAYER ME2 ;
  RECT 317.387 0.000 317.707 0.600 ;
  LAYER ME1 ;
  RECT 317.387 0.000 317.707 0.600 ;
 END
 ANTENNAPARTIALMETALAREA                  1.058 LAYER ME2 ;
 ANTENNAGATEAREA                          0.072 LAYER ME2 ;
 ANTENNAGATEAREA                          0.072 LAYER ME3 ;
 ANTENNAGATEAREA                          0.072 LAYER ME4 ;
 ANTENNADIFFAREA                          0.160 LAYER ME2 ;
 ANTENNADIFFAREA                          0.160 LAYER ME3 ;
 ANTENNADIFFAREA                          0.160 LAYER ME4 ;
 ANTENNAMAXAREACAR                       21.782 LAYER ME2 ;
 ANTENNAMAXAREACAR                       24.449 LAYER ME3 ;
 ANTENNAMAXAREACAR                       27.116 LAYER ME4 ;
END DI69
PIN DO69
  DIRECTION OUTPUT ;
 PORT
  LAYER ME4 ;
  RECT 316.825 0.000 317.145 0.600 ;
  LAYER ME3 ;
  RECT 316.825 0.000 317.145 0.600 ;
  LAYER ME2 ;
  RECT 316.825 0.000 317.145 0.600 ;
  LAYER ME1 ;
  RECT 316.825 0.000 317.145 0.600 ;
 END
 ANTENNAPARTIALMETALAREA                  5.273 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME3 ;
 ANTENNADIFFAREA                          1.293 LAYER ME4 ;
END DO69
PIN DI68
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 313.383 0.000 313.703 0.600 ;
  LAYER ME3 ;
  RECT 313.383 0.000 313.703 0.600 ;
  LAYER ME2 ;
  RECT 313.383 0.000 313.703 0.600 ;
  LAYER ME1 ;
  RECT 313.383 0.000 313.703 0.600 ;
 END
 ANTENNAPARTIALMETALAREA                  1.058 LAYER ME2 ;
 ANTENNAGATEAREA                          0.072 LAYER ME2 ;
 ANTENNAGATEAREA                          0.072 LAYER ME3 ;
 ANTENNAGATEAREA                          0.072 LAYER ME4 ;
 ANTENNADIFFAREA                          0.160 LAYER ME2 ;
 ANTENNADIFFAREA                          0.160 LAYER ME3 ;
 ANTENNADIFFAREA                          0.160 LAYER ME4 ;
 ANTENNAMAXAREACAR                       21.782 LAYER ME2 ;
 ANTENNAMAXAREACAR                       24.449 LAYER ME3 ;
 ANTENNAMAXAREACAR                       27.116 LAYER ME4 ;
END DI68
PIN DO68
  DIRECTION OUTPUT ;
 PORT
  LAYER ME4 ;
  RECT 312.821 0.000 313.141 0.600 ;
  LAYER ME3 ;
  RECT 312.821 0.000 313.141 0.600 ;
  LAYER ME2 ;
  RECT 312.821 0.000 313.141 0.600 ;
  LAYER ME1 ;
  RECT 312.821 0.000 313.141 0.600 ;
 END
 ANTENNAPARTIALMETALAREA                  5.273 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME3 ;
 ANTENNADIFFAREA                          1.293 LAYER ME4 ;
END DO68
PIN DI67
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 309.379 0.000 309.699 0.600 ;
  LAYER ME3 ;
  RECT 309.379 0.000 309.699 0.600 ;
  LAYER ME2 ;
  RECT 309.379 0.000 309.699 0.600 ;
  LAYER ME1 ;
  RECT 309.379 0.000 309.699 0.600 ;
 END
 ANTENNAPARTIALMETALAREA                  1.058 LAYER ME2 ;
 ANTENNAGATEAREA                          0.072 LAYER ME2 ;
 ANTENNAGATEAREA                          0.072 LAYER ME3 ;
 ANTENNAGATEAREA                          0.072 LAYER ME4 ;
 ANTENNADIFFAREA                          0.160 LAYER ME2 ;
 ANTENNADIFFAREA                          0.160 LAYER ME3 ;
 ANTENNADIFFAREA                          0.160 LAYER ME4 ;
 ANTENNAMAXAREACAR                       21.782 LAYER ME2 ;
 ANTENNAMAXAREACAR                       24.449 LAYER ME3 ;
 ANTENNAMAXAREACAR                       27.116 LAYER ME4 ;
END DI67
PIN DO67
  DIRECTION OUTPUT ;
 PORT
  LAYER ME4 ;
  RECT 308.817 0.000 309.137 0.600 ;
  LAYER ME3 ;
  RECT 308.817 0.000 309.137 0.600 ;
  LAYER ME2 ;
  RECT 308.817 0.000 309.137 0.600 ;
  LAYER ME1 ;
  RECT 308.817 0.000 309.137 0.600 ;
 END
 ANTENNAPARTIALMETALAREA                  5.273 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME3 ;
 ANTENNADIFFAREA                          1.293 LAYER ME4 ;
END DO67
PIN DI66
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 304.813 0.000 305.133 0.600 ;
  LAYER ME3 ;
  RECT 304.813 0.000 305.133 0.600 ;
  LAYER ME2 ;
  RECT 304.813 0.000 305.133 0.600 ;
  LAYER ME1 ;
  RECT 304.813 0.000 305.133 0.600 ;
 END
 ANTENNAPARTIALMETALAREA                  0.346 LAYER ME1 ;
 ANTENNAPARTIALMETALAREA                  1.466 LAYER ME2 ;
 ANTENNAPARTIALMETALAREA                  0.508 LAYER ME3 ;
 ANTENNAGATEAREA                          0.072 LAYER ME3 ;
 ANTENNAGATEAREA                          0.072 LAYER ME4 ;
 ANTENNADIFFAREA                          0.218 LAYER ME1 ;
 ANTENNADIFFAREA                          0.218 LAYER ME2 ;
 ANTENNADIFFAREA                          0.218 LAYER ME3 ;
 ANTENNADIFFAREA                          0.218 LAYER ME4 ;
 ANTENNAMAXAREACAR                       17.267 LAYER ME3 ;
 ANTENNAMAXAREACAR                       19.933 LAYER ME4 ;
END DI66
PIN DO66
  DIRECTION OUTPUT ;
 PORT
  LAYER ME4 ;
  RECT 305.375 0.000 305.695 0.600 ;
  LAYER ME3 ;
  RECT 305.375 0.000 305.695 0.600 ;
  LAYER ME2 ;
  RECT 305.375 0.000 305.695 0.600 ;
  LAYER ME1 ;
  RECT 305.375 0.000 305.695 0.600 ;
 END
 ANTENNAPARTIALMETALAREA                  5.602 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME3 ;
 ANTENNADIFFAREA                          1.293 LAYER ME4 ;
END DO66
PIN WEB6
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 303.373 0.000 303.693 0.600 ;
  LAYER ME3 ;
  RECT 303.373 0.000 303.693 0.600 ;
  LAYER ME2 ;
  RECT 303.373 0.000 303.693 0.600 ;
  LAYER ME1 ;
  RECT 303.373 0.000 303.693 0.600 ;
 END
 ANTENNAPARTIALMETALAREA                  1.036 LAYER ME2 ;
 ANTENNAGATEAREA                          0.288 LAYER ME2 ;
 ANTENNAGATEAREA                          0.288 LAYER ME3 ;
 ANTENNAGATEAREA                          0.288 LAYER ME4 ;
 ANTENNADIFFAREA                          0.206 LAYER ME2 ;
 ANTENNADIFFAREA                          0.206 LAYER ME3 ;
 ANTENNADIFFAREA                          0.206 LAYER ME4 ;
 ANTENNAMAXAREACAR                        5.844 LAYER ME2 ;
 ANTENNAMAXAREACAR                        6.511 LAYER ME3 ;
 ANTENNAMAXAREACAR                        7.178 LAYER ME4 ;
END WEB6
PIN DI65
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 301.371 0.000 301.691 0.600 ;
  LAYER ME3 ;
  RECT 301.371 0.000 301.691 0.600 ;
  LAYER ME2 ;
  RECT 301.371 0.000 301.691 0.600 ;
  LAYER ME1 ;
  RECT 301.371 0.000 301.691 0.600 ;
 END
 ANTENNAPARTIALMETALAREA                  1.058 LAYER ME2 ;
 ANTENNAGATEAREA                          0.072 LAYER ME2 ;
 ANTENNAGATEAREA                          0.072 LAYER ME3 ;
 ANTENNAGATEAREA                          0.072 LAYER ME4 ;
 ANTENNADIFFAREA                          0.160 LAYER ME2 ;
 ANTENNADIFFAREA                          0.160 LAYER ME3 ;
 ANTENNADIFFAREA                          0.160 LAYER ME4 ;
 ANTENNAMAXAREACAR                       21.782 LAYER ME2 ;
 ANTENNAMAXAREACAR                       24.449 LAYER ME3 ;
 ANTENNAMAXAREACAR                       27.116 LAYER ME4 ;
END DI65
PIN DO65
  DIRECTION OUTPUT ;
 PORT
  LAYER ME4 ;
  RECT 300.809 0.000 301.129 0.600 ;
  LAYER ME3 ;
  RECT 300.809 0.000 301.129 0.600 ;
  LAYER ME2 ;
  RECT 300.809 0.000 301.129 0.600 ;
  LAYER ME1 ;
  RECT 300.809 0.000 301.129 0.600 ;
 END
 ANTENNAPARTIALMETALAREA                  5.273 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME3 ;
 ANTENNADIFFAREA                          1.293 LAYER ME4 ;
END DO65
PIN DI64
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 297.367 0.000 297.687 0.600 ;
  LAYER ME3 ;
  RECT 297.367 0.000 297.687 0.600 ;
  LAYER ME2 ;
  RECT 297.367 0.000 297.687 0.600 ;
  LAYER ME1 ;
  RECT 297.367 0.000 297.687 0.600 ;
 END
 ANTENNAPARTIALMETALAREA                  1.058 LAYER ME2 ;
 ANTENNAGATEAREA                          0.072 LAYER ME2 ;
 ANTENNAGATEAREA                          0.072 LAYER ME3 ;
 ANTENNAGATEAREA                          0.072 LAYER ME4 ;
 ANTENNADIFFAREA                          0.160 LAYER ME2 ;
 ANTENNADIFFAREA                          0.160 LAYER ME3 ;
 ANTENNADIFFAREA                          0.160 LAYER ME4 ;
 ANTENNAMAXAREACAR                       21.782 LAYER ME2 ;
 ANTENNAMAXAREACAR                       24.449 LAYER ME3 ;
 ANTENNAMAXAREACAR                       27.116 LAYER ME4 ;
END DI64
PIN DO64
  DIRECTION OUTPUT ;
 PORT
  LAYER ME4 ;
  RECT 296.805 0.000 297.125 0.600 ;
  LAYER ME3 ;
  RECT 296.805 0.000 297.125 0.600 ;
  LAYER ME2 ;
  RECT 296.805 0.000 297.125 0.600 ;
  LAYER ME1 ;
  RECT 296.805 0.000 297.125 0.600 ;
 END
 ANTENNAPARTIALMETALAREA                  5.273 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME3 ;
 ANTENNADIFFAREA                          1.293 LAYER ME4 ;
END DO64
PIN DI63
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 293.363 0.000 293.683 0.600 ;
  LAYER ME3 ;
  RECT 293.363 0.000 293.683 0.600 ;
  LAYER ME2 ;
  RECT 293.363 0.000 293.683 0.600 ;
  LAYER ME1 ;
  RECT 293.363 0.000 293.683 0.600 ;
 END
 ANTENNAPARTIALMETALAREA                  1.058 LAYER ME2 ;
 ANTENNAGATEAREA                          0.072 LAYER ME2 ;
 ANTENNAGATEAREA                          0.072 LAYER ME3 ;
 ANTENNAGATEAREA                          0.072 LAYER ME4 ;
 ANTENNADIFFAREA                          0.160 LAYER ME2 ;
 ANTENNADIFFAREA                          0.160 LAYER ME3 ;
 ANTENNADIFFAREA                          0.160 LAYER ME4 ;
 ANTENNAMAXAREACAR                       21.782 LAYER ME2 ;
 ANTENNAMAXAREACAR                       24.449 LAYER ME3 ;
 ANTENNAMAXAREACAR                       27.116 LAYER ME4 ;
END DI63
PIN DO63
  DIRECTION OUTPUT ;
 PORT
  LAYER ME4 ;
  RECT 292.801 0.000 293.121 0.600 ;
  LAYER ME3 ;
  RECT 292.801 0.000 293.121 0.600 ;
  LAYER ME2 ;
  RECT 292.801 0.000 293.121 0.600 ;
  LAYER ME1 ;
  RECT 292.801 0.000 293.121 0.600 ;
 END
 ANTENNAPARTIALMETALAREA                  5.273 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME3 ;
 ANTENNADIFFAREA                          1.293 LAYER ME4 ;
END DO63
PIN DI62
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 289.359 0.000 289.679 0.600 ;
  LAYER ME3 ;
  RECT 289.359 0.000 289.679 0.600 ;
  LAYER ME2 ;
  RECT 289.359 0.000 289.679 0.600 ;
  LAYER ME1 ;
  RECT 289.359 0.000 289.679 0.600 ;
 END
 ANTENNAPARTIALMETALAREA                  1.058 LAYER ME2 ;
 ANTENNAGATEAREA                          0.072 LAYER ME2 ;
 ANTENNAGATEAREA                          0.072 LAYER ME3 ;
 ANTENNAGATEAREA                          0.072 LAYER ME4 ;
 ANTENNADIFFAREA                          0.160 LAYER ME2 ;
 ANTENNADIFFAREA                          0.160 LAYER ME3 ;
 ANTENNADIFFAREA                          0.160 LAYER ME4 ;
 ANTENNAMAXAREACAR                       21.782 LAYER ME2 ;
 ANTENNAMAXAREACAR                       24.449 LAYER ME3 ;
 ANTENNAMAXAREACAR                       27.116 LAYER ME4 ;
END DI62
PIN DO62
  DIRECTION OUTPUT ;
 PORT
  LAYER ME4 ;
  RECT 288.797 0.000 289.117 0.600 ;
  LAYER ME3 ;
  RECT 288.797 0.000 289.117 0.600 ;
  LAYER ME2 ;
  RECT 288.797 0.000 289.117 0.600 ;
  LAYER ME1 ;
  RECT 288.797 0.000 289.117 0.600 ;
 END
 ANTENNAPARTIALMETALAREA                  5.273 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME3 ;
 ANTENNADIFFAREA                          1.293 LAYER ME4 ;
END DO62
PIN DI61
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 285.355 0.000 285.675 0.600 ;
  LAYER ME3 ;
  RECT 285.355 0.000 285.675 0.600 ;
  LAYER ME2 ;
  RECT 285.355 0.000 285.675 0.600 ;
  LAYER ME1 ;
  RECT 285.355 0.000 285.675 0.600 ;
 END
 ANTENNAPARTIALMETALAREA                  1.058 LAYER ME2 ;
 ANTENNAGATEAREA                          0.072 LAYER ME2 ;
 ANTENNAGATEAREA                          0.072 LAYER ME3 ;
 ANTENNAGATEAREA                          0.072 LAYER ME4 ;
 ANTENNADIFFAREA                          0.160 LAYER ME2 ;
 ANTENNADIFFAREA                          0.160 LAYER ME3 ;
 ANTENNADIFFAREA                          0.160 LAYER ME4 ;
 ANTENNAMAXAREACAR                       21.782 LAYER ME2 ;
 ANTENNAMAXAREACAR                       24.449 LAYER ME3 ;
 ANTENNAMAXAREACAR                       27.116 LAYER ME4 ;
END DI61
PIN DO61
  DIRECTION OUTPUT ;
 PORT
  LAYER ME4 ;
  RECT 284.793 0.000 285.113 0.600 ;
  LAYER ME3 ;
  RECT 284.793 0.000 285.113 0.600 ;
  LAYER ME2 ;
  RECT 284.793 0.000 285.113 0.600 ;
  LAYER ME1 ;
  RECT 284.793 0.000 285.113 0.600 ;
 END
 ANTENNAPARTIALMETALAREA                  5.273 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME3 ;
 ANTENNADIFFAREA                          1.293 LAYER ME4 ;
END DO61
PIN DI60
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 281.351 0.000 281.671 0.600 ;
  LAYER ME3 ;
  RECT 281.351 0.000 281.671 0.600 ;
  LAYER ME2 ;
  RECT 281.351 0.000 281.671 0.600 ;
  LAYER ME1 ;
  RECT 281.351 0.000 281.671 0.600 ;
 END
 ANTENNAPARTIALMETALAREA                  1.058 LAYER ME2 ;
 ANTENNAGATEAREA                          0.072 LAYER ME2 ;
 ANTENNAGATEAREA                          0.072 LAYER ME3 ;
 ANTENNAGATEAREA                          0.072 LAYER ME4 ;
 ANTENNADIFFAREA                          0.160 LAYER ME2 ;
 ANTENNADIFFAREA                          0.160 LAYER ME3 ;
 ANTENNADIFFAREA                          0.160 LAYER ME4 ;
 ANTENNAMAXAREACAR                       21.782 LAYER ME2 ;
 ANTENNAMAXAREACAR                       24.449 LAYER ME3 ;
 ANTENNAMAXAREACAR                       27.116 LAYER ME4 ;
END DI60
PIN DO60
  DIRECTION OUTPUT ;
 PORT
  LAYER ME4 ;
  RECT 280.789 0.000 281.109 0.600 ;
  LAYER ME3 ;
  RECT 280.789 0.000 281.109 0.600 ;
  LAYER ME2 ;
  RECT 280.789 0.000 281.109 0.600 ;
  LAYER ME1 ;
  RECT 280.789 0.000 281.109 0.600 ;
 END
 ANTENNAPARTIALMETALAREA                  5.273 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME3 ;
 ANTENNADIFFAREA                          1.293 LAYER ME4 ;
END DO60
PIN DI59
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 277.347 0.000 277.667 0.600 ;
  LAYER ME3 ;
  RECT 277.347 0.000 277.667 0.600 ;
  LAYER ME2 ;
  RECT 277.347 0.000 277.667 0.600 ;
  LAYER ME1 ;
  RECT 277.347 0.000 277.667 0.600 ;
 END
 ANTENNAPARTIALMETALAREA                  1.058 LAYER ME2 ;
 ANTENNAGATEAREA                          0.072 LAYER ME2 ;
 ANTENNAGATEAREA                          0.072 LAYER ME3 ;
 ANTENNAGATEAREA                          0.072 LAYER ME4 ;
 ANTENNADIFFAREA                          0.160 LAYER ME2 ;
 ANTENNADIFFAREA                          0.160 LAYER ME3 ;
 ANTENNADIFFAREA                          0.160 LAYER ME4 ;
 ANTENNAMAXAREACAR                       21.782 LAYER ME2 ;
 ANTENNAMAXAREACAR                       24.449 LAYER ME3 ;
 ANTENNAMAXAREACAR                       27.116 LAYER ME4 ;
END DI59
PIN DO59
  DIRECTION OUTPUT ;
 PORT
  LAYER ME4 ;
  RECT 276.785 0.000 277.105 0.600 ;
  LAYER ME3 ;
  RECT 276.785 0.000 277.105 0.600 ;
  LAYER ME2 ;
  RECT 276.785 0.000 277.105 0.600 ;
  LAYER ME1 ;
  RECT 276.785 0.000 277.105 0.600 ;
 END
 ANTENNAPARTIALMETALAREA                  5.273 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME3 ;
 ANTENNADIFFAREA                          1.293 LAYER ME4 ;
END DO59
PIN DI58
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 273.343 0.000 273.663 0.600 ;
  LAYER ME3 ;
  RECT 273.343 0.000 273.663 0.600 ;
  LAYER ME2 ;
  RECT 273.343 0.000 273.663 0.600 ;
  LAYER ME1 ;
  RECT 273.343 0.000 273.663 0.600 ;
 END
 ANTENNAPARTIALMETALAREA                  1.058 LAYER ME2 ;
 ANTENNAGATEAREA                          0.072 LAYER ME2 ;
 ANTENNAGATEAREA                          0.072 LAYER ME3 ;
 ANTENNAGATEAREA                          0.072 LAYER ME4 ;
 ANTENNADIFFAREA                          0.160 LAYER ME2 ;
 ANTENNADIFFAREA                          0.160 LAYER ME3 ;
 ANTENNADIFFAREA                          0.160 LAYER ME4 ;
 ANTENNAMAXAREACAR                       21.782 LAYER ME2 ;
 ANTENNAMAXAREACAR                       24.449 LAYER ME3 ;
 ANTENNAMAXAREACAR                       27.116 LAYER ME4 ;
END DI58
PIN DO58
  DIRECTION OUTPUT ;
 PORT
  LAYER ME4 ;
  RECT 272.781 0.000 273.101 0.600 ;
  LAYER ME3 ;
  RECT 272.781 0.000 273.101 0.600 ;
  LAYER ME2 ;
  RECT 272.781 0.000 273.101 0.600 ;
  LAYER ME1 ;
  RECT 272.781 0.000 273.101 0.600 ;
 END
 ANTENNAPARTIALMETALAREA                  5.273 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME3 ;
 ANTENNADIFFAREA                          1.293 LAYER ME4 ;
END DO58
PIN DI57
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 269.339 0.000 269.659 0.600 ;
  LAYER ME3 ;
  RECT 269.339 0.000 269.659 0.600 ;
  LAYER ME2 ;
  RECT 269.339 0.000 269.659 0.600 ;
  LAYER ME1 ;
  RECT 269.339 0.000 269.659 0.600 ;
 END
 ANTENNAPARTIALMETALAREA                  1.058 LAYER ME2 ;
 ANTENNAGATEAREA                          0.072 LAYER ME2 ;
 ANTENNAGATEAREA                          0.072 LAYER ME3 ;
 ANTENNAGATEAREA                          0.072 LAYER ME4 ;
 ANTENNADIFFAREA                          0.160 LAYER ME2 ;
 ANTENNADIFFAREA                          0.160 LAYER ME3 ;
 ANTENNADIFFAREA                          0.160 LAYER ME4 ;
 ANTENNAMAXAREACAR                       21.782 LAYER ME2 ;
 ANTENNAMAXAREACAR                       24.449 LAYER ME3 ;
 ANTENNAMAXAREACAR                       27.116 LAYER ME4 ;
END DI57
PIN DO57
  DIRECTION OUTPUT ;
 PORT
  LAYER ME4 ;
  RECT 268.777 0.000 269.097 0.600 ;
  LAYER ME3 ;
  RECT 268.777 0.000 269.097 0.600 ;
  LAYER ME2 ;
  RECT 268.777 0.000 269.097 0.600 ;
  LAYER ME1 ;
  RECT 268.777 0.000 269.097 0.600 ;
 END
 ANTENNAPARTIALMETALAREA                  5.273 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME3 ;
 ANTENNADIFFAREA                          1.293 LAYER ME4 ;
END DO57
PIN DI56
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 265.335 0.000 265.655 0.600 ;
  LAYER ME3 ;
  RECT 265.335 0.000 265.655 0.600 ;
  LAYER ME2 ;
  RECT 265.335 0.000 265.655 0.600 ;
  LAYER ME1 ;
  RECT 265.335 0.000 265.655 0.600 ;
 END
 ANTENNAPARTIALMETALAREA                  1.058 LAYER ME2 ;
 ANTENNAGATEAREA                          0.072 LAYER ME2 ;
 ANTENNAGATEAREA                          0.072 LAYER ME3 ;
 ANTENNAGATEAREA                          0.072 LAYER ME4 ;
 ANTENNADIFFAREA                          0.160 LAYER ME2 ;
 ANTENNADIFFAREA                          0.160 LAYER ME3 ;
 ANTENNADIFFAREA                          0.160 LAYER ME4 ;
 ANTENNAMAXAREACAR                       21.782 LAYER ME2 ;
 ANTENNAMAXAREACAR                       24.449 LAYER ME3 ;
 ANTENNAMAXAREACAR                       27.116 LAYER ME4 ;
END DI56
PIN DO56
  DIRECTION OUTPUT ;
 PORT
  LAYER ME4 ;
  RECT 264.773 0.000 265.093 0.600 ;
  LAYER ME3 ;
  RECT 264.773 0.000 265.093 0.600 ;
  LAYER ME2 ;
  RECT 264.773 0.000 265.093 0.600 ;
  LAYER ME1 ;
  RECT 264.773 0.000 265.093 0.600 ;
 END
 ANTENNAPARTIALMETALAREA                  5.273 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME3 ;
 ANTENNADIFFAREA                          1.293 LAYER ME4 ;
END DO56
PIN DI55
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 260.769 0.000 261.089 0.600 ;
  LAYER ME3 ;
  RECT 260.769 0.000 261.089 0.600 ;
  LAYER ME2 ;
  RECT 260.769 0.000 261.089 0.600 ;
  LAYER ME1 ;
  RECT 260.769 0.000 261.089 0.600 ;
 END
 ANTENNAPARTIALMETALAREA                  0.346 LAYER ME1 ;
 ANTENNAPARTIALMETALAREA                  1.466 LAYER ME2 ;
 ANTENNAPARTIALMETALAREA                  0.508 LAYER ME3 ;
 ANTENNAGATEAREA                          0.072 LAYER ME3 ;
 ANTENNAGATEAREA                          0.072 LAYER ME4 ;
 ANTENNADIFFAREA                          0.218 LAYER ME1 ;
 ANTENNADIFFAREA                          0.218 LAYER ME2 ;
 ANTENNADIFFAREA                          0.218 LAYER ME3 ;
 ANTENNADIFFAREA                          0.218 LAYER ME4 ;
 ANTENNAMAXAREACAR                       17.267 LAYER ME3 ;
 ANTENNAMAXAREACAR                       19.933 LAYER ME4 ;
END DI55
PIN DO55
  DIRECTION OUTPUT ;
 PORT
  LAYER ME4 ;
  RECT 261.331 0.000 261.651 0.600 ;
  LAYER ME3 ;
  RECT 261.331 0.000 261.651 0.600 ;
  LAYER ME2 ;
  RECT 261.331 0.000 261.651 0.600 ;
  LAYER ME1 ;
  RECT 261.331 0.000 261.651 0.600 ;
 END
 ANTENNAPARTIALMETALAREA                  5.602 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME3 ;
 ANTENNADIFFAREA                          1.293 LAYER ME4 ;
END DO55
PIN WEB5
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 259.329 0.000 259.649 0.600 ;
  LAYER ME3 ;
  RECT 259.329 0.000 259.649 0.600 ;
  LAYER ME2 ;
  RECT 259.329 0.000 259.649 0.600 ;
  LAYER ME1 ;
  RECT 259.329 0.000 259.649 0.600 ;
 END
 ANTENNAPARTIALMETALAREA                  1.036 LAYER ME2 ;
 ANTENNAGATEAREA                          0.288 LAYER ME2 ;
 ANTENNAGATEAREA                          0.288 LAYER ME3 ;
 ANTENNAGATEAREA                          0.288 LAYER ME4 ;
 ANTENNADIFFAREA                          0.206 LAYER ME2 ;
 ANTENNADIFFAREA                          0.206 LAYER ME3 ;
 ANTENNADIFFAREA                          0.206 LAYER ME4 ;
 ANTENNAMAXAREACAR                        5.844 LAYER ME2 ;
 ANTENNAMAXAREACAR                        6.511 LAYER ME3 ;
 ANTENNAMAXAREACAR                        7.178 LAYER ME4 ;
END WEB5
PIN DI54
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 257.327 0.000 257.647 0.600 ;
  LAYER ME3 ;
  RECT 257.327 0.000 257.647 0.600 ;
  LAYER ME2 ;
  RECT 257.327 0.000 257.647 0.600 ;
  LAYER ME1 ;
  RECT 257.327 0.000 257.647 0.600 ;
 END
 ANTENNAPARTIALMETALAREA                  1.058 LAYER ME2 ;
 ANTENNAGATEAREA                          0.072 LAYER ME2 ;
 ANTENNAGATEAREA                          0.072 LAYER ME3 ;
 ANTENNAGATEAREA                          0.072 LAYER ME4 ;
 ANTENNADIFFAREA                          0.160 LAYER ME2 ;
 ANTENNADIFFAREA                          0.160 LAYER ME3 ;
 ANTENNADIFFAREA                          0.160 LAYER ME4 ;
 ANTENNAMAXAREACAR                       21.782 LAYER ME2 ;
 ANTENNAMAXAREACAR                       24.449 LAYER ME3 ;
 ANTENNAMAXAREACAR                       27.116 LAYER ME4 ;
END DI54
PIN DO54
  DIRECTION OUTPUT ;
 PORT
  LAYER ME4 ;
  RECT 256.765 0.000 257.085 0.600 ;
  LAYER ME3 ;
  RECT 256.765 0.000 257.085 0.600 ;
  LAYER ME2 ;
  RECT 256.765 0.000 257.085 0.600 ;
  LAYER ME1 ;
  RECT 256.765 0.000 257.085 0.600 ;
 END
 ANTENNAPARTIALMETALAREA                  5.273 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME3 ;
 ANTENNADIFFAREA                          1.293 LAYER ME4 ;
END DO54
PIN DI53
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 253.323 0.000 253.643 0.600 ;
  LAYER ME3 ;
  RECT 253.323 0.000 253.643 0.600 ;
  LAYER ME2 ;
  RECT 253.323 0.000 253.643 0.600 ;
  LAYER ME1 ;
  RECT 253.323 0.000 253.643 0.600 ;
 END
 ANTENNAPARTIALMETALAREA                  1.058 LAYER ME2 ;
 ANTENNAGATEAREA                          0.072 LAYER ME2 ;
 ANTENNAGATEAREA                          0.072 LAYER ME3 ;
 ANTENNAGATEAREA                          0.072 LAYER ME4 ;
 ANTENNADIFFAREA                          0.160 LAYER ME2 ;
 ANTENNADIFFAREA                          0.160 LAYER ME3 ;
 ANTENNADIFFAREA                          0.160 LAYER ME4 ;
 ANTENNAMAXAREACAR                       21.782 LAYER ME2 ;
 ANTENNAMAXAREACAR                       24.449 LAYER ME3 ;
 ANTENNAMAXAREACAR                       27.116 LAYER ME4 ;
END DI53
PIN DO53
  DIRECTION OUTPUT ;
 PORT
  LAYER ME4 ;
  RECT 252.761 0.000 253.081 0.600 ;
  LAYER ME3 ;
  RECT 252.761 0.000 253.081 0.600 ;
  LAYER ME2 ;
  RECT 252.761 0.000 253.081 0.600 ;
  LAYER ME1 ;
  RECT 252.761 0.000 253.081 0.600 ;
 END
 ANTENNAPARTIALMETALAREA                  5.273 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME3 ;
 ANTENNADIFFAREA                          1.293 LAYER ME4 ;
END DO53
PIN DI52
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 249.319 0.000 249.639 0.600 ;
  LAYER ME3 ;
  RECT 249.319 0.000 249.639 0.600 ;
  LAYER ME2 ;
  RECT 249.319 0.000 249.639 0.600 ;
  LAYER ME1 ;
  RECT 249.319 0.000 249.639 0.600 ;
 END
 ANTENNAPARTIALMETALAREA                  1.058 LAYER ME2 ;
 ANTENNAGATEAREA                          0.072 LAYER ME2 ;
 ANTENNAGATEAREA                          0.072 LAYER ME3 ;
 ANTENNAGATEAREA                          0.072 LAYER ME4 ;
 ANTENNADIFFAREA                          0.160 LAYER ME2 ;
 ANTENNADIFFAREA                          0.160 LAYER ME3 ;
 ANTENNADIFFAREA                          0.160 LAYER ME4 ;
 ANTENNAMAXAREACAR                       21.782 LAYER ME2 ;
 ANTENNAMAXAREACAR                       24.449 LAYER ME3 ;
 ANTENNAMAXAREACAR                       27.116 LAYER ME4 ;
END DI52
PIN DO52
  DIRECTION OUTPUT ;
 PORT
  LAYER ME4 ;
  RECT 248.757 0.000 249.077 0.600 ;
  LAYER ME3 ;
  RECT 248.757 0.000 249.077 0.600 ;
  LAYER ME2 ;
  RECT 248.757 0.000 249.077 0.600 ;
  LAYER ME1 ;
  RECT 248.757 0.000 249.077 0.600 ;
 END
 ANTENNAPARTIALMETALAREA                  5.273 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME3 ;
 ANTENNADIFFAREA                          1.293 LAYER ME4 ;
END DO52
PIN DI51
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 245.315 0.000 245.635 0.600 ;
  LAYER ME3 ;
  RECT 245.315 0.000 245.635 0.600 ;
  LAYER ME2 ;
  RECT 245.315 0.000 245.635 0.600 ;
  LAYER ME1 ;
  RECT 245.315 0.000 245.635 0.600 ;
 END
 ANTENNAPARTIALMETALAREA                  1.058 LAYER ME2 ;
 ANTENNAGATEAREA                          0.072 LAYER ME2 ;
 ANTENNAGATEAREA                          0.072 LAYER ME3 ;
 ANTENNAGATEAREA                          0.072 LAYER ME4 ;
 ANTENNADIFFAREA                          0.160 LAYER ME2 ;
 ANTENNADIFFAREA                          0.160 LAYER ME3 ;
 ANTENNADIFFAREA                          0.160 LAYER ME4 ;
 ANTENNAMAXAREACAR                       21.782 LAYER ME2 ;
 ANTENNAMAXAREACAR                       24.449 LAYER ME3 ;
 ANTENNAMAXAREACAR                       27.116 LAYER ME4 ;
END DI51
PIN DO51
  DIRECTION OUTPUT ;
 PORT
  LAYER ME4 ;
  RECT 244.753 0.000 245.073 0.600 ;
  LAYER ME3 ;
  RECT 244.753 0.000 245.073 0.600 ;
  LAYER ME2 ;
  RECT 244.753 0.000 245.073 0.600 ;
  LAYER ME1 ;
  RECT 244.753 0.000 245.073 0.600 ;
 END
 ANTENNAPARTIALMETALAREA                  5.273 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME3 ;
 ANTENNADIFFAREA                          1.293 LAYER ME4 ;
END DO51
PIN DI50
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 241.311 0.000 241.631 0.600 ;
  LAYER ME3 ;
  RECT 241.311 0.000 241.631 0.600 ;
  LAYER ME2 ;
  RECT 241.311 0.000 241.631 0.600 ;
  LAYER ME1 ;
  RECT 241.311 0.000 241.631 0.600 ;
 END
 ANTENNAPARTIALMETALAREA                  1.058 LAYER ME2 ;
 ANTENNAGATEAREA                          0.072 LAYER ME2 ;
 ANTENNAGATEAREA                          0.072 LAYER ME3 ;
 ANTENNAGATEAREA                          0.072 LAYER ME4 ;
 ANTENNADIFFAREA                          0.160 LAYER ME2 ;
 ANTENNADIFFAREA                          0.160 LAYER ME3 ;
 ANTENNADIFFAREA                          0.160 LAYER ME4 ;
 ANTENNAMAXAREACAR                       21.782 LAYER ME2 ;
 ANTENNAMAXAREACAR                       24.449 LAYER ME3 ;
 ANTENNAMAXAREACAR                       27.116 LAYER ME4 ;
END DI50
PIN DO50
  DIRECTION OUTPUT ;
 PORT
  LAYER ME4 ;
  RECT 240.749 0.000 241.069 0.600 ;
  LAYER ME3 ;
  RECT 240.749 0.000 241.069 0.600 ;
  LAYER ME2 ;
  RECT 240.749 0.000 241.069 0.600 ;
  LAYER ME1 ;
  RECT 240.749 0.000 241.069 0.600 ;
 END
 ANTENNAPARTIALMETALAREA                  5.273 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME3 ;
 ANTENNADIFFAREA                          1.293 LAYER ME4 ;
END DO50
PIN DI49
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 237.307 0.000 237.627 0.600 ;
  LAYER ME3 ;
  RECT 237.307 0.000 237.627 0.600 ;
  LAYER ME2 ;
  RECT 237.307 0.000 237.627 0.600 ;
  LAYER ME1 ;
  RECT 237.307 0.000 237.627 0.600 ;
 END
 ANTENNAPARTIALMETALAREA                  1.058 LAYER ME2 ;
 ANTENNAGATEAREA                          0.072 LAYER ME2 ;
 ANTENNAGATEAREA                          0.072 LAYER ME3 ;
 ANTENNAGATEAREA                          0.072 LAYER ME4 ;
 ANTENNADIFFAREA                          0.160 LAYER ME2 ;
 ANTENNADIFFAREA                          0.160 LAYER ME3 ;
 ANTENNADIFFAREA                          0.160 LAYER ME4 ;
 ANTENNAMAXAREACAR                       21.782 LAYER ME2 ;
 ANTENNAMAXAREACAR                       24.449 LAYER ME3 ;
 ANTENNAMAXAREACAR                       27.116 LAYER ME4 ;
END DI49
PIN DO49
  DIRECTION OUTPUT ;
 PORT
  LAYER ME4 ;
  RECT 236.745 0.000 237.065 0.600 ;
  LAYER ME3 ;
  RECT 236.745 0.000 237.065 0.600 ;
  LAYER ME2 ;
  RECT 236.745 0.000 237.065 0.600 ;
  LAYER ME1 ;
  RECT 236.745 0.000 237.065 0.600 ;
 END
 ANTENNAPARTIALMETALAREA                  5.273 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME3 ;
 ANTENNADIFFAREA                          1.293 LAYER ME4 ;
END DO49
PIN DI48
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 233.303 0.000 233.623 0.600 ;
  LAYER ME3 ;
  RECT 233.303 0.000 233.623 0.600 ;
  LAYER ME2 ;
  RECT 233.303 0.000 233.623 0.600 ;
  LAYER ME1 ;
  RECT 233.303 0.000 233.623 0.600 ;
 END
 ANTENNAPARTIALMETALAREA                  1.058 LAYER ME2 ;
 ANTENNAGATEAREA                          0.072 LAYER ME2 ;
 ANTENNAGATEAREA                          0.072 LAYER ME3 ;
 ANTENNAGATEAREA                          0.072 LAYER ME4 ;
 ANTENNADIFFAREA                          0.160 LAYER ME2 ;
 ANTENNADIFFAREA                          0.160 LAYER ME3 ;
 ANTENNADIFFAREA                          0.160 LAYER ME4 ;
 ANTENNAMAXAREACAR                       21.782 LAYER ME2 ;
 ANTENNAMAXAREACAR                       24.449 LAYER ME3 ;
 ANTENNAMAXAREACAR                       27.116 LAYER ME4 ;
END DI48
PIN DO48
  DIRECTION OUTPUT ;
 PORT
  LAYER ME4 ;
  RECT 232.741 0.000 233.061 0.600 ;
  LAYER ME3 ;
  RECT 232.741 0.000 233.061 0.600 ;
  LAYER ME2 ;
  RECT 232.741 0.000 233.061 0.600 ;
  LAYER ME1 ;
  RECT 232.741 0.000 233.061 0.600 ;
 END
 ANTENNAPARTIALMETALAREA                  5.273 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME3 ;
 ANTENNADIFFAREA                          1.293 LAYER ME4 ;
END DO48
PIN DI47
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 229.299 0.000 229.619 0.600 ;
  LAYER ME3 ;
  RECT 229.299 0.000 229.619 0.600 ;
  LAYER ME2 ;
  RECT 229.299 0.000 229.619 0.600 ;
  LAYER ME1 ;
  RECT 229.299 0.000 229.619 0.600 ;
 END
 ANTENNAPARTIALMETALAREA                  1.058 LAYER ME2 ;
 ANTENNAGATEAREA                          0.072 LAYER ME2 ;
 ANTENNAGATEAREA                          0.072 LAYER ME3 ;
 ANTENNAGATEAREA                          0.072 LAYER ME4 ;
 ANTENNADIFFAREA                          0.160 LAYER ME2 ;
 ANTENNADIFFAREA                          0.160 LAYER ME3 ;
 ANTENNADIFFAREA                          0.160 LAYER ME4 ;
 ANTENNAMAXAREACAR                       21.782 LAYER ME2 ;
 ANTENNAMAXAREACAR                       24.449 LAYER ME3 ;
 ANTENNAMAXAREACAR                       27.116 LAYER ME4 ;
END DI47
PIN DO47
  DIRECTION OUTPUT ;
 PORT
  LAYER ME4 ;
  RECT 228.737 0.000 229.057 0.600 ;
  LAYER ME3 ;
  RECT 228.737 0.000 229.057 0.600 ;
  LAYER ME2 ;
  RECT 228.737 0.000 229.057 0.600 ;
  LAYER ME1 ;
  RECT 228.737 0.000 229.057 0.600 ;
 END
 ANTENNAPARTIALMETALAREA                  5.273 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME3 ;
 ANTENNADIFFAREA                          1.293 LAYER ME4 ;
END DO47
PIN DI46
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 225.295 0.000 225.615 0.600 ;
  LAYER ME3 ;
  RECT 225.295 0.000 225.615 0.600 ;
  LAYER ME2 ;
  RECT 225.295 0.000 225.615 0.600 ;
  LAYER ME1 ;
  RECT 225.295 0.000 225.615 0.600 ;
 END
 ANTENNAPARTIALMETALAREA                  1.058 LAYER ME2 ;
 ANTENNAGATEAREA                          0.072 LAYER ME2 ;
 ANTENNAGATEAREA                          0.072 LAYER ME3 ;
 ANTENNAGATEAREA                          0.072 LAYER ME4 ;
 ANTENNADIFFAREA                          0.160 LAYER ME2 ;
 ANTENNADIFFAREA                          0.160 LAYER ME3 ;
 ANTENNADIFFAREA                          0.160 LAYER ME4 ;
 ANTENNAMAXAREACAR                       21.782 LAYER ME2 ;
 ANTENNAMAXAREACAR                       24.449 LAYER ME3 ;
 ANTENNAMAXAREACAR                       27.116 LAYER ME4 ;
END DI46
PIN DO46
  DIRECTION OUTPUT ;
 PORT
  LAYER ME4 ;
  RECT 224.733 0.000 225.053 0.600 ;
  LAYER ME3 ;
  RECT 224.733 0.000 225.053 0.600 ;
  LAYER ME2 ;
  RECT 224.733 0.000 225.053 0.600 ;
  LAYER ME1 ;
  RECT 224.733 0.000 225.053 0.600 ;
 END
 ANTENNAPARTIALMETALAREA                  5.273 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME3 ;
 ANTENNADIFFAREA                          1.293 LAYER ME4 ;
END DO46
PIN DI45
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 221.291 0.000 221.611 0.600 ;
  LAYER ME3 ;
  RECT 221.291 0.000 221.611 0.600 ;
  LAYER ME2 ;
  RECT 221.291 0.000 221.611 0.600 ;
  LAYER ME1 ;
  RECT 221.291 0.000 221.611 0.600 ;
 END
 ANTENNAPARTIALMETALAREA                  1.058 LAYER ME2 ;
 ANTENNAGATEAREA                          0.072 LAYER ME2 ;
 ANTENNAGATEAREA                          0.072 LAYER ME3 ;
 ANTENNAGATEAREA                          0.072 LAYER ME4 ;
 ANTENNADIFFAREA                          0.160 LAYER ME2 ;
 ANTENNADIFFAREA                          0.160 LAYER ME3 ;
 ANTENNADIFFAREA                          0.160 LAYER ME4 ;
 ANTENNAMAXAREACAR                       21.782 LAYER ME2 ;
 ANTENNAMAXAREACAR                       24.449 LAYER ME3 ;
 ANTENNAMAXAREACAR                       27.116 LAYER ME4 ;
END DI45
PIN DO45
  DIRECTION OUTPUT ;
 PORT
  LAYER ME4 ;
  RECT 220.729 0.000 221.049 0.600 ;
  LAYER ME3 ;
  RECT 220.729 0.000 221.049 0.600 ;
  LAYER ME2 ;
  RECT 220.729 0.000 221.049 0.600 ;
  LAYER ME1 ;
  RECT 220.729 0.000 221.049 0.600 ;
 END
 ANTENNAPARTIALMETALAREA                  5.273 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME3 ;
 ANTENNADIFFAREA                          1.293 LAYER ME4 ;
END DO45
PIN DI44
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 216.725 0.000 217.045 0.600 ;
  LAYER ME3 ;
  RECT 216.725 0.000 217.045 0.600 ;
  LAYER ME2 ;
  RECT 216.725 0.000 217.045 0.600 ;
  LAYER ME1 ;
  RECT 216.725 0.000 217.045 0.600 ;
 END
 ANTENNAPARTIALMETALAREA                  0.346 LAYER ME1 ;
 ANTENNAPARTIALMETALAREA                  1.466 LAYER ME2 ;
 ANTENNAPARTIALMETALAREA                  0.508 LAYER ME3 ;
 ANTENNAGATEAREA                          0.072 LAYER ME3 ;
 ANTENNAGATEAREA                          0.072 LAYER ME4 ;
 ANTENNADIFFAREA                          0.218 LAYER ME1 ;
 ANTENNADIFFAREA                          0.218 LAYER ME2 ;
 ANTENNADIFFAREA                          0.218 LAYER ME3 ;
 ANTENNADIFFAREA                          0.218 LAYER ME4 ;
 ANTENNAMAXAREACAR                       17.267 LAYER ME3 ;
 ANTENNAMAXAREACAR                       19.933 LAYER ME4 ;
END DI44
PIN DO44
  DIRECTION OUTPUT ;
 PORT
  LAYER ME4 ;
  RECT 217.287 0.000 217.607 0.600 ;
  LAYER ME3 ;
  RECT 217.287 0.000 217.607 0.600 ;
  LAYER ME2 ;
  RECT 217.287 0.000 217.607 0.600 ;
  LAYER ME1 ;
  RECT 217.287 0.000 217.607 0.600 ;
 END
 ANTENNAPARTIALMETALAREA                  5.602 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME3 ;
 ANTENNADIFFAREA                          1.293 LAYER ME4 ;
END DO44
PIN WEB4
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 215.285 0.000 215.605 0.600 ;
  LAYER ME3 ;
  RECT 215.285 0.000 215.605 0.600 ;
  LAYER ME2 ;
  RECT 215.285 0.000 215.605 0.600 ;
  LAYER ME1 ;
  RECT 215.285 0.000 215.605 0.600 ;
 END
 ANTENNAPARTIALMETALAREA                  1.036 LAYER ME2 ;
 ANTENNAGATEAREA                          0.288 LAYER ME2 ;
 ANTENNAGATEAREA                          0.288 LAYER ME3 ;
 ANTENNAGATEAREA                          0.288 LAYER ME4 ;
 ANTENNADIFFAREA                          0.206 LAYER ME2 ;
 ANTENNADIFFAREA                          0.206 LAYER ME3 ;
 ANTENNADIFFAREA                          0.206 LAYER ME4 ;
 ANTENNAMAXAREACAR                        5.844 LAYER ME2 ;
 ANTENNAMAXAREACAR                        6.511 LAYER ME3 ;
 ANTENNAMAXAREACAR                        7.178 LAYER ME4 ;
END WEB4
OBS
  LAYER ME3 SPACING 0.260 ;
  RECT 0.000 0.000 394.251 66.831 ;
  LAYER ME2 SPACING 0.260 ;
  RECT 0.000 0.000 394.251 66.831 ;
  LAYER ME1 SPACING 0.260 ;
  RECT 0.000 0.000 394.251 66.831 ;
  LAYER ME4 SPACING 0.260 ;
  RECT 0.000 0.000 190.318 66.831 ;
  LAYER ME4 SPACING 0.260 ;
  RECT 191.972 0.000 193.092 66.831 ;
  LAYER ME4 SPACING 0.260 ;
  RECT 194.687 0.000 195.407 66.831 ;
  LAYER ME4 SPACING 0.260 ;
  RECT 196.137 0.000 196.857 66.831 ;
  LAYER ME4 SPACING 0.260 ;
  RECT 198.917 0.000 199.517 66.831 ;
  LAYER ME4 SPACING 0.260 ;
  RECT 202.131 0.000 203.817 66.831 ;
  LAYER ME4 SPACING 0.260 ;
  RECT 205.207 0.000 206.327 66.831 ;
  LAYER ME4 SPACING 0.260 ;
  RECT 207.602 0.000 208.322 66.831 ;
  LAYER ME4 SPACING 0.260 ;
  RECT 209.317 0.000 210.037 66.831 ;
  LAYER ME4 SPACING 0.260 ;
  RECT 211.237 0.000 394.251 66.831 ;
END
END SYKB110_32X11X8CM2
END LIBRARY





