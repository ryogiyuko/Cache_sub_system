# ________________________________________________________________________________________________
# 
# 
#             Synchronous One-Port Register File Compiler
# 
#                 UMC 0.11um LL AE Logic Process
# 
# ________________________________________________________________________________________________
# 
#               
#         Copyright (C) 2024 Faraday Technology Corporation. All Rights Reserved.       
#                
#         This source code is an unpublished work belongs to Faraday Technology Corporation       
#         It is considered a trade secret and is not to be divulged or       
#         used by parties who have not received written authorization from       
#         Faraday Technology Corporation       
#                
#         Faraday's home page can be found at: http://www.faraday-tech.com/       
#                
# ________________________________________________________________________________________________
# 
#        IP Name            :  FSR0K_B_SY                
#        IP Version         :  1.4.0                     
#        IP Release Status  :  Active                    
#        Word               :  1024                      
#        Bit                :  8                         
#        Byte               :  8                         
#        Mux                :  4                         
#        Output Loading     :  0.01                      
#        Clock Input Slew   :  0.016                     
#        Data Input Slew    :  0.016                     
#        Ring Type          :  Ringless Model            
#        Ring Width         :  0                         
#        Bus Format         :  0                         
#        Memaker Path       :  /home/mem/Desktop/memlib  
#        GUI Version        :  m20230904                 
#        Date               :  2024/10/18 14:57:08       
# ________________________________________________________________________________________________
# 

VERSION 5.5 ;
NAMESCASESENSITIVE ON ;
MACRO SYKB110_1024X8X8CM4
CLASS BLOCK ;
FOREIGN SYKB110_1024X8X8CM4 0.000 0.000 ;
ORIGIN 0.000 0.000 ;
SIZE 557.611 BY 280.651 ;
SYMMETRY x y r90 ;
SITE core ;
PIN VCC
  DIRECTION INOUT ;
  USE POWER ;
 PORT
  LAYER ME4 ;
  RECT 303.089 0.000 303.809 33.870 ;
 END
 PORT
  LAYER ME4 ;
  RECT 299.085 0.000 299.805 33.870 ;
 END
 PORT
  LAYER ME4 ;
  RECT 311.097 0.000 311.817 33.870 ;
 END
 PORT
  LAYER ME4 ;
  RECT 307.093 0.000 307.813 33.870 ;
 END
 PORT
  LAYER ME4 ;
  RECT 319.105 0.000 319.825 33.870 ;
 END
 PORT
  LAYER ME4 ;
  RECT 315.101 0.000 315.821 33.870 ;
 END
 PORT
  LAYER ME4 ;
  RECT 327.113 0.000 327.833 33.870 ;
 END
 PORT
  LAYER ME4 ;
  RECT 323.109 0.000 323.829 33.870 ;
 END
 PORT
  LAYER ME4 ;
  RECT 335.121 0.000 335.841 33.870 ;
 END
 PORT
  LAYER ME4 ;
  RECT 331.117 0.000 331.837 33.870 ;
 END
 PORT
  LAYER ME4 ;
  RECT 343.129 0.000 343.849 33.870 ;
 END
 PORT
  LAYER ME4 ;
  RECT 339.125 0.000 339.845 33.870 ;
 END
 PORT
  LAYER ME4 ;
  RECT 351.137 0.000 351.857 33.870 ;
 END
 PORT
  LAYER ME4 ;
  RECT 347.133 0.000 347.853 33.870 ;
 END
 PORT
  LAYER ME4 ;
  RECT 359.145 0.000 359.865 33.870 ;
 END
 PORT
  LAYER ME4 ;
  RECT 355.141 0.000 355.861 33.870 ;
 END
 PORT
  LAYER ME4 ;
  RECT 367.153 0.000 367.873 33.870 ;
 END
 PORT
  LAYER ME4 ;
  RECT 363.149 0.000 363.869 33.870 ;
 END
 PORT
  LAYER ME4 ;
  RECT 375.161 0.000 375.881 33.870 ;
 END
 PORT
  LAYER ME4 ;
  RECT 371.157 0.000 371.877 33.870 ;
 END
 PORT
  LAYER ME4 ;
  RECT 383.169 0.000 383.889 33.870 ;
 END
 PORT
  LAYER ME4 ;
  RECT 379.165 0.000 379.885 33.870 ;
 END
 PORT
  LAYER ME4 ;
  RECT 391.177 0.000 391.897 33.870 ;
 END
 PORT
  LAYER ME4 ;
  RECT 387.173 0.000 387.893 33.870 ;
 END
 PORT
  LAYER ME4 ;
  RECT 399.185 0.000 399.905 33.870 ;
 END
 PORT
  LAYER ME4 ;
  RECT 395.181 0.000 395.901 33.870 ;
 END
 PORT
  LAYER ME4 ;
  RECT 407.193 0.000 407.913 33.870 ;
 END
 PORT
  LAYER ME4 ;
  RECT 403.189 0.000 403.909 33.870 ;
 END
 PORT
  LAYER ME4 ;
  RECT 415.201 0.000 415.921 33.870 ;
 END
 PORT
  LAYER ME4 ;
  RECT 411.197 0.000 411.917 33.870 ;
 END
 PORT
  LAYER ME4 ;
  RECT 423.209 0.000 423.929 33.870 ;
 END
 PORT
  LAYER ME4 ;
  RECT 419.205 0.000 419.925 33.870 ;
 END
 PORT
  LAYER ME4 ;
  RECT 431.217 0.000 431.937 33.870 ;
 END
 PORT
  LAYER ME4 ;
  RECT 427.213 0.000 427.933 33.870 ;
 END
 PORT
  LAYER ME4 ;
  RECT 439.225 0.000 439.945 33.870 ;
 END
 PORT
  LAYER ME4 ;
  RECT 435.221 0.000 435.941 33.870 ;
 END
 PORT
  LAYER ME4 ;
  RECT 447.233 0.000 447.953 33.870 ;
 END
 PORT
  LAYER ME4 ;
  RECT 443.229 0.000 443.949 33.870 ;
 END
 PORT
  LAYER ME4 ;
  RECT 455.241 0.000 455.961 33.870 ;
 END
 PORT
  LAYER ME4 ;
  RECT 451.237 0.000 451.957 33.870 ;
 END
 PORT
  LAYER ME4 ;
  RECT 463.249 0.000 463.969 33.870 ;
 END
 PORT
  LAYER ME4 ;
  RECT 459.245 0.000 459.965 33.870 ;
 END
 PORT
  LAYER ME4 ;
  RECT 471.257 0.000 471.977 33.870 ;
 END
 PORT
  LAYER ME4 ;
  RECT 467.253 0.000 467.973 33.870 ;
 END
 PORT
  LAYER ME4 ;
  RECT 479.265 0.000 479.985 33.870 ;
 END
 PORT
  LAYER ME4 ;
  RECT 475.261 0.000 475.981 33.870 ;
 END
 PORT
  LAYER ME4 ;
  RECT 487.273 0.000 487.993 33.870 ;
 END
 PORT
  LAYER ME4 ;
  RECT 483.269 0.000 483.989 33.870 ;
 END
 PORT
  LAYER ME4 ;
  RECT 495.281 0.000 496.001 33.870 ;
 END
 PORT
  LAYER ME4 ;
  RECT 491.277 0.000 491.997 33.870 ;
 END
 PORT
  LAYER ME4 ;
  RECT 503.289 0.000 504.009 33.870 ;
 END
 PORT
  LAYER ME4 ;
  RECT 499.285 0.000 500.005 33.870 ;
 END
 PORT
  LAYER ME4 ;
  RECT 511.297 0.000 512.017 33.870 ;
 END
 PORT
  LAYER ME4 ;
  RECT 507.293 0.000 508.013 33.870 ;
 END
 PORT
  LAYER ME4 ;
  RECT 519.305 0.000 520.025 33.870 ;
 END
 PORT
  LAYER ME4 ;
  RECT 515.301 0.000 516.021 33.870 ;
 END
 PORT
  LAYER ME4 ;
  RECT 527.313 0.000 528.033 33.870 ;
 END
 PORT
  LAYER ME4 ;
  RECT 523.309 0.000 524.029 33.870 ;
 END
 PORT
  LAYER ME4 ;
  RECT 535.321 0.000 536.041 33.870 ;
 END
 PORT
  LAYER ME4 ;
  RECT 531.317 0.000 532.037 33.870 ;
 END
 PORT
  LAYER ME4 ;
  RECT 543.329 0.000 544.049 33.870 ;
 END
 PORT
  LAYER ME4 ;
  RECT 539.325 0.000 540.045 33.870 ;
 END
 PORT
  LAYER ME4 ;
  RECT 551.337 0.000 552.057 33.870 ;
 END
 PORT
  LAYER ME4 ;
  RECT 547.333 0.000 548.053 33.870 ;
 END
 PORT
  LAYER ME4 ;
  RECT 556.311 0.000 556.691 280.651 ;
 END
 PORT
  LAYER ME4 ;
  RECT 282.197 0.000 282.797 280.651 ;
 END
 PORT
  LAYER ME4 ;
  RECT 286.377 0.000 287.097 280.651 ;
 END
 PORT
  LAYER ME4 ;
  RECT 288.487 0.000 289.607 280.651 ;
 END
 PORT
  LAYER ME4 ;
  RECT 294.517 0.000 295.237 280.651 ;
 END
 PORT
  LAYER ME4 ;
  RECT 296.453 0.921 296.833 280.651 ;
 END
 PORT
  LAYER ME4 ;
  RECT 275.252 0.000 276.372 280.651 ;
 END
 PORT
  LAYER ME4 ;
  RECT 277.967 0.000 278.687 280.651 ;
 END
 PORT
  LAYER ME4 ;
  RECT 272.878 0.000 273.598 279.771 ;
 END
 PORT
  LAYER ME4 ;
  RECT 270.838 0.921 271.558 280.651 ;
 END
 PORT
  LAYER ME4 ;
  RECT 268.718 0.000 269.438 280.651 ;
 END
 PORT
  LAYER ME4 ;
  RECT 266.678 0.921 267.398 280.651 ;
 END
 PORT
  LAYER ME4 ;
  RECT 264.558 0.000 265.278 280.651 ;
 END
 PORT
  LAYER ME4 ;
  RECT 262.518 0.921 263.238 280.651 ;
 END
 PORT
  LAYER ME4 ;
  RECT 0.920 0.000 1.300 280.651 ;
 END
 PORT
  LAYER ME4 ;
  RECT 7.556 0.000 8.276 33.870 ;
 END
 PORT
  LAYER ME4 ;
  RECT 3.552 0.000 4.272 33.870 ;
 END
 PORT
  LAYER ME4 ;
  RECT 15.564 0.000 16.284 33.870 ;
 END
 PORT
  LAYER ME4 ;
  RECT 11.560 0.000 12.280 33.870 ;
 END
 PORT
  LAYER ME4 ;
  RECT 23.572 0.000 24.292 33.870 ;
 END
 PORT
  LAYER ME4 ;
  RECT 19.568 0.000 20.288 33.870 ;
 END
 PORT
  LAYER ME4 ;
  RECT 31.580 0.000 32.300 33.870 ;
 END
 PORT
  LAYER ME4 ;
  RECT 27.576 0.000 28.296 33.870 ;
 END
 PORT
  LAYER ME4 ;
  RECT 39.588 0.000 40.308 33.870 ;
 END
 PORT
  LAYER ME4 ;
  RECT 35.584 0.000 36.304 33.870 ;
 END
 PORT
  LAYER ME4 ;
  RECT 47.596 0.000 48.316 33.870 ;
 END
 PORT
  LAYER ME4 ;
  RECT 43.592 0.000 44.312 33.870 ;
 END
 PORT
  LAYER ME4 ;
  RECT 55.604 0.000 56.324 33.870 ;
 END
 PORT
  LAYER ME4 ;
  RECT 51.600 0.000 52.320 33.870 ;
 END
 PORT
  LAYER ME4 ;
  RECT 63.612 0.000 64.332 33.870 ;
 END
 PORT
  LAYER ME4 ;
  RECT 59.608 0.000 60.328 33.870 ;
 END
 PORT
  LAYER ME4 ;
  RECT 71.620 0.000 72.340 33.870 ;
 END
 PORT
  LAYER ME4 ;
  RECT 67.616 0.000 68.336 33.870 ;
 END
 PORT
  LAYER ME4 ;
  RECT 79.628 0.000 80.348 33.870 ;
 END
 PORT
  LAYER ME4 ;
  RECT 75.624 0.000 76.344 33.870 ;
 END
 PORT
  LAYER ME4 ;
  RECT 87.636 0.000 88.356 33.870 ;
 END
 PORT
  LAYER ME4 ;
  RECT 83.632 0.000 84.352 33.870 ;
 END
 PORT
  LAYER ME4 ;
  RECT 95.644 0.000 96.364 33.870 ;
 END
 PORT
  LAYER ME4 ;
  RECT 91.640 0.000 92.360 33.870 ;
 END
 PORT
  LAYER ME4 ;
  RECT 103.652 0.000 104.372 33.870 ;
 END
 PORT
  LAYER ME4 ;
  RECT 99.648 0.000 100.368 33.870 ;
 END
 PORT
  LAYER ME4 ;
  RECT 111.660 0.000 112.380 33.870 ;
 END
 PORT
  LAYER ME4 ;
  RECT 107.656 0.000 108.376 33.870 ;
 END
 PORT
  LAYER ME4 ;
  RECT 119.668 0.000 120.388 33.870 ;
 END
 PORT
  LAYER ME4 ;
  RECT 115.664 0.000 116.384 33.870 ;
 END
 PORT
  LAYER ME4 ;
  RECT 127.676 0.000 128.396 33.870 ;
 END
 PORT
  LAYER ME4 ;
  RECT 123.672 0.000 124.392 33.870 ;
 END
 PORT
  LAYER ME4 ;
  RECT 135.684 0.000 136.404 33.870 ;
 END
 PORT
  LAYER ME4 ;
  RECT 131.680 0.000 132.400 33.870 ;
 END
 PORT
  LAYER ME4 ;
  RECT 143.692 0.000 144.412 33.870 ;
 END
 PORT
  LAYER ME4 ;
  RECT 139.688 0.000 140.408 33.870 ;
 END
 PORT
  LAYER ME4 ;
  RECT 151.700 0.000 152.420 33.870 ;
 END
 PORT
  LAYER ME4 ;
  RECT 147.696 0.000 148.416 33.870 ;
 END
 PORT
  LAYER ME4 ;
  RECT 159.708 0.000 160.428 33.870 ;
 END
 PORT
  LAYER ME4 ;
  RECT 155.704 0.000 156.424 33.870 ;
 END
 PORT
  LAYER ME4 ;
  RECT 167.716 0.000 168.436 33.870 ;
 END
 PORT
  LAYER ME4 ;
  RECT 163.712 0.000 164.432 33.870 ;
 END
 PORT
  LAYER ME4 ;
  RECT 175.724 0.000 176.444 33.870 ;
 END
 PORT
  LAYER ME4 ;
  RECT 171.720 0.000 172.440 33.870 ;
 END
 PORT
  LAYER ME4 ;
  RECT 183.732 0.000 184.452 33.870 ;
 END
 PORT
  LAYER ME4 ;
  RECT 179.728 0.000 180.448 33.870 ;
 END
 PORT
  LAYER ME4 ;
  RECT 191.740 0.000 192.460 33.870 ;
 END
 PORT
  LAYER ME4 ;
  RECT 187.736 0.000 188.456 33.870 ;
 END
 PORT
  LAYER ME4 ;
  RECT 199.748 0.000 200.468 33.870 ;
 END
 PORT
  LAYER ME4 ;
  RECT 195.744 0.000 196.464 33.870 ;
 END
 PORT
  LAYER ME4 ;
  RECT 207.756 0.000 208.476 33.870 ;
 END
 PORT
  LAYER ME4 ;
  RECT 203.752 0.000 204.472 33.870 ;
 END
 PORT
  LAYER ME4 ;
  RECT 215.764 0.000 216.484 33.870 ;
 END
 PORT
  LAYER ME4 ;
  RECT 211.760 0.000 212.480 33.870 ;
 END
 PORT
  LAYER ME4 ;
  RECT 223.772 0.000 224.492 33.870 ;
 END
 PORT
  LAYER ME4 ;
  RECT 219.768 0.000 220.488 33.870 ;
 END
 PORT
  LAYER ME4 ;
  RECT 231.780 0.000 232.500 33.870 ;
 END
 PORT
  LAYER ME4 ;
  RECT 227.776 0.000 228.496 33.870 ;
 END
 PORT
  LAYER ME4 ;
  RECT 239.788 0.000 240.508 33.870 ;
 END
 PORT
  LAYER ME4 ;
  RECT 235.784 0.000 236.504 33.870 ;
 END
 PORT
  LAYER ME4 ;
  RECT 247.796 0.000 248.516 33.870 ;
 END
 PORT
  LAYER ME4 ;
  RECT 243.792 0.000 244.512 33.870 ;
 END
 PORT
  LAYER ME4 ;
  RECT 255.804 0.000 256.524 33.870 ;
 END
 PORT
  LAYER ME4 ;
  RECT 251.800 0.000 252.520 33.870 ;
 END
 PORT
  LAYER ME4 ;
  RECT 260.778 0.000 261.158 280.651 ;
 END
 PORT
  LAYER ME4 ;
  RECT 305.281 35.220 305.621 280.651 ;
 END
 PORT
  LAYER ME4 ;
  RECT 303.279 35.220 303.619 280.651 ;
 END
 PORT
  LAYER ME4 ;
  RECT 301.277 35.220 301.617 280.651 ;
 END
 PORT
  LAYER ME4 ;
  RECT 299.275 35.220 299.615 280.651 ;
 END
 PORT
  LAYER ME4 ;
  RECT 313.289 35.220 313.629 280.651 ;
 END
 PORT
  LAYER ME4 ;
  RECT 311.287 35.220 311.627 280.651 ;
 END
 PORT
  LAYER ME4 ;
  RECT 309.285 35.220 309.625 280.651 ;
 END
 PORT
  LAYER ME4 ;
  RECT 307.283 35.220 307.623 280.651 ;
 END
 PORT
  LAYER ME4 ;
  RECT 321.297 35.220 321.637 280.651 ;
 END
 PORT
  LAYER ME4 ;
  RECT 319.295 35.220 319.635 280.651 ;
 END
 PORT
  LAYER ME4 ;
  RECT 317.293 35.220 317.633 280.651 ;
 END
 PORT
  LAYER ME4 ;
  RECT 315.291 35.220 315.631 280.651 ;
 END
 PORT
  LAYER ME4 ;
  RECT 329.305 35.220 329.645 280.651 ;
 END
 PORT
  LAYER ME4 ;
  RECT 327.303 35.220 327.643 280.651 ;
 END
 PORT
  LAYER ME4 ;
  RECT 325.301 35.220 325.641 280.651 ;
 END
 PORT
  LAYER ME4 ;
  RECT 323.299 35.220 323.639 280.651 ;
 END
 PORT
  LAYER ME4 ;
  RECT 337.313 35.220 337.653 280.651 ;
 END
 PORT
  LAYER ME4 ;
  RECT 335.311 35.220 335.651 280.651 ;
 END
 PORT
  LAYER ME4 ;
  RECT 333.309 35.220 333.649 280.651 ;
 END
 PORT
  LAYER ME4 ;
  RECT 331.307 35.220 331.647 280.651 ;
 END
 PORT
  LAYER ME4 ;
  RECT 345.321 35.220 345.661 280.651 ;
 END
 PORT
  LAYER ME4 ;
  RECT 343.319 35.220 343.659 280.651 ;
 END
 PORT
  LAYER ME4 ;
  RECT 341.317 35.220 341.657 280.651 ;
 END
 PORT
  LAYER ME4 ;
  RECT 339.315 35.220 339.655 280.651 ;
 END
 PORT
  LAYER ME4 ;
  RECT 353.329 35.220 353.669 280.651 ;
 END
 PORT
  LAYER ME4 ;
  RECT 351.327 35.220 351.667 280.651 ;
 END
 PORT
  LAYER ME4 ;
  RECT 349.325 35.220 349.665 280.651 ;
 END
 PORT
  LAYER ME4 ;
  RECT 347.323 35.220 347.663 280.651 ;
 END
 PORT
  LAYER ME4 ;
  RECT 361.337 35.220 361.677 280.651 ;
 END
 PORT
  LAYER ME4 ;
  RECT 359.335 35.220 359.675 280.651 ;
 END
 PORT
  LAYER ME4 ;
  RECT 357.333 35.220 357.673 280.651 ;
 END
 PORT
  LAYER ME4 ;
  RECT 355.331 35.220 355.671 280.651 ;
 END
 PORT
  LAYER ME4 ;
  RECT 369.345 35.220 369.685 280.651 ;
 END
 PORT
  LAYER ME4 ;
  RECT 367.343 35.220 367.683 280.651 ;
 END
 PORT
  LAYER ME4 ;
  RECT 365.341 35.220 365.681 280.651 ;
 END
 PORT
  LAYER ME4 ;
  RECT 363.339 35.220 363.679 280.651 ;
 END
 PORT
  LAYER ME4 ;
  RECT 377.353 35.220 377.693 280.651 ;
 END
 PORT
  LAYER ME4 ;
  RECT 375.351 35.220 375.691 280.651 ;
 END
 PORT
  LAYER ME4 ;
  RECT 373.349 35.220 373.689 280.651 ;
 END
 PORT
  LAYER ME4 ;
  RECT 371.347 35.220 371.687 280.651 ;
 END
 PORT
  LAYER ME4 ;
  RECT 385.361 35.220 385.701 280.651 ;
 END
 PORT
  LAYER ME4 ;
  RECT 383.359 35.220 383.699 280.651 ;
 END
 PORT
  LAYER ME4 ;
  RECT 381.357 35.220 381.697 280.651 ;
 END
 PORT
  LAYER ME4 ;
  RECT 379.355 35.220 379.695 280.651 ;
 END
 PORT
  LAYER ME4 ;
  RECT 393.369 35.220 393.709 280.651 ;
 END
 PORT
  LAYER ME4 ;
  RECT 391.367 35.220 391.707 280.651 ;
 END
 PORT
  LAYER ME4 ;
  RECT 389.365 35.220 389.705 280.651 ;
 END
 PORT
  LAYER ME4 ;
  RECT 387.363 35.220 387.703 280.651 ;
 END
 PORT
  LAYER ME4 ;
  RECT 401.377 35.220 401.717 280.651 ;
 END
 PORT
  LAYER ME4 ;
  RECT 399.375 35.220 399.715 280.651 ;
 END
 PORT
  LAYER ME4 ;
  RECT 397.373 35.220 397.713 280.651 ;
 END
 PORT
  LAYER ME4 ;
  RECT 395.371 35.220 395.711 280.651 ;
 END
 PORT
  LAYER ME4 ;
  RECT 409.385 35.220 409.725 280.651 ;
 END
 PORT
  LAYER ME4 ;
  RECT 407.383 35.220 407.723 280.651 ;
 END
 PORT
  LAYER ME4 ;
  RECT 405.381 35.220 405.721 280.651 ;
 END
 PORT
  LAYER ME4 ;
  RECT 403.379 35.220 403.719 280.651 ;
 END
 PORT
  LAYER ME4 ;
  RECT 417.393 35.220 417.733 280.651 ;
 END
 PORT
  LAYER ME4 ;
  RECT 415.391 35.220 415.731 280.651 ;
 END
 PORT
  LAYER ME4 ;
  RECT 413.389 35.220 413.729 280.651 ;
 END
 PORT
  LAYER ME4 ;
  RECT 411.387 35.220 411.727 280.651 ;
 END
 PORT
  LAYER ME4 ;
  RECT 425.401 35.220 425.741 280.651 ;
 END
 PORT
  LAYER ME4 ;
  RECT 423.399 35.220 423.739 280.651 ;
 END
 PORT
  LAYER ME4 ;
  RECT 421.397 35.220 421.737 280.651 ;
 END
 PORT
  LAYER ME4 ;
  RECT 419.395 35.220 419.735 280.651 ;
 END
 PORT
  LAYER ME4 ;
  RECT 433.409 35.220 433.749 280.651 ;
 END
 PORT
  LAYER ME4 ;
  RECT 431.407 35.220 431.747 280.651 ;
 END
 PORT
  LAYER ME4 ;
  RECT 429.405 35.220 429.745 280.651 ;
 END
 PORT
  LAYER ME4 ;
  RECT 427.403 35.220 427.743 280.651 ;
 END
 PORT
  LAYER ME4 ;
  RECT 441.417 35.220 441.757 280.651 ;
 END
 PORT
  LAYER ME4 ;
  RECT 439.415 35.220 439.755 280.651 ;
 END
 PORT
  LAYER ME4 ;
  RECT 437.413 35.220 437.753 280.651 ;
 END
 PORT
  LAYER ME4 ;
  RECT 435.411 35.220 435.751 280.651 ;
 END
 PORT
  LAYER ME4 ;
  RECT 449.425 35.220 449.765 280.651 ;
 END
 PORT
  LAYER ME4 ;
  RECT 447.423 35.220 447.763 280.651 ;
 END
 PORT
  LAYER ME4 ;
  RECT 445.421 35.220 445.761 280.651 ;
 END
 PORT
  LAYER ME4 ;
  RECT 443.419 35.220 443.759 280.651 ;
 END
 PORT
  LAYER ME4 ;
  RECT 457.433 35.220 457.773 280.651 ;
 END
 PORT
  LAYER ME4 ;
  RECT 455.431 35.220 455.771 280.651 ;
 END
 PORT
  LAYER ME4 ;
  RECT 453.429 35.220 453.769 280.651 ;
 END
 PORT
  LAYER ME4 ;
  RECT 451.427 35.220 451.767 280.651 ;
 END
 PORT
  LAYER ME4 ;
  RECT 465.441 35.220 465.781 280.651 ;
 END
 PORT
  LAYER ME4 ;
  RECT 463.439 35.220 463.779 280.651 ;
 END
 PORT
  LAYER ME4 ;
  RECT 461.437 35.220 461.777 280.651 ;
 END
 PORT
  LAYER ME4 ;
  RECT 459.435 35.220 459.775 280.651 ;
 END
 PORT
  LAYER ME4 ;
  RECT 473.449 35.220 473.789 280.651 ;
 END
 PORT
  LAYER ME4 ;
  RECT 471.447 35.220 471.787 280.651 ;
 END
 PORT
  LAYER ME4 ;
  RECT 469.445 35.220 469.785 280.651 ;
 END
 PORT
  LAYER ME4 ;
  RECT 467.443 35.220 467.783 280.651 ;
 END
 PORT
  LAYER ME4 ;
  RECT 481.457 35.220 481.797 280.651 ;
 END
 PORT
  LAYER ME4 ;
  RECT 479.455 35.220 479.795 280.651 ;
 END
 PORT
  LAYER ME4 ;
  RECT 477.453 35.220 477.793 280.651 ;
 END
 PORT
  LAYER ME4 ;
  RECT 475.451 35.220 475.791 280.651 ;
 END
 PORT
  LAYER ME4 ;
  RECT 489.465 35.220 489.805 280.651 ;
 END
 PORT
  LAYER ME4 ;
  RECT 487.463 35.220 487.803 280.651 ;
 END
 PORT
  LAYER ME4 ;
  RECT 485.461 35.220 485.801 280.651 ;
 END
 PORT
  LAYER ME4 ;
  RECT 483.459 35.220 483.799 280.651 ;
 END
 PORT
  LAYER ME4 ;
  RECT 497.473 35.220 497.813 280.651 ;
 END
 PORT
  LAYER ME4 ;
  RECT 495.471 35.220 495.811 280.651 ;
 END
 PORT
  LAYER ME4 ;
  RECT 493.469 35.220 493.809 280.651 ;
 END
 PORT
  LAYER ME4 ;
  RECT 491.467 35.220 491.807 280.651 ;
 END
 PORT
  LAYER ME4 ;
  RECT 505.481 35.220 505.821 280.651 ;
 END
 PORT
  LAYER ME4 ;
  RECT 503.479 35.220 503.819 280.651 ;
 END
 PORT
  LAYER ME4 ;
  RECT 501.477 35.220 501.817 280.651 ;
 END
 PORT
  LAYER ME4 ;
  RECT 499.475 35.220 499.815 280.651 ;
 END
 PORT
  LAYER ME4 ;
  RECT 513.489 35.220 513.829 280.651 ;
 END
 PORT
  LAYER ME4 ;
  RECT 511.487 35.220 511.827 280.651 ;
 END
 PORT
  LAYER ME4 ;
  RECT 509.485 35.220 509.825 280.651 ;
 END
 PORT
  LAYER ME4 ;
  RECT 507.483 35.220 507.823 280.651 ;
 END
 PORT
  LAYER ME4 ;
  RECT 521.497 35.220 521.837 280.651 ;
 END
 PORT
  LAYER ME4 ;
  RECT 519.495 35.220 519.835 280.651 ;
 END
 PORT
  LAYER ME4 ;
  RECT 517.493 35.220 517.833 280.651 ;
 END
 PORT
  LAYER ME4 ;
  RECT 515.491 35.220 515.831 280.651 ;
 END
 PORT
  LAYER ME4 ;
  RECT 529.505 35.220 529.845 280.651 ;
 END
 PORT
  LAYER ME4 ;
  RECT 527.503 35.220 527.843 280.651 ;
 END
 PORT
  LAYER ME4 ;
  RECT 525.501 35.220 525.841 280.651 ;
 END
 PORT
  LAYER ME4 ;
  RECT 523.499 35.220 523.839 280.651 ;
 END
 PORT
  LAYER ME4 ;
  RECT 537.513 35.220 537.853 280.651 ;
 END
 PORT
  LAYER ME4 ;
  RECT 535.511 35.220 535.851 280.651 ;
 END
 PORT
  LAYER ME4 ;
  RECT 533.509 35.220 533.849 280.651 ;
 END
 PORT
  LAYER ME4 ;
  RECT 531.507 35.220 531.847 280.651 ;
 END
 PORT
  LAYER ME4 ;
  RECT 545.521 35.220 545.861 280.651 ;
 END
 PORT
  LAYER ME4 ;
  RECT 543.519 35.220 543.859 280.651 ;
 END
 PORT
  LAYER ME4 ;
  RECT 541.517 35.220 541.857 280.651 ;
 END
 PORT
  LAYER ME4 ;
  RECT 539.515 35.220 539.855 280.651 ;
 END
 PORT
  LAYER ME4 ;
  RECT 553.529 35.220 553.869 280.651 ;
 END
 PORT
  LAYER ME4 ;
  RECT 551.527 35.220 551.867 280.651 ;
 END
 PORT
  LAYER ME4 ;
  RECT 549.525 35.220 549.865 280.651 ;
 END
 PORT
  LAYER ME4 ;
  RECT 547.523 35.220 547.863 280.651 ;
 END
 PORT
  LAYER ME4 ;
  RECT 9.748 35.220 10.088 280.651 ;
 END
 PORT
  LAYER ME4 ;
  RECT 7.746 35.220 8.086 280.651 ;
 END
 PORT
  LAYER ME4 ;
  RECT 5.744 35.220 6.084 280.651 ;
 END
 PORT
  LAYER ME4 ;
  RECT 3.742 35.220 4.082 280.651 ;
 END
 PORT
  LAYER ME4 ;
  RECT 17.756 35.220 18.096 280.651 ;
 END
 PORT
  LAYER ME4 ;
  RECT 15.754 35.220 16.094 280.651 ;
 END
 PORT
  LAYER ME4 ;
  RECT 13.752 35.220 14.092 280.651 ;
 END
 PORT
  LAYER ME4 ;
  RECT 11.750 35.220 12.090 280.651 ;
 END
 PORT
  LAYER ME4 ;
  RECT 25.764 35.220 26.104 280.651 ;
 END
 PORT
  LAYER ME4 ;
  RECT 23.762 35.220 24.102 280.651 ;
 END
 PORT
  LAYER ME4 ;
  RECT 21.760 35.220 22.100 280.651 ;
 END
 PORT
  LAYER ME4 ;
  RECT 19.758 35.220 20.098 280.651 ;
 END
 PORT
  LAYER ME4 ;
  RECT 33.772 35.220 34.112 280.651 ;
 END
 PORT
  LAYER ME4 ;
  RECT 31.770 35.220 32.110 280.651 ;
 END
 PORT
  LAYER ME4 ;
  RECT 29.768 35.220 30.108 280.651 ;
 END
 PORT
  LAYER ME4 ;
  RECT 27.766 35.220 28.106 280.651 ;
 END
 PORT
  LAYER ME4 ;
  RECT 41.780 35.220 42.120 280.651 ;
 END
 PORT
  LAYER ME4 ;
  RECT 39.778 35.220 40.118 280.651 ;
 END
 PORT
  LAYER ME4 ;
  RECT 37.776 35.220 38.116 280.651 ;
 END
 PORT
  LAYER ME4 ;
  RECT 35.774 35.220 36.114 280.651 ;
 END
 PORT
  LAYER ME4 ;
  RECT 49.788 35.220 50.128 280.651 ;
 END
 PORT
  LAYER ME4 ;
  RECT 47.786 35.220 48.126 280.651 ;
 END
 PORT
  LAYER ME4 ;
  RECT 45.784 35.220 46.124 280.651 ;
 END
 PORT
  LAYER ME4 ;
  RECT 43.782 35.220 44.122 280.651 ;
 END
 PORT
  LAYER ME4 ;
  RECT 57.796 35.220 58.136 280.651 ;
 END
 PORT
  LAYER ME4 ;
  RECT 55.794 35.220 56.134 280.651 ;
 END
 PORT
  LAYER ME4 ;
  RECT 53.792 35.220 54.132 280.651 ;
 END
 PORT
  LAYER ME4 ;
  RECT 51.790 35.220 52.130 280.651 ;
 END
 PORT
  LAYER ME4 ;
  RECT 65.804 35.220 66.144 280.651 ;
 END
 PORT
  LAYER ME4 ;
  RECT 63.802 35.220 64.142 280.651 ;
 END
 PORT
  LAYER ME4 ;
  RECT 61.800 35.220 62.140 280.651 ;
 END
 PORT
  LAYER ME4 ;
  RECT 59.798 35.220 60.138 280.651 ;
 END
 PORT
  LAYER ME4 ;
  RECT 73.812 35.220 74.152 280.651 ;
 END
 PORT
  LAYER ME4 ;
  RECT 71.810 35.220 72.150 280.651 ;
 END
 PORT
  LAYER ME4 ;
  RECT 69.808 35.220 70.148 280.651 ;
 END
 PORT
  LAYER ME4 ;
  RECT 67.806 35.220 68.146 280.651 ;
 END
 PORT
  LAYER ME4 ;
  RECT 81.820 35.220 82.160 280.651 ;
 END
 PORT
  LAYER ME4 ;
  RECT 79.818 35.220 80.158 280.651 ;
 END
 PORT
  LAYER ME4 ;
  RECT 77.816 35.220 78.156 280.651 ;
 END
 PORT
  LAYER ME4 ;
  RECT 75.814 35.220 76.154 280.651 ;
 END
 PORT
  LAYER ME4 ;
  RECT 89.828 35.220 90.168 280.651 ;
 END
 PORT
  LAYER ME4 ;
  RECT 87.826 35.220 88.166 280.651 ;
 END
 PORT
  LAYER ME4 ;
  RECT 85.824 35.220 86.164 280.651 ;
 END
 PORT
  LAYER ME4 ;
  RECT 83.822 35.220 84.162 280.651 ;
 END
 PORT
  LAYER ME4 ;
  RECT 97.836 35.220 98.176 280.651 ;
 END
 PORT
  LAYER ME4 ;
  RECT 95.834 35.220 96.174 280.651 ;
 END
 PORT
  LAYER ME4 ;
  RECT 93.832 35.220 94.172 280.651 ;
 END
 PORT
  LAYER ME4 ;
  RECT 91.830 35.220 92.170 280.651 ;
 END
 PORT
  LAYER ME4 ;
  RECT 105.844 35.220 106.184 280.651 ;
 END
 PORT
  LAYER ME4 ;
  RECT 103.842 35.220 104.182 280.651 ;
 END
 PORT
  LAYER ME4 ;
  RECT 101.840 35.220 102.180 280.651 ;
 END
 PORT
  LAYER ME4 ;
  RECT 99.838 35.220 100.178 280.651 ;
 END
 PORT
  LAYER ME4 ;
  RECT 113.852 35.220 114.192 280.651 ;
 END
 PORT
  LAYER ME4 ;
  RECT 111.850 35.220 112.190 280.651 ;
 END
 PORT
  LAYER ME4 ;
  RECT 109.848 35.220 110.188 280.651 ;
 END
 PORT
  LAYER ME4 ;
  RECT 107.846 35.220 108.186 280.651 ;
 END
 PORT
  LAYER ME4 ;
  RECT 121.860 35.220 122.200 280.651 ;
 END
 PORT
  LAYER ME4 ;
  RECT 119.858 35.220 120.198 280.651 ;
 END
 PORT
  LAYER ME4 ;
  RECT 117.856 35.220 118.196 280.651 ;
 END
 PORT
  LAYER ME4 ;
  RECT 115.854 35.220 116.194 280.651 ;
 END
 PORT
  LAYER ME4 ;
  RECT 129.868 35.220 130.208 280.651 ;
 END
 PORT
  LAYER ME4 ;
  RECT 127.866 35.220 128.206 280.651 ;
 END
 PORT
  LAYER ME4 ;
  RECT 125.864 35.220 126.204 280.651 ;
 END
 PORT
  LAYER ME4 ;
  RECT 123.862 35.220 124.202 280.651 ;
 END
 PORT
  LAYER ME4 ;
  RECT 137.876 35.220 138.216 280.651 ;
 END
 PORT
  LAYER ME4 ;
  RECT 135.874 35.220 136.214 280.651 ;
 END
 PORT
  LAYER ME4 ;
  RECT 133.872 35.220 134.212 280.651 ;
 END
 PORT
  LAYER ME4 ;
  RECT 131.870 35.220 132.210 280.651 ;
 END
 PORT
  LAYER ME4 ;
  RECT 145.884 35.220 146.224 280.651 ;
 END
 PORT
  LAYER ME4 ;
  RECT 143.882 35.220 144.222 280.651 ;
 END
 PORT
  LAYER ME4 ;
  RECT 141.880 35.220 142.220 280.651 ;
 END
 PORT
  LAYER ME4 ;
  RECT 139.878 35.220 140.218 280.651 ;
 END
 PORT
  LAYER ME4 ;
  RECT 153.892 35.220 154.232 280.651 ;
 END
 PORT
  LAYER ME4 ;
  RECT 151.890 35.220 152.230 280.651 ;
 END
 PORT
  LAYER ME4 ;
  RECT 149.888 35.220 150.228 280.651 ;
 END
 PORT
  LAYER ME4 ;
  RECT 147.886 35.220 148.226 280.651 ;
 END
 PORT
  LAYER ME4 ;
  RECT 161.900 35.220 162.240 280.651 ;
 END
 PORT
  LAYER ME4 ;
  RECT 159.898 35.220 160.238 280.651 ;
 END
 PORT
  LAYER ME4 ;
  RECT 157.896 35.220 158.236 280.651 ;
 END
 PORT
  LAYER ME4 ;
  RECT 155.894 35.220 156.234 280.651 ;
 END
 PORT
  LAYER ME4 ;
  RECT 169.908 35.220 170.248 280.651 ;
 END
 PORT
  LAYER ME4 ;
  RECT 167.906 35.220 168.246 280.651 ;
 END
 PORT
  LAYER ME4 ;
  RECT 165.904 35.220 166.244 280.651 ;
 END
 PORT
  LAYER ME4 ;
  RECT 163.902 35.220 164.242 280.651 ;
 END
 PORT
  LAYER ME4 ;
  RECT 177.916 35.220 178.256 280.651 ;
 END
 PORT
  LAYER ME4 ;
  RECT 175.914 35.220 176.254 280.651 ;
 END
 PORT
  LAYER ME4 ;
  RECT 173.912 35.220 174.252 280.651 ;
 END
 PORT
  LAYER ME4 ;
  RECT 171.910 35.220 172.250 280.651 ;
 END
 PORT
  LAYER ME4 ;
  RECT 185.924 35.220 186.264 280.651 ;
 END
 PORT
  LAYER ME4 ;
  RECT 183.922 35.220 184.262 280.651 ;
 END
 PORT
  LAYER ME4 ;
  RECT 181.920 35.220 182.260 280.651 ;
 END
 PORT
  LAYER ME4 ;
  RECT 179.918 35.220 180.258 280.651 ;
 END
 PORT
  LAYER ME4 ;
  RECT 193.932 35.220 194.272 280.651 ;
 END
 PORT
  LAYER ME4 ;
  RECT 191.930 35.220 192.270 280.651 ;
 END
 PORT
  LAYER ME4 ;
  RECT 189.928 35.220 190.268 280.651 ;
 END
 PORT
  LAYER ME4 ;
  RECT 187.926 35.220 188.266 280.651 ;
 END
 PORT
  LAYER ME4 ;
  RECT 201.940 35.220 202.280 280.651 ;
 END
 PORT
  LAYER ME4 ;
  RECT 199.938 35.220 200.278 280.651 ;
 END
 PORT
  LAYER ME4 ;
  RECT 197.936 35.220 198.276 280.651 ;
 END
 PORT
  LAYER ME4 ;
  RECT 195.934 35.220 196.274 280.651 ;
 END
 PORT
  LAYER ME4 ;
  RECT 209.948 35.220 210.288 280.651 ;
 END
 PORT
  LAYER ME4 ;
  RECT 207.946 35.220 208.286 280.651 ;
 END
 PORT
  LAYER ME4 ;
  RECT 205.944 35.220 206.284 280.651 ;
 END
 PORT
  LAYER ME4 ;
  RECT 203.942 35.220 204.282 280.651 ;
 END
 PORT
  LAYER ME4 ;
  RECT 217.956 35.220 218.296 280.651 ;
 END
 PORT
  LAYER ME4 ;
  RECT 215.954 35.220 216.294 280.651 ;
 END
 PORT
  LAYER ME4 ;
  RECT 213.952 35.220 214.292 280.651 ;
 END
 PORT
  LAYER ME4 ;
  RECT 211.950 35.220 212.290 280.651 ;
 END
 PORT
  LAYER ME4 ;
  RECT 225.964 35.220 226.304 280.651 ;
 END
 PORT
  LAYER ME4 ;
  RECT 223.962 35.220 224.302 280.651 ;
 END
 PORT
  LAYER ME4 ;
  RECT 221.960 35.220 222.300 280.651 ;
 END
 PORT
  LAYER ME4 ;
  RECT 219.958 35.220 220.298 280.651 ;
 END
 PORT
  LAYER ME4 ;
  RECT 233.972 35.220 234.312 280.651 ;
 END
 PORT
  LAYER ME4 ;
  RECT 231.970 35.220 232.310 280.651 ;
 END
 PORT
  LAYER ME4 ;
  RECT 229.968 35.220 230.308 280.651 ;
 END
 PORT
  LAYER ME4 ;
  RECT 227.966 35.220 228.306 280.651 ;
 END
 PORT
  LAYER ME4 ;
  RECT 241.980 35.220 242.320 280.651 ;
 END
 PORT
  LAYER ME4 ;
  RECT 239.978 35.220 240.318 280.651 ;
 END
 PORT
  LAYER ME4 ;
  RECT 237.976 35.220 238.316 280.651 ;
 END
 PORT
  LAYER ME4 ;
  RECT 235.974 35.220 236.314 280.651 ;
 END
 PORT
  LAYER ME4 ;
  RECT 249.988 35.220 250.328 280.651 ;
 END
 PORT
  LAYER ME4 ;
  RECT 247.986 35.220 248.326 280.651 ;
 END
 PORT
  LAYER ME4 ;
  RECT 245.984 35.220 246.324 280.651 ;
 END
 PORT
  LAYER ME4 ;
  RECT 243.982 35.220 244.322 280.651 ;
 END
 PORT
  LAYER ME4 ;
  RECT 257.996 35.220 258.336 280.651 ;
 END
 PORT
  LAYER ME4 ;
  RECT 255.994 35.220 256.334 280.651 ;
 END
 PORT
  LAYER ME4 ;
  RECT 253.992 35.220 254.332 280.651 ;
 END
 PORT
  LAYER ME4 ;
  RECT 251.990 35.220 252.330 280.651 ;
 END
END VCC
PIN GND
  DIRECTION INOUT ;
  USE GROUND ;
 PORT
  LAYER ME4 ;
  RECT 298.274 0.921 298.614 280.651 ;
 END
 PORT
  LAYER ME4 ;
  RECT 305.091 0.000 305.811 31.570 ;
 END
 PORT
  LAYER ME4 ;
  RECT 306.282 0.000 306.622 280.651 ;
 END
 PORT
  LAYER ME4 ;
  RECT 300.276 0.000 300.616 280.651 ;
 END
 PORT
  LAYER ME4 ;
  RECT 301.087 0.000 301.807 31.570 ;
 END
 PORT
  LAYER ME4 ;
  RECT 302.278 0.921 302.618 280.651 ;
 END
 PORT
  LAYER ME4 ;
  RECT 304.280 0.921 304.620 280.651 ;
 END
 PORT
  LAYER ME4 ;
  RECT 313.099 0.000 313.819 31.570 ;
 END
 PORT
  LAYER ME4 ;
  RECT 314.290 0.000 314.630 280.651 ;
 END
 PORT
  LAYER ME4 ;
  RECT 308.284 0.000 308.624 280.651 ;
 END
 PORT
  LAYER ME4 ;
  RECT 309.095 0.000 309.815 31.570 ;
 END
 PORT
  LAYER ME4 ;
  RECT 310.286 0.921 310.626 280.651 ;
 END
 PORT
  LAYER ME4 ;
  RECT 312.288 0.921 312.628 280.651 ;
 END
 PORT
  LAYER ME4 ;
  RECT 321.107 0.000 321.827 31.570 ;
 END
 PORT
  LAYER ME4 ;
  RECT 322.298 0.000 322.638 280.651 ;
 END
 PORT
  LAYER ME4 ;
  RECT 316.292 0.000 316.632 280.651 ;
 END
 PORT
  LAYER ME4 ;
  RECT 317.103 0.000 317.823 31.570 ;
 END
 PORT
  LAYER ME4 ;
  RECT 318.294 0.921 318.634 280.651 ;
 END
 PORT
  LAYER ME4 ;
  RECT 320.296 0.921 320.636 280.651 ;
 END
 PORT
  LAYER ME4 ;
  RECT 329.115 0.000 329.835 31.570 ;
 END
 PORT
  LAYER ME4 ;
  RECT 330.306 0.000 330.646 280.651 ;
 END
 PORT
  LAYER ME4 ;
  RECT 324.300 0.000 324.640 280.651 ;
 END
 PORT
  LAYER ME4 ;
  RECT 325.111 0.000 325.831 31.570 ;
 END
 PORT
  LAYER ME4 ;
  RECT 326.302 0.921 326.642 280.651 ;
 END
 PORT
  LAYER ME4 ;
  RECT 328.304 0.921 328.644 280.651 ;
 END
 PORT
  LAYER ME4 ;
  RECT 337.123 0.000 337.843 31.570 ;
 END
 PORT
  LAYER ME4 ;
  RECT 338.314 0.000 338.654 280.651 ;
 END
 PORT
  LAYER ME4 ;
  RECT 332.308 0.000 332.648 280.651 ;
 END
 PORT
  LAYER ME4 ;
  RECT 333.119 0.000 333.839 31.570 ;
 END
 PORT
  LAYER ME4 ;
  RECT 334.310 0.921 334.650 280.651 ;
 END
 PORT
  LAYER ME4 ;
  RECT 336.312 0.921 336.652 280.651 ;
 END
 PORT
  LAYER ME4 ;
  RECT 345.131 0.000 345.851 31.570 ;
 END
 PORT
  LAYER ME4 ;
  RECT 346.322 0.000 346.662 280.651 ;
 END
 PORT
  LAYER ME4 ;
  RECT 340.316 0.000 340.656 280.651 ;
 END
 PORT
  LAYER ME4 ;
  RECT 341.127 0.000 341.847 31.570 ;
 END
 PORT
  LAYER ME4 ;
  RECT 342.318 0.921 342.658 280.651 ;
 END
 PORT
  LAYER ME4 ;
  RECT 344.320 0.921 344.660 280.651 ;
 END
 PORT
  LAYER ME4 ;
  RECT 353.139 0.000 353.859 31.570 ;
 END
 PORT
  LAYER ME4 ;
  RECT 354.330 0.000 354.670 280.651 ;
 END
 PORT
  LAYER ME4 ;
  RECT 348.324 0.000 348.664 280.651 ;
 END
 PORT
  LAYER ME4 ;
  RECT 349.135 0.000 349.855 31.570 ;
 END
 PORT
  LAYER ME4 ;
  RECT 350.326 0.921 350.666 280.651 ;
 END
 PORT
  LAYER ME4 ;
  RECT 352.328 0.921 352.668 280.651 ;
 END
 PORT
  LAYER ME4 ;
  RECT 361.147 0.000 361.867 31.570 ;
 END
 PORT
  LAYER ME4 ;
  RECT 362.338 0.000 362.678 280.651 ;
 END
 PORT
  LAYER ME4 ;
  RECT 356.332 0.000 356.672 280.651 ;
 END
 PORT
  LAYER ME4 ;
  RECT 357.143 0.000 357.863 31.570 ;
 END
 PORT
  LAYER ME4 ;
  RECT 358.334 0.921 358.674 280.651 ;
 END
 PORT
  LAYER ME4 ;
  RECT 360.336 0.921 360.676 280.651 ;
 END
 PORT
  LAYER ME4 ;
  RECT 369.155 0.000 369.875 31.570 ;
 END
 PORT
  LAYER ME4 ;
  RECT 370.346 0.000 370.686 280.651 ;
 END
 PORT
  LAYER ME4 ;
  RECT 364.340 0.000 364.680 280.651 ;
 END
 PORT
  LAYER ME4 ;
  RECT 365.151 0.000 365.871 31.570 ;
 END
 PORT
  LAYER ME4 ;
  RECT 366.342 0.921 366.682 280.651 ;
 END
 PORT
  LAYER ME4 ;
  RECT 368.344 0.921 368.684 280.651 ;
 END
 PORT
  LAYER ME4 ;
  RECT 377.163 0.000 377.883 31.570 ;
 END
 PORT
  LAYER ME4 ;
  RECT 378.354 0.000 378.694 280.651 ;
 END
 PORT
  LAYER ME4 ;
  RECT 372.348 0.000 372.688 280.651 ;
 END
 PORT
  LAYER ME4 ;
  RECT 373.159 0.000 373.879 31.570 ;
 END
 PORT
  LAYER ME4 ;
  RECT 374.350 0.921 374.690 280.651 ;
 END
 PORT
  LAYER ME4 ;
  RECT 376.352 0.921 376.692 280.651 ;
 END
 PORT
  LAYER ME4 ;
  RECT 385.171 0.000 385.891 31.570 ;
 END
 PORT
  LAYER ME4 ;
  RECT 386.362 0.000 386.702 280.651 ;
 END
 PORT
  LAYER ME4 ;
  RECT 380.356 0.000 380.696 280.651 ;
 END
 PORT
  LAYER ME4 ;
  RECT 381.167 0.000 381.887 31.570 ;
 END
 PORT
  LAYER ME4 ;
  RECT 382.358 0.921 382.698 280.651 ;
 END
 PORT
  LAYER ME4 ;
  RECT 384.360 0.921 384.700 280.651 ;
 END
 PORT
  LAYER ME4 ;
  RECT 393.179 0.000 393.899 31.570 ;
 END
 PORT
  LAYER ME4 ;
  RECT 394.370 0.000 394.710 280.651 ;
 END
 PORT
  LAYER ME4 ;
  RECT 388.364 0.000 388.704 280.651 ;
 END
 PORT
  LAYER ME4 ;
  RECT 389.175 0.000 389.895 31.570 ;
 END
 PORT
  LAYER ME4 ;
  RECT 390.366 0.921 390.706 280.651 ;
 END
 PORT
  LAYER ME4 ;
  RECT 392.368 0.921 392.708 280.651 ;
 END
 PORT
  LAYER ME4 ;
  RECT 401.187 0.000 401.907 31.570 ;
 END
 PORT
  LAYER ME4 ;
  RECT 402.378 0.000 402.718 280.651 ;
 END
 PORT
  LAYER ME4 ;
  RECT 396.372 0.000 396.712 280.651 ;
 END
 PORT
  LAYER ME4 ;
  RECT 397.183 0.000 397.903 31.570 ;
 END
 PORT
  LAYER ME4 ;
  RECT 398.374 0.921 398.714 280.651 ;
 END
 PORT
  LAYER ME4 ;
  RECT 400.376 0.921 400.716 280.651 ;
 END
 PORT
  LAYER ME4 ;
  RECT 409.195 0.000 409.915 31.570 ;
 END
 PORT
  LAYER ME4 ;
  RECT 410.386 0.000 410.726 280.651 ;
 END
 PORT
  LAYER ME4 ;
  RECT 404.380 0.000 404.720 280.651 ;
 END
 PORT
  LAYER ME4 ;
  RECT 405.191 0.000 405.911 31.570 ;
 END
 PORT
  LAYER ME4 ;
  RECT 406.382 0.921 406.722 280.651 ;
 END
 PORT
  LAYER ME4 ;
  RECT 408.384 0.921 408.724 280.651 ;
 END
 PORT
  LAYER ME4 ;
  RECT 417.203 0.000 417.923 31.570 ;
 END
 PORT
  LAYER ME4 ;
  RECT 418.394 0.000 418.734 280.651 ;
 END
 PORT
  LAYER ME4 ;
  RECT 412.388 0.000 412.728 280.651 ;
 END
 PORT
  LAYER ME4 ;
  RECT 413.199 0.000 413.919 31.570 ;
 END
 PORT
  LAYER ME4 ;
  RECT 414.390 0.921 414.730 280.651 ;
 END
 PORT
  LAYER ME4 ;
  RECT 416.392 0.921 416.732 280.651 ;
 END
 PORT
  LAYER ME4 ;
  RECT 425.211 0.000 425.931 31.570 ;
 END
 PORT
  LAYER ME4 ;
  RECT 426.402 0.000 426.742 280.651 ;
 END
 PORT
  LAYER ME4 ;
  RECT 420.396 0.000 420.736 280.651 ;
 END
 PORT
  LAYER ME4 ;
  RECT 421.207 0.000 421.927 31.570 ;
 END
 PORT
  LAYER ME4 ;
  RECT 422.398 0.921 422.738 280.651 ;
 END
 PORT
  LAYER ME4 ;
  RECT 424.400 0.921 424.740 280.651 ;
 END
 PORT
  LAYER ME4 ;
  RECT 433.219 0.000 433.939 31.570 ;
 END
 PORT
  LAYER ME4 ;
  RECT 434.410 0.000 434.750 280.651 ;
 END
 PORT
  LAYER ME4 ;
  RECT 428.404 0.000 428.744 280.651 ;
 END
 PORT
  LAYER ME4 ;
  RECT 429.215 0.000 429.935 31.570 ;
 END
 PORT
  LAYER ME4 ;
  RECT 430.406 0.921 430.746 280.651 ;
 END
 PORT
  LAYER ME4 ;
  RECT 432.408 0.921 432.748 280.651 ;
 END
 PORT
  LAYER ME4 ;
  RECT 441.227 0.000 441.947 31.570 ;
 END
 PORT
  LAYER ME4 ;
  RECT 442.418 0.000 442.758 280.651 ;
 END
 PORT
  LAYER ME4 ;
  RECT 436.412 0.000 436.752 280.651 ;
 END
 PORT
  LAYER ME4 ;
  RECT 437.223 0.000 437.943 31.570 ;
 END
 PORT
  LAYER ME4 ;
  RECT 438.414 0.921 438.754 280.651 ;
 END
 PORT
  LAYER ME4 ;
  RECT 440.416 0.921 440.756 280.651 ;
 END
 PORT
  LAYER ME4 ;
  RECT 449.235 0.000 449.955 31.570 ;
 END
 PORT
  LAYER ME4 ;
  RECT 450.426 0.000 450.766 280.651 ;
 END
 PORT
  LAYER ME4 ;
  RECT 444.420 0.000 444.760 280.651 ;
 END
 PORT
  LAYER ME4 ;
  RECT 445.231 0.000 445.951 31.570 ;
 END
 PORT
  LAYER ME4 ;
  RECT 446.422 0.921 446.762 280.651 ;
 END
 PORT
  LAYER ME4 ;
  RECT 448.424 0.921 448.764 280.651 ;
 END
 PORT
  LAYER ME4 ;
  RECT 457.243 0.000 457.963 31.570 ;
 END
 PORT
  LAYER ME4 ;
  RECT 458.434 0.000 458.774 280.651 ;
 END
 PORT
  LAYER ME4 ;
  RECT 452.428 0.000 452.768 280.651 ;
 END
 PORT
  LAYER ME4 ;
  RECT 453.239 0.000 453.959 31.570 ;
 END
 PORT
  LAYER ME4 ;
  RECT 454.430 0.921 454.770 280.651 ;
 END
 PORT
  LAYER ME4 ;
  RECT 456.432 0.921 456.772 280.651 ;
 END
 PORT
  LAYER ME4 ;
  RECT 465.251 0.000 465.971 31.570 ;
 END
 PORT
  LAYER ME4 ;
  RECT 466.442 0.000 466.782 280.651 ;
 END
 PORT
  LAYER ME4 ;
  RECT 460.436 0.000 460.776 280.651 ;
 END
 PORT
  LAYER ME4 ;
  RECT 461.247 0.000 461.967 31.570 ;
 END
 PORT
  LAYER ME4 ;
  RECT 462.438 0.921 462.778 280.651 ;
 END
 PORT
  LAYER ME4 ;
  RECT 464.440 0.921 464.780 280.651 ;
 END
 PORT
  LAYER ME4 ;
  RECT 473.259 0.000 473.979 31.570 ;
 END
 PORT
  LAYER ME4 ;
  RECT 474.450 0.000 474.790 280.651 ;
 END
 PORT
  LAYER ME4 ;
  RECT 468.444 0.000 468.784 280.651 ;
 END
 PORT
  LAYER ME4 ;
  RECT 469.255 0.000 469.975 31.570 ;
 END
 PORT
  LAYER ME4 ;
  RECT 470.446 0.921 470.786 280.651 ;
 END
 PORT
  LAYER ME4 ;
  RECT 472.448 0.921 472.788 280.651 ;
 END
 PORT
  LAYER ME4 ;
  RECT 481.267 0.000 481.987 31.570 ;
 END
 PORT
  LAYER ME4 ;
  RECT 482.458 0.000 482.798 280.651 ;
 END
 PORT
  LAYER ME4 ;
  RECT 476.452 0.000 476.792 280.651 ;
 END
 PORT
  LAYER ME4 ;
  RECT 477.263 0.000 477.983 31.570 ;
 END
 PORT
  LAYER ME4 ;
  RECT 478.454 0.921 478.794 280.651 ;
 END
 PORT
  LAYER ME4 ;
  RECT 480.456 0.921 480.796 280.651 ;
 END
 PORT
  LAYER ME4 ;
  RECT 489.275 0.000 489.995 31.570 ;
 END
 PORT
  LAYER ME4 ;
  RECT 490.466 0.000 490.806 280.651 ;
 END
 PORT
  LAYER ME4 ;
  RECT 484.460 0.000 484.800 280.651 ;
 END
 PORT
  LAYER ME4 ;
  RECT 485.271 0.000 485.991 31.570 ;
 END
 PORT
  LAYER ME4 ;
  RECT 486.462 0.921 486.802 280.651 ;
 END
 PORT
  LAYER ME4 ;
  RECT 488.464 0.921 488.804 280.651 ;
 END
 PORT
  LAYER ME4 ;
  RECT 497.283 0.000 498.003 31.570 ;
 END
 PORT
  LAYER ME4 ;
  RECT 498.474 0.000 498.814 280.651 ;
 END
 PORT
  LAYER ME4 ;
  RECT 492.468 0.000 492.808 280.651 ;
 END
 PORT
  LAYER ME4 ;
  RECT 493.279 0.000 493.999 31.570 ;
 END
 PORT
  LAYER ME4 ;
  RECT 494.470 0.921 494.810 280.651 ;
 END
 PORT
  LAYER ME4 ;
  RECT 496.472 0.921 496.812 280.651 ;
 END
 PORT
  LAYER ME4 ;
  RECT 505.291 0.000 506.011 31.570 ;
 END
 PORT
  LAYER ME4 ;
  RECT 506.482 0.000 506.822 280.651 ;
 END
 PORT
  LAYER ME4 ;
  RECT 500.476 0.000 500.816 280.651 ;
 END
 PORT
  LAYER ME4 ;
  RECT 501.287 0.000 502.007 31.570 ;
 END
 PORT
  LAYER ME4 ;
  RECT 502.478 0.921 502.818 280.651 ;
 END
 PORT
  LAYER ME4 ;
  RECT 504.480 0.921 504.820 280.651 ;
 END
 PORT
  LAYER ME4 ;
  RECT 513.299 0.000 514.019 31.570 ;
 END
 PORT
  LAYER ME4 ;
  RECT 514.490 0.000 514.830 280.651 ;
 END
 PORT
  LAYER ME4 ;
  RECT 508.484 0.000 508.824 280.651 ;
 END
 PORT
  LAYER ME4 ;
  RECT 509.295 0.000 510.015 31.570 ;
 END
 PORT
  LAYER ME4 ;
  RECT 510.486 0.921 510.826 280.651 ;
 END
 PORT
  LAYER ME4 ;
  RECT 512.488 0.921 512.828 280.651 ;
 END
 PORT
  LAYER ME4 ;
  RECT 521.307 0.000 522.027 31.570 ;
 END
 PORT
  LAYER ME4 ;
  RECT 522.498 0.000 522.838 280.651 ;
 END
 PORT
  LAYER ME4 ;
  RECT 516.492 0.000 516.832 280.651 ;
 END
 PORT
  LAYER ME4 ;
  RECT 517.303 0.000 518.023 31.570 ;
 END
 PORT
  LAYER ME4 ;
  RECT 518.494 0.921 518.834 280.651 ;
 END
 PORT
  LAYER ME4 ;
  RECT 520.496 0.921 520.836 280.651 ;
 END
 PORT
  LAYER ME4 ;
  RECT 529.315 0.000 530.035 31.570 ;
 END
 PORT
  LAYER ME4 ;
  RECT 530.506 0.000 530.846 280.651 ;
 END
 PORT
  LAYER ME4 ;
  RECT 524.500 0.000 524.840 280.651 ;
 END
 PORT
  LAYER ME4 ;
  RECT 525.311 0.000 526.031 31.570 ;
 END
 PORT
  LAYER ME4 ;
  RECT 526.502 0.921 526.842 280.651 ;
 END
 PORT
  LAYER ME4 ;
  RECT 528.504 0.921 528.844 280.651 ;
 END
 PORT
  LAYER ME4 ;
  RECT 537.323 0.000 538.043 31.570 ;
 END
 PORT
  LAYER ME4 ;
  RECT 538.514 0.000 538.854 280.651 ;
 END
 PORT
  LAYER ME4 ;
  RECT 532.508 0.000 532.848 280.651 ;
 END
 PORT
  LAYER ME4 ;
  RECT 533.319 0.000 534.039 31.570 ;
 END
 PORT
  LAYER ME4 ;
  RECT 534.510 0.921 534.850 280.651 ;
 END
 PORT
  LAYER ME4 ;
  RECT 536.512 0.921 536.852 280.651 ;
 END
 PORT
  LAYER ME4 ;
  RECT 545.331 0.000 546.051 31.570 ;
 END
 PORT
  LAYER ME4 ;
  RECT 546.522 0.000 546.862 280.651 ;
 END
 PORT
  LAYER ME4 ;
  RECT 540.516 0.000 540.856 280.651 ;
 END
 PORT
  LAYER ME4 ;
  RECT 541.327 0.000 542.047 31.570 ;
 END
 PORT
  LAYER ME4 ;
  RECT 542.518 0.921 542.858 280.651 ;
 END
 PORT
  LAYER ME4 ;
  RECT 544.520 0.921 544.860 280.651 ;
 END
 PORT
  LAYER ME4 ;
  RECT 553.339 0.000 554.059 31.570 ;
 END
 PORT
  LAYER ME4 ;
  RECT 554.530 0.000 554.870 280.651 ;
 END
 PORT
  LAYER ME4 ;
  RECT 548.524 0.000 548.864 280.651 ;
 END
 PORT
  LAYER ME4 ;
  RECT 549.335 0.000 550.055 31.570 ;
 END
 PORT
  LAYER ME4 ;
  RECT 550.526 0.921 550.866 280.651 ;
 END
 PORT
  LAYER ME4 ;
  RECT 552.528 0.921 552.868 280.651 ;
 END
 PORT
  LAYER ME4 ;
  RECT 555.531 0.000 555.871 280.651 ;
 END
 PORT
  LAYER ME4 ;
  RECT 279.417 0.000 280.137 280.651 ;
 END
 PORT
  LAYER ME4 ;
  RECT 285.411 0.000 286.131 280.651 ;
 END
 PORT
  LAYER ME4 ;
  RECT 290.882 0.000 291.602 280.651 ;
 END
 PORT
  LAYER ME4 ;
  RECT 292.597 0.000 293.317 280.651 ;
 END
 PORT
  LAYER ME4 ;
  RECT 295.593 0.000 296.193 280.651 ;
 END
 PORT
  LAYER ME4 ;
  RECT 297.273 0.921 297.613 280.651 ;
 END
 PORT
  LAYER ME4 ;
  RECT 271.858 0.000 272.578 280.651 ;
 END
 PORT
  LAYER ME4 ;
  RECT 269.818 0.921 270.538 279.771 ;
 END
 PORT
  LAYER ME4 ;
  RECT 267.698 0.000 268.418 280.651 ;
 END
 PORT
  LAYER ME4 ;
  RECT 265.658 0.921 266.378 280.651 ;
 END
 PORT
  LAYER ME4 ;
  RECT 263.538 0.000 264.258 280.651 ;
 END
 PORT
  LAYER ME4 ;
  RECT 261.498 0.921 262.218 280.651 ;
 END
 PORT
  LAYER ME4 ;
  RECT 1.740 0.000 2.080 280.651 ;
 END
 PORT
  LAYER ME4 ;
  RECT 2.741 0.921 3.081 280.651 ;
 END
 PORT
  LAYER ME4 ;
  RECT 9.558 0.000 10.278 31.570 ;
 END
 PORT
  LAYER ME4 ;
  RECT 10.749 0.000 11.089 280.651 ;
 END
 PORT
  LAYER ME4 ;
  RECT 4.743 0.000 5.083 280.651 ;
 END
 PORT
  LAYER ME4 ;
  RECT 5.554 0.000 6.274 31.570 ;
 END
 PORT
  LAYER ME4 ;
  RECT 6.745 0.921 7.085 280.651 ;
 END
 PORT
  LAYER ME4 ;
  RECT 8.747 0.921 9.087 280.651 ;
 END
 PORT
  LAYER ME4 ;
  RECT 17.566 0.000 18.286 31.570 ;
 END
 PORT
  LAYER ME4 ;
  RECT 18.757 0.000 19.097 280.651 ;
 END
 PORT
  LAYER ME4 ;
  RECT 12.751 0.000 13.091 280.651 ;
 END
 PORT
  LAYER ME4 ;
  RECT 13.562 0.000 14.282 31.570 ;
 END
 PORT
  LAYER ME4 ;
  RECT 14.753 0.921 15.093 280.651 ;
 END
 PORT
  LAYER ME4 ;
  RECT 16.755 0.921 17.095 280.651 ;
 END
 PORT
  LAYER ME4 ;
  RECT 25.574 0.000 26.294 31.570 ;
 END
 PORT
  LAYER ME4 ;
  RECT 26.765 0.000 27.105 280.651 ;
 END
 PORT
  LAYER ME4 ;
  RECT 20.759 0.000 21.099 280.651 ;
 END
 PORT
  LAYER ME4 ;
  RECT 21.570 0.000 22.290 31.570 ;
 END
 PORT
  LAYER ME4 ;
  RECT 22.761 0.921 23.101 280.651 ;
 END
 PORT
  LAYER ME4 ;
  RECT 24.763 0.921 25.103 280.651 ;
 END
 PORT
  LAYER ME4 ;
  RECT 33.582 0.000 34.302 31.570 ;
 END
 PORT
  LAYER ME4 ;
  RECT 34.773 0.000 35.113 280.651 ;
 END
 PORT
  LAYER ME4 ;
  RECT 28.767 0.000 29.107 280.651 ;
 END
 PORT
  LAYER ME4 ;
  RECT 29.578 0.000 30.298 31.570 ;
 END
 PORT
  LAYER ME4 ;
  RECT 30.769 0.921 31.109 280.651 ;
 END
 PORT
  LAYER ME4 ;
  RECT 32.771 0.921 33.111 280.651 ;
 END
 PORT
  LAYER ME4 ;
  RECT 41.590 0.000 42.310 31.570 ;
 END
 PORT
  LAYER ME4 ;
  RECT 42.781 0.000 43.121 280.651 ;
 END
 PORT
  LAYER ME4 ;
  RECT 36.775 0.000 37.115 280.651 ;
 END
 PORT
  LAYER ME4 ;
  RECT 37.586 0.000 38.306 31.570 ;
 END
 PORT
  LAYER ME4 ;
  RECT 38.777 0.921 39.117 280.651 ;
 END
 PORT
  LAYER ME4 ;
  RECT 40.779 0.921 41.119 280.651 ;
 END
 PORT
  LAYER ME4 ;
  RECT 49.598 0.000 50.318 31.570 ;
 END
 PORT
  LAYER ME4 ;
  RECT 50.789 0.000 51.129 280.651 ;
 END
 PORT
  LAYER ME4 ;
  RECT 44.783 0.000 45.123 280.651 ;
 END
 PORT
  LAYER ME4 ;
  RECT 45.594 0.000 46.314 31.570 ;
 END
 PORT
  LAYER ME4 ;
  RECT 46.785 0.921 47.125 280.651 ;
 END
 PORT
  LAYER ME4 ;
  RECT 48.787 0.921 49.127 280.651 ;
 END
 PORT
  LAYER ME4 ;
  RECT 57.606 0.000 58.326 31.570 ;
 END
 PORT
  LAYER ME4 ;
  RECT 58.797 0.000 59.137 280.651 ;
 END
 PORT
  LAYER ME4 ;
  RECT 52.791 0.000 53.131 280.651 ;
 END
 PORT
  LAYER ME4 ;
  RECT 53.602 0.000 54.322 31.570 ;
 END
 PORT
  LAYER ME4 ;
  RECT 54.793 0.921 55.133 280.651 ;
 END
 PORT
  LAYER ME4 ;
  RECT 56.795 0.921 57.135 280.651 ;
 END
 PORT
  LAYER ME4 ;
  RECT 65.614 0.000 66.334 31.570 ;
 END
 PORT
  LAYER ME4 ;
  RECT 66.805 0.000 67.145 280.651 ;
 END
 PORT
  LAYER ME4 ;
  RECT 60.799 0.000 61.139 280.651 ;
 END
 PORT
  LAYER ME4 ;
  RECT 61.610 0.000 62.330 31.570 ;
 END
 PORT
  LAYER ME4 ;
  RECT 62.801 0.921 63.141 280.651 ;
 END
 PORT
  LAYER ME4 ;
  RECT 64.803 0.921 65.143 280.651 ;
 END
 PORT
  LAYER ME4 ;
  RECT 73.622 0.000 74.342 31.570 ;
 END
 PORT
  LAYER ME4 ;
  RECT 74.813 0.000 75.153 280.651 ;
 END
 PORT
  LAYER ME4 ;
  RECT 68.807 0.000 69.147 280.651 ;
 END
 PORT
  LAYER ME4 ;
  RECT 69.618 0.000 70.338 31.570 ;
 END
 PORT
  LAYER ME4 ;
  RECT 70.809 0.921 71.149 280.651 ;
 END
 PORT
  LAYER ME4 ;
  RECT 72.811 0.921 73.151 280.651 ;
 END
 PORT
  LAYER ME4 ;
  RECT 81.630 0.000 82.350 31.570 ;
 END
 PORT
  LAYER ME4 ;
  RECT 82.821 0.000 83.161 280.651 ;
 END
 PORT
  LAYER ME4 ;
  RECT 76.815 0.000 77.155 280.651 ;
 END
 PORT
  LAYER ME4 ;
  RECT 77.626 0.000 78.346 31.570 ;
 END
 PORT
  LAYER ME4 ;
  RECT 78.817 0.921 79.157 280.651 ;
 END
 PORT
  LAYER ME4 ;
  RECT 80.819 0.921 81.159 280.651 ;
 END
 PORT
  LAYER ME4 ;
  RECT 89.638 0.000 90.358 31.570 ;
 END
 PORT
  LAYER ME4 ;
  RECT 90.829 0.000 91.169 280.651 ;
 END
 PORT
  LAYER ME4 ;
  RECT 84.823 0.000 85.163 280.651 ;
 END
 PORT
  LAYER ME4 ;
  RECT 85.634 0.000 86.354 31.570 ;
 END
 PORT
  LAYER ME4 ;
  RECT 86.825 0.921 87.165 280.651 ;
 END
 PORT
  LAYER ME4 ;
  RECT 88.827 0.921 89.167 280.651 ;
 END
 PORT
  LAYER ME4 ;
  RECT 97.646 0.000 98.366 31.570 ;
 END
 PORT
  LAYER ME4 ;
  RECT 98.837 0.000 99.177 280.651 ;
 END
 PORT
  LAYER ME4 ;
  RECT 92.831 0.000 93.171 280.651 ;
 END
 PORT
  LAYER ME4 ;
  RECT 93.642 0.000 94.362 31.570 ;
 END
 PORT
  LAYER ME4 ;
  RECT 94.833 0.921 95.173 280.651 ;
 END
 PORT
  LAYER ME4 ;
  RECT 96.835 0.921 97.175 280.651 ;
 END
 PORT
  LAYER ME4 ;
  RECT 105.654 0.000 106.374 31.570 ;
 END
 PORT
  LAYER ME4 ;
  RECT 106.845 0.000 107.185 280.651 ;
 END
 PORT
  LAYER ME4 ;
  RECT 100.839 0.000 101.179 280.651 ;
 END
 PORT
  LAYER ME4 ;
  RECT 101.650 0.000 102.370 31.570 ;
 END
 PORT
  LAYER ME4 ;
  RECT 102.841 0.921 103.181 280.651 ;
 END
 PORT
  LAYER ME4 ;
  RECT 104.843 0.921 105.183 280.651 ;
 END
 PORT
  LAYER ME4 ;
  RECT 113.662 0.000 114.382 31.570 ;
 END
 PORT
  LAYER ME4 ;
  RECT 114.853 0.000 115.193 280.651 ;
 END
 PORT
  LAYER ME4 ;
  RECT 108.847 0.000 109.187 280.651 ;
 END
 PORT
  LAYER ME4 ;
  RECT 109.658 0.000 110.378 31.570 ;
 END
 PORT
  LAYER ME4 ;
  RECT 110.849 0.921 111.189 280.651 ;
 END
 PORT
  LAYER ME4 ;
  RECT 112.851 0.921 113.191 280.651 ;
 END
 PORT
  LAYER ME4 ;
  RECT 121.670 0.000 122.390 31.570 ;
 END
 PORT
  LAYER ME4 ;
  RECT 122.861 0.000 123.201 280.651 ;
 END
 PORT
  LAYER ME4 ;
  RECT 116.855 0.000 117.195 280.651 ;
 END
 PORT
  LAYER ME4 ;
  RECT 117.666 0.000 118.386 31.570 ;
 END
 PORT
  LAYER ME4 ;
  RECT 118.857 0.921 119.197 280.651 ;
 END
 PORT
  LAYER ME4 ;
  RECT 120.859 0.921 121.199 280.651 ;
 END
 PORT
  LAYER ME4 ;
  RECT 129.678 0.000 130.398 31.570 ;
 END
 PORT
  LAYER ME4 ;
  RECT 130.869 0.000 131.209 280.651 ;
 END
 PORT
  LAYER ME4 ;
  RECT 124.863 0.000 125.203 280.651 ;
 END
 PORT
  LAYER ME4 ;
  RECT 125.674 0.000 126.394 31.570 ;
 END
 PORT
  LAYER ME4 ;
  RECT 126.865 0.921 127.205 280.651 ;
 END
 PORT
  LAYER ME4 ;
  RECT 128.867 0.921 129.207 280.651 ;
 END
 PORT
  LAYER ME4 ;
  RECT 137.686 0.000 138.406 31.570 ;
 END
 PORT
  LAYER ME4 ;
  RECT 138.877 0.000 139.217 280.651 ;
 END
 PORT
  LAYER ME4 ;
  RECT 132.871 0.000 133.211 280.651 ;
 END
 PORT
  LAYER ME4 ;
  RECT 133.682 0.000 134.402 31.570 ;
 END
 PORT
  LAYER ME4 ;
  RECT 134.873 0.921 135.213 280.651 ;
 END
 PORT
  LAYER ME4 ;
  RECT 136.875 0.921 137.215 280.651 ;
 END
 PORT
  LAYER ME4 ;
  RECT 145.694 0.000 146.414 31.570 ;
 END
 PORT
  LAYER ME4 ;
  RECT 146.885 0.000 147.225 280.651 ;
 END
 PORT
  LAYER ME4 ;
  RECT 140.879 0.000 141.219 280.651 ;
 END
 PORT
  LAYER ME4 ;
  RECT 141.690 0.000 142.410 31.570 ;
 END
 PORT
  LAYER ME4 ;
  RECT 142.881 0.921 143.221 280.651 ;
 END
 PORT
  LAYER ME4 ;
  RECT 144.883 0.921 145.223 280.651 ;
 END
 PORT
  LAYER ME4 ;
  RECT 153.702 0.000 154.422 31.570 ;
 END
 PORT
  LAYER ME4 ;
  RECT 154.893 0.000 155.233 280.651 ;
 END
 PORT
  LAYER ME4 ;
  RECT 148.887 0.000 149.227 280.651 ;
 END
 PORT
  LAYER ME4 ;
  RECT 149.698 0.000 150.418 31.570 ;
 END
 PORT
  LAYER ME4 ;
  RECT 150.889 0.921 151.229 280.651 ;
 END
 PORT
  LAYER ME4 ;
  RECT 152.891 0.921 153.231 280.651 ;
 END
 PORT
  LAYER ME4 ;
  RECT 161.710 0.000 162.430 31.570 ;
 END
 PORT
  LAYER ME4 ;
  RECT 162.901 0.000 163.241 280.651 ;
 END
 PORT
  LAYER ME4 ;
  RECT 156.895 0.000 157.235 280.651 ;
 END
 PORT
  LAYER ME4 ;
  RECT 157.706 0.000 158.426 31.570 ;
 END
 PORT
  LAYER ME4 ;
  RECT 158.897 0.921 159.237 280.651 ;
 END
 PORT
  LAYER ME4 ;
  RECT 160.899 0.921 161.239 280.651 ;
 END
 PORT
  LAYER ME4 ;
  RECT 169.718 0.000 170.438 31.570 ;
 END
 PORT
  LAYER ME4 ;
  RECT 170.909 0.000 171.249 280.651 ;
 END
 PORT
  LAYER ME4 ;
  RECT 164.903 0.000 165.243 280.651 ;
 END
 PORT
  LAYER ME4 ;
  RECT 165.714 0.000 166.434 31.570 ;
 END
 PORT
  LAYER ME4 ;
  RECT 166.905 0.921 167.245 280.651 ;
 END
 PORT
  LAYER ME4 ;
  RECT 168.907 0.921 169.247 280.651 ;
 END
 PORT
  LAYER ME4 ;
  RECT 177.726 0.000 178.446 31.570 ;
 END
 PORT
  LAYER ME4 ;
  RECT 178.917 0.000 179.257 280.651 ;
 END
 PORT
  LAYER ME4 ;
  RECT 172.911 0.000 173.251 280.651 ;
 END
 PORT
  LAYER ME4 ;
  RECT 173.722 0.000 174.442 31.570 ;
 END
 PORT
  LAYER ME4 ;
  RECT 174.913 0.921 175.253 280.651 ;
 END
 PORT
  LAYER ME4 ;
  RECT 176.915 0.921 177.255 280.651 ;
 END
 PORT
  LAYER ME4 ;
  RECT 185.734 0.000 186.454 31.570 ;
 END
 PORT
  LAYER ME4 ;
  RECT 186.925 0.000 187.265 280.651 ;
 END
 PORT
  LAYER ME4 ;
  RECT 180.919 0.000 181.259 280.651 ;
 END
 PORT
  LAYER ME4 ;
  RECT 181.730 0.000 182.450 31.570 ;
 END
 PORT
  LAYER ME4 ;
  RECT 182.921 0.921 183.261 280.651 ;
 END
 PORT
  LAYER ME4 ;
  RECT 184.923 0.921 185.263 280.651 ;
 END
 PORT
  LAYER ME4 ;
  RECT 193.742 0.000 194.462 31.570 ;
 END
 PORT
  LAYER ME4 ;
  RECT 194.933 0.000 195.273 280.651 ;
 END
 PORT
  LAYER ME4 ;
  RECT 188.927 0.000 189.267 280.651 ;
 END
 PORT
  LAYER ME4 ;
  RECT 189.738 0.000 190.458 31.570 ;
 END
 PORT
  LAYER ME4 ;
  RECT 190.929 0.921 191.269 280.651 ;
 END
 PORT
  LAYER ME4 ;
  RECT 192.931 0.921 193.271 280.651 ;
 END
 PORT
  LAYER ME4 ;
  RECT 201.750 0.000 202.470 31.570 ;
 END
 PORT
  LAYER ME4 ;
  RECT 202.941 0.000 203.281 280.651 ;
 END
 PORT
  LAYER ME4 ;
  RECT 196.935 0.000 197.275 280.651 ;
 END
 PORT
  LAYER ME4 ;
  RECT 197.746 0.000 198.466 31.570 ;
 END
 PORT
  LAYER ME4 ;
  RECT 198.937 0.921 199.277 280.651 ;
 END
 PORT
  LAYER ME4 ;
  RECT 200.939 0.921 201.279 280.651 ;
 END
 PORT
  LAYER ME4 ;
  RECT 209.758 0.000 210.478 31.570 ;
 END
 PORT
  LAYER ME4 ;
  RECT 210.949 0.000 211.289 280.651 ;
 END
 PORT
  LAYER ME4 ;
  RECT 204.943 0.000 205.283 280.651 ;
 END
 PORT
  LAYER ME4 ;
  RECT 205.754 0.000 206.474 31.570 ;
 END
 PORT
  LAYER ME4 ;
  RECT 206.945 0.921 207.285 280.651 ;
 END
 PORT
  LAYER ME4 ;
  RECT 208.947 0.921 209.287 280.651 ;
 END
 PORT
  LAYER ME4 ;
  RECT 217.766 0.000 218.486 31.570 ;
 END
 PORT
  LAYER ME4 ;
  RECT 218.957 0.000 219.297 280.651 ;
 END
 PORT
  LAYER ME4 ;
  RECT 212.951 0.000 213.291 280.651 ;
 END
 PORT
  LAYER ME4 ;
  RECT 213.762 0.000 214.482 31.570 ;
 END
 PORT
  LAYER ME4 ;
  RECT 214.953 0.921 215.293 280.651 ;
 END
 PORT
  LAYER ME4 ;
  RECT 216.955 0.921 217.295 280.651 ;
 END
 PORT
  LAYER ME4 ;
  RECT 225.774 0.000 226.494 31.570 ;
 END
 PORT
  LAYER ME4 ;
  RECT 226.965 0.000 227.305 280.651 ;
 END
 PORT
  LAYER ME4 ;
  RECT 220.959 0.000 221.299 280.651 ;
 END
 PORT
  LAYER ME4 ;
  RECT 221.770 0.000 222.490 31.570 ;
 END
 PORT
  LAYER ME4 ;
  RECT 222.961 0.921 223.301 280.651 ;
 END
 PORT
  LAYER ME4 ;
  RECT 224.963 0.921 225.303 280.651 ;
 END
 PORT
  LAYER ME4 ;
  RECT 233.782 0.000 234.502 31.570 ;
 END
 PORT
  LAYER ME4 ;
  RECT 234.973 0.000 235.313 280.651 ;
 END
 PORT
  LAYER ME4 ;
  RECT 228.967 0.000 229.307 280.651 ;
 END
 PORT
  LAYER ME4 ;
  RECT 229.778 0.000 230.498 31.570 ;
 END
 PORT
  LAYER ME4 ;
  RECT 230.969 0.921 231.309 280.651 ;
 END
 PORT
  LAYER ME4 ;
  RECT 232.971 0.921 233.311 280.651 ;
 END
 PORT
  LAYER ME4 ;
  RECT 241.790 0.000 242.510 31.570 ;
 END
 PORT
  LAYER ME4 ;
  RECT 242.981 0.000 243.321 280.651 ;
 END
 PORT
  LAYER ME4 ;
  RECT 236.975 0.000 237.315 280.651 ;
 END
 PORT
  LAYER ME4 ;
  RECT 237.786 0.000 238.506 31.570 ;
 END
 PORT
  LAYER ME4 ;
  RECT 238.977 0.921 239.317 280.651 ;
 END
 PORT
  LAYER ME4 ;
  RECT 240.979 0.921 241.319 280.651 ;
 END
 PORT
  LAYER ME4 ;
  RECT 249.798 0.000 250.518 31.570 ;
 END
 PORT
  LAYER ME4 ;
  RECT 250.989 0.000 251.329 280.651 ;
 END
 PORT
  LAYER ME4 ;
  RECT 244.983 0.000 245.323 280.651 ;
 END
 PORT
  LAYER ME4 ;
  RECT 245.794 0.000 246.514 31.570 ;
 END
 PORT
  LAYER ME4 ;
  RECT 246.985 0.921 247.325 280.651 ;
 END
 PORT
  LAYER ME4 ;
  RECT 248.987 0.921 249.327 280.651 ;
 END
 PORT
  LAYER ME4 ;
  RECT 257.806 0.000 258.526 31.570 ;
 END
 PORT
  LAYER ME4 ;
  RECT 258.997 0.000 259.337 280.651 ;
 END
 PORT
  LAYER ME4 ;
  RECT 252.991 0.000 253.331 280.651 ;
 END
 PORT
  LAYER ME4 ;
  RECT 253.802 0.000 254.522 31.570 ;
 END
 PORT
  LAYER ME4 ;
  RECT 254.993 0.921 255.333 280.651 ;
 END
 PORT
  LAYER ME4 ;
  RECT 256.995 0.921 257.335 280.651 ;
 END
 PORT
  LAYER ME4 ;
  RECT 259.998 0.000 260.338 280.651 ;
 END
END GND
PIN DI31
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 256.854 0.000 257.134 0.720 ;
  LAYER ME3 ;
  RECT 256.854 0.000 257.134 0.720 ;
  LAYER ME2 ;
  RECT 256.854 0.000 257.134 0.720 ;
  LAYER ME1 ;
  RECT 256.854 0.000 257.134 0.720 ;
 END
 ANTENNAPARTIALMETALAREA                  0.805 LAYER ME1 ;
 ANTENNAGATEAREA                          0.072 LAYER ME1 ;
 ANTENNAGATEAREA                          0.072 LAYER ME2 ;
 ANTENNAGATEAREA                          0.072 LAYER ME3 ;
 ANTENNAGATEAREA                          0.072 LAYER ME4 ;
 ANTENNADIFFAREA                          0.218 LAYER ME1 ;
 ANTENNADIFFAREA                          0.218 LAYER ME2 ;
 ANTENNADIFFAREA                          0.218 LAYER ME3 ;
 ANTENNADIFFAREA                          0.218 LAYER ME4 ;
 ANTENNAMAXAREACAR                       13.984 LAYER ME1 ;
 ANTENNAMAXAREACAR                       16.784 LAYER ME2 ;
 ANTENNAMAXAREACAR                       19.584 LAYER ME3 ;
 ANTENNAMAXAREACAR                       22.384 LAYER ME4 ;
END DI31
PIN DO31
  DIRECTION OUTPUT ;
 PORT
  LAYER ME4 ;
  RECT 254.876 0.000 255.156 0.720 ;
  LAYER ME3 ;
  RECT 254.876 0.000 255.156 0.720 ;
  LAYER ME2 ;
  RECT 254.876 0.000 255.156 0.720 ;
  LAYER ME1 ;
  RECT 254.876 0.000 255.156 0.720 ;
 END
 ANTENNAPARTIALMETALAREA                  2.030 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME3 ;
 ANTENNADIFFAREA                          1.293 LAYER ME4 ;
END DO31
PIN DI30
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 248.846 0.000 249.126 0.720 ;
  LAYER ME3 ;
  RECT 248.846 0.000 249.126 0.720 ;
  LAYER ME2 ;
  RECT 248.846 0.000 249.126 0.720 ;
  LAYER ME1 ;
  RECT 248.846 0.000 249.126 0.720 ;
 END
 ANTENNAPARTIALMETALAREA                  0.805 LAYER ME1 ;
 ANTENNAGATEAREA                          0.072 LAYER ME1 ;
 ANTENNAGATEAREA                          0.072 LAYER ME2 ;
 ANTENNAGATEAREA                          0.072 LAYER ME3 ;
 ANTENNAGATEAREA                          0.072 LAYER ME4 ;
 ANTENNADIFFAREA                          0.218 LAYER ME1 ;
 ANTENNADIFFAREA                          0.218 LAYER ME2 ;
 ANTENNADIFFAREA                          0.218 LAYER ME3 ;
 ANTENNADIFFAREA                          0.218 LAYER ME4 ;
 ANTENNAMAXAREACAR                       13.984 LAYER ME1 ;
 ANTENNAMAXAREACAR                       16.784 LAYER ME2 ;
 ANTENNAMAXAREACAR                       19.584 LAYER ME3 ;
 ANTENNAMAXAREACAR                       22.384 LAYER ME4 ;
END DI30
PIN DO30
  DIRECTION OUTPUT ;
 PORT
  LAYER ME4 ;
  RECT 246.868 0.000 247.148 0.720 ;
  LAYER ME3 ;
  RECT 246.868 0.000 247.148 0.720 ;
  LAYER ME2 ;
  RECT 246.868 0.000 247.148 0.720 ;
  LAYER ME1 ;
  RECT 246.868 0.000 247.148 0.720 ;
 END
 ANTENNAPARTIALMETALAREA                  2.030 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME3 ;
 ANTENNADIFFAREA                          1.293 LAYER ME4 ;
END DO30
PIN DI29
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 240.838 0.000 241.118 0.720 ;
  LAYER ME3 ;
  RECT 240.838 0.000 241.118 0.720 ;
  LAYER ME2 ;
  RECT 240.838 0.000 241.118 0.720 ;
  LAYER ME1 ;
  RECT 240.838 0.000 241.118 0.720 ;
 END
 ANTENNAPARTIALMETALAREA                  0.805 LAYER ME1 ;
 ANTENNAGATEAREA                          0.072 LAYER ME1 ;
 ANTENNAGATEAREA                          0.072 LAYER ME2 ;
 ANTENNAGATEAREA                          0.072 LAYER ME3 ;
 ANTENNAGATEAREA                          0.072 LAYER ME4 ;
 ANTENNADIFFAREA                          0.218 LAYER ME1 ;
 ANTENNADIFFAREA                          0.218 LAYER ME2 ;
 ANTENNADIFFAREA                          0.218 LAYER ME3 ;
 ANTENNADIFFAREA                          0.218 LAYER ME4 ;
 ANTENNAMAXAREACAR                       13.984 LAYER ME1 ;
 ANTENNAMAXAREACAR                       16.784 LAYER ME2 ;
 ANTENNAMAXAREACAR                       19.584 LAYER ME3 ;
 ANTENNAMAXAREACAR                       22.384 LAYER ME4 ;
END DI29
PIN DO29
  DIRECTION OUTPUT ;
 PORT
  LAYER ME4 ;
  RECT 238.860 0.000 239.140 0.720 ;
  LAYER ME3 ;
  RECT 238.860 0.000 239.140 0.720 ;
  LAYER ME2 ;
  RECT 238.860 0.000 239.140 0.720 ;
  LAYER ME1 ;
  RECT 238.860 0.000 239.140 0.720 ;
 END
 ANTENNAPARTIALMETALAREA                  2.030 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME3 ;
 ANTENNADIFFAREA                          1.293 LAYER ME4 ;
END DO29
PIN DI28
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 232.830 0.000 233.110 0.720 ;
  LAYER ME3 ;
  RECT 232.830 0.000 233.110 0.720 ;
  LAYER ME2 ;
  RECT 232.830 0.000 233.110 0.720 ;
  LAYER ME1 ;
  RECT 232.830 0.000 233.110 0.720 ;
 END
 ANTENNAPARTIALMETALAREA                  0.805 LAYER ME1 ;
 ANTENNAGATEAREA                          0.072 LAYER ME1 ;
 ANTENNAGATEAREA                          0.072 LAYER ME2 ;
 ANTENNAGATEAREA                          0.072 LAYER ME3 ;
 ANTENNAGATEAREA                          0.072 LAYER ME4 ;
 ANTENNADIFFAREA                          0.218 LAYER ME1 ;
 ANTENNADIFFAREA                          0.218 LAYER ME2 ;
 ANTENNADIFFAREA                          0.218 LAYER ME3 ;
 ANTENNADIFFAREA                          0.218 LAYER ME4 ;
 ANTENNAMAXAREACAR                       13.984 LAYER ME1 ;
 ANTENNAMAXAREACAR                       16.784 LAYER ME2 ;
 ANTENNAMAXAREACAR                       19.584 LAYER ME3 ;
 ANTENNAMAXAREACAR                       22.384 LAYER ME4 ;
END DI28
PIN DO28
  DIRECTION OUTPUT ;
 PORT
  LAYER ME4 ;
  RECT 230.852 0.000 231.132 0.720 ;
  LAYER ME3 ;
  RECT 230.852 0.000 231.132 0.720 ;
  LAYER ME2 ;
  RECT 230.852 0.000 231.132 0.720 ;
  LAYER ME1 ;
  RECT 230.852 0.000 231.132 0.720 ;
 END
 ANTENNAPARTIALMETALAREA                  2.030 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME3 ;
 ANTENNADIFFAREA                          1.293 LAYER ME4 ;
END DO28
PIN DI27
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 224.822 0.000 225.102 0.720 ;
  LAYER ME3 ;
  RECT 224.822 0.000 225.102 0.720 ;
  LAYER ME2 ;
  RECT 224.822 0.000 225.102 0.720 ;
  LAYER ME1 ;
  RECT 224.822 0.000 225.102 0.720 ;
 END
 ANTENNAPARTIALMETALAREA                  0.805 LAYER ME1 ;
 ANTENNAGATEAREA                          0.072 LAYER ME1 ;
 ANTENNAGATEAREA                          0.072 LAYER ME2 ;
 ANTENNAGATEAREA                          0.072 LAYER ME3 ;
 ANTENNAGATEAREA                          0.072 LAYER ME4 ;
 ANTENNADIFFAREA                          0.218 LAYER ME1 ;
 ANTENNADIFFAREA                          0.218 LAYER ME2 ;
 ANTENNADIFFAREA                          0.218 LAYER ME3 ;
 ANTENNADIFFAREA                          0.218 LAYER ME4 ;
 ANTENNAMAXAREACAR                       13.984 LAYER ME1 ;
 ANTENNAMAXAREACAR                       16.784 LAYER ME2 ;
 ANTENNAMAXAREACAR                       19.584 LAYER ME3 ;
 ANTENNAMAXAREACAR                       22.384 LAYER ME4 ;
END DI27
PIN DO27
  DIRECTION OUTPUT ;
 PORT
  LAYER ME4 ;
  RECT 222.844 0.000 223.124 0.720 ;
  LAYER ME3 ;
  RECT 222.844 0.000 223.124 0.720 ;
  LAYER ME2 ;
  RECT 222.844 0.000 223.124 0.720 ;
  LAYER ME1 ;
  RECT 222.844 0.000 223.124 0.720 ;
 END
 ANTENNAPARTIALMETALAREA                  2.030 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME3 ;
 ANTENNADIFFAREA                          1.293 LAYER ME4 ;
END DO27
PIN DI26
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 216.814 0.000 217.094 0.720 ;
  LAYER ME3 ;
  RECT 216.814 0.000 217.094 0.720 ;
  LAYER ME2 ;
  RECT 216.814 0.000 217.094 0.720 ;
  LAYER ME1 ;
  RECT 216.814 0.000 217.094 0.720 ;
 END
 ANTENNAPARTIALMETALAREA                  0.805 LAYER ME1 ;
 ANTENNAGATEAREA                          0.072 LAYER ME1 ;
 ANTENNAGATEAREA                          0.072 LAYER ME2 ;
 ANTENNAGATEAREA                          0.072 LAYER ME3 ;
 ANTENNAGATEAREA                          0.072 LAYER ME4 ;
 ANTENNADIFFAREA                          0.218 LAYER ME1 ;
 ANTENNADIFFAREA                          0.218 LAYER ME2 ;
 ANTENNADIFFAREA                          0.218 LAYER ME3 ;
 ANTENNADIFFAREA                          0.218 LAYER ME4 ;
 ANTENNAMAXAREACAR                       13.984 LAYER ME1 ;
 ANTENNAMAXAREACAR                       16.784 LAYER ME2 ;
 ANTENNAMAXAREACAR                       19.584 LAYER ME3 ;
 ANTENNAMAXAREACAR                       22.384 LAYER ME4 ;
END DI26
PIN DO26
  DIRECTION OUTPUT ;
 PORT
  LAYER ME4 ;
  RECT 214.836 0.000 215.116 0.720 ;
  LAYER ME3 ;
  RECT 214.836 0.000 215.116 0.720 ;
  LAYER ME2 ;
  RECT 214.836 0.000 215.116 0.720 ;
  LAYER ME1 ;
  RECT 214.836 0.000 215.116 0.720 ;
 END
 ANTENNAPARTIALMETALAREA                  2.030 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME3 ;
 ANTENNADIFFAREA                          1.293 LAYER ME4 ;
END DO26
PIN DI25
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 208.806 0.000 209.086 0.720 ;
  LAYER ME3 ;
  RECT 208.806 0.000 209.086 0.720 ;
  LAYER ME2 ;
  RECT 208.806 0.000 209.086 0.720 ;
  LAYER ME1 ;
  RECT 208.806 0.000 209.086 0.720 ;
 END
 ANTENNAPARTIALMETALAREA                  0.805 LAYER ME1 ;
 ANTENNAGATEAREA                          0.072 LAYER ME1 ;
 ANTENNAGATEAREA                          0.072 LAYER ME2 ;
 ANTENNAGATEAREA                          0.072 LAYER ME3 ;
 ANTENNAGATEAREA                          0.072 LAYER ME4 ;
 ANTENNADIFFAREA                          0.218 LAYER ME1 ;
 ANTENNADIFFAREA                          0.218 LAYER ME2 ;
 ANTENNADIFFAREA                          0.218 LAYER ME3 ;
 ANTENNADIFFAREA                          0.218 LAYER ME4 ;
 ANTENNAMAXAREACAR                       13.984 LAYER ME1 ;
 ANTENNAMAXAREACAR                       16.784 LAYER ME2 ;
 ANTENNAMAXAREACAR                       19.584 LAYER ME3 ;
 ANTENNAMAXAREACAR                       22.384 LAYER ME4 ;
END DI25
PIN DO25
  DIRECTION OUTPUT ;
 PORT
  LAYER ME4 ;
  RECT 206.828 0.000 207.108 0.720 ;
  LAYER ME3 ;
  RECT 206.828 0.000 207.108 0.720 ;
  LAYER ME2 ;
  RECT 206.828 0.000 207.108 0.720 ;
  LAYER ME1 ;
  RECT 206.828 0.000 207.108 0.720 ;
 END
 ANTENNAPARTIALMETALAREA                  2.030 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME3 ;
 ANTENNADIFFAREA                          1.293 LAYER ME4 ;
END DO25
PIN DI24
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 200.798 0.000 201.078 0.720 ;
  LAYER ME3 ;
  RECT 200.798 0.000 201.078 0.720 ;
  LAYER ME2 ;
  RECT 200.798 0.000 201.078 0.720 ;
  LAYER ME1 ;
  RECT 200.798 0.000 201.078 0.720 ;
 END
 ANTENNAPARTIALMETALAREA                  0.522 LAYER ME1 ;
 ANTENNAGATEAREA                          0.072 LAYER ME1 ;
 ANTENNAGATEAREA                          0.072 LAYER ME2 ;
 ANTENNAGATEAREA                          0.072 LAYER ME3 ;
 ANTENNAGATEAREA                          0.072 LAYER ME4 ;
 ANTENNADIFFAREA                          0.218 LAYER ME1 ;
 ANTENNADIFFAREA                          0.218 LAYER ME2 ;
 ANTENNADIFFAREA                          0.218 LAYER ME3 ;
 ANTENNADIFFAREA                          0.218 LAYER ME4 ;
 ANTENNAMAXAREACAR                       10.048 LAYER ME1 ;
 ANTENNAMAXAREACAR                       12.848 LAYER ME2 ;
 ANTENNAMAXAREACAR                       15.648 LAYER ME3 ;
 ANTENNAMAXAREACAR                       18.448 LAYER ME4 ;
END DI24
PIN DO24
  DIRECTION OUTPUT ;
 PORT
  LAYER ME4 ;
  RECT 198.740 0.000 199.020 0.720 ;
  LAYER ME3 ;
  RECT 198.740 0.000 199.020 0.720 ;
  LAYER ME2 ;
  RECT 198.740 0.000 199.020 0.720 ;
  LAYER ME1 ;
  RECT 198.740 0.000 199.020 0.720 ;
 END
 ANTENNAPARTIALMETALAREA                  2.030 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME3 ;
 ANTENNADIFFAREA                          1.293 LAYER ME4 ;
END DO24
PIN WEB3
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 199.220 0.000 199.500 0.720 ;
  LAYER ME3 ;
  RECT 199.220 0.000 199.500 0.720 ;
  LAYER ME2 ;
  RECT 199.220 0.000 199.500 0.720 ;
  LAYER ME1 ;
  RECT 199.220 0.000 199.500 0.720 ;
 END
 ANTENNAPARTIALMETALAREA                  0.436 LAYER ME2 ;
 ANTENNAGATEAREA                          0.288 LAYER ME2 ;
 ANTENNAGATEAREA                          0.288 LAYER ME3 ;
 ANTENNAGATEAREA                          0.288 LAYER ME4 ;
 ANTENNADIFFAREA                          0.218 LAYER ME2 ;
 ANTENNADIFFAREA                          0.218 LAYER ME3 ;
 ANTENNADIFFAREA                          0.218 LAYER ME4 ;
 ANTENNAMAXAREACAR                        4.602 LAYER ME2 ;
 ANTENNAMAXAREACAR                        5.302 LAYER ME3 ;
 ANTENNAMAXAREACAR                        6.002 LAYER ME4 ;
END WEB3
PIN DI23
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 192.790 0.000 193.070 0.720 ;
  LAYER ME3 ;
  RECT 192.790 0.000 193.070 0.720 ;
  LAYER ME2 ;
  RECT 192.790 0.000 193.070 0.720 ;
  LAYER ME1 ;
  RECT 192.790 0.000 193.070 0.720 ;
 END
 ANTENNAPARTIALMETALAREA                  0.805 LAYER ME1 ;
 ANTENNAGATEAREA                          0.072 LAYER ME1 ;
 ANTENNAGATEAREA                          0.072 LAYER ME2 ;
 ANTENNAGATEAREA                          0.072 LAYER ME3 ;
 ANTENNAGATEAREA                          0.072 LAYER ME4 ;
 ANTENNADIFFAREA                          0.218 LAYER ME1 ;
 ANTENNADIFFAREA                          0.218 LAYER ME2 ;
 ANTENNADIFFAREA                          0.218 LAYER ME3 ;
 ANTENNADIFFAREA                          0.218 LAYER ME4 ;
 ANTENNAMAXAREACAR                       13.984 LAYER ME1 ;
 ANTENNAMAXAREACAR                       16.784 LAYER ME2 ;
 ANTENNAMAXAREACAR                       19.584 LAYER ME3 ;
 ANTENNAMAXAREACAR                       22.384 LAYER ME4 ;
END DI23
PIN DO23
  DIRECTION OUTPUT ;
 PORT
  LAYER ME4 ;
  RECT 190.812 0.000 191.092 0.720 ;
  LAYER ME3 ;
  RECT 190.812 0.000 191.092 0.720 ;
  LAYER ME2 ;
  RECT 190.812 0.000 191.092 0.720 ;
  LAYER ME1 ;
  RECT 190.812 0.000 191.092 0.720 ;
 END
 ANTENNAPARTIALMETALAREA                  2.030 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME3 ;
 ANTENNADIFFAREA                          1.293 LAYER ME4 ;
END DO23
PIN DI22
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 184.782 0.000 185.062 0.720 ;
  LAYER ME3 ;
  RECT 184.782 0.000 185.062 0.720 ;
  LAYER ME2 ;
  RECT 184.782 0.000 185.062 0.720 ;
  LAYER ME1 ;
  RECT 184.782 0.000 185.062 0.720 ;
 END
 ANTENNAPARTIALMETALAREA                  0.805 LAYER ME1 ;
 ANTENNAGATEAREA                          0.072 LAYER ME1 ;
 ANTENNAGATEAREA                          0.072 LAYER ME2 ;
 ANTENNAGATEAREA                          0.072 LAYER ME3 ;
 ANTENNAGATEAREA                          0.072 LAYER ME4 ;
 ANTENNADIFFAREA                          0.218 LAYER ME1 ;
 ANTENNADIFFAREA                          0.218 LAYER ME2 ;
 ANTENNADIFFAREA                          0.218 LAYER ME3 ;
 ANTENNADIFFAREA                          0.218 LAYER ME4 ;
 ANTENNAMAXAREACAR                       13.984 LAYER ME1 ;
 ANTENNAMAXAREACAR                       16.784 LAYER ME2 ;
 ANTENNAMAXAREACAR                       19.584 LAYER ME3 ;
 ANTENNAMAXAREACAR                       22.384 LAYER ME4 ;
END DI22
PIN DO22
  DIRECTION OUTPUT ;
 PORT
  LAYER ME4 ;
  RECT 182.804 0.000 183.084 0.720 ;
  LAYER ME3 ;
  RECT 182.804 0.000 183.084 0.720 ;
  LAYER ME2 ;
  RECT 182.804 0.000 183.084 0.720 ;
  LAYER ME1 ;
  RECT 182.804 0.000 183.084 0.720 ;
 END
 ANTENNAPARTIALMETALAREA                  2.030 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME3 ;
 ANTENNADIFFAREA                          1.293 LAYER ME4 ;
END DO22
PIN DI21
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 176.774 0.000 177.054 0.720 ;
  LAYER ME3 ;
  RECT 176.774 0.000 177.054 0.720 ;
  LAYER ME2 ;
  RECT 176.774 0.000 177.054 0.720 ;
  LAYER ME1 ;
  RECT 176.774 0.000 177.054 0.720 ;
 END
 ANTENNAPARTIALMETALAREA                  0.805 LAYER ME1 ;
 ANTENNAGATEAREA                          0.072 LAYER ME1 ;
 ANTENNAGATEAREA                          0.072 LAYER ME2 ;
 ANTENNAGATEAREA                          0.072 LAYER ME3 ;
 ANTENNAGATEAREA                          0.072 LAYER ME4 ;
 ANTENNADIFFAREA                          0.218 LAYER ME1 ;
 ANTENNADIFFAREA                          0.218 LAYER ME2 ;
 ANTENNADIFFAREA                          0.218 LAYER ME3 ;
 ANTENNADIFFAREA                          0.218 LAYER ME4 ;
 ANTENNAMAXAREACAR                       13.984 LAYER ME1 ;
 ANTENNAMAXAREACAR                       16.784 LAYER ME2 ;
 ANTENNAMAXAREACAR                       19.584 LAYER ME3 ;
 ANTENNAMAXAREACAR                       22.384 LAYER ME4 ;
END DI21
PIN DO21
  DIRECTION OUTPUT ;
 PORT
  LAYER ME4 ;
  RECT 174.796 0.000 175.076 0.720 ;
  LAYER ME3 ;
  RECT 174.796 0.000 175.076 0.720 ;
  LAYER ME2 ;
  RECT 174.796 0.000 175.076 0.720 ;
  LAYER ME1 ;
  RECT 174.796 0.000 175.076 0.720 ;
 END
 ANTENNAPARTIALMETALAREA                  2.030 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME3 ;
 ANTENNADIFFAREA                          1.293 LAYER ME4 ;
END DO21
PIN DI20
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 168.766 0.000 169.046 0.720 ;
  LAYER ME3 ;
  RECT 168.766 0.000 169.046 0.720 ;
  LAYER ME2 ;
  RECT 168.766 0.000 169.046 0.720 ;
  LAYER ME1 ;
  RECT 168.766 0.000 169.046 0.720 ;
 END
 ANTENNAPARTIALMETALAREA                  0.805 LAYER ME1 ;
 ANTENNAGATEAREA                          0.072 LAYER ME1 ;
 ANTENNAGATEAREA                          0.072 LAYER ME2 ;
 ANTENNAGATEAREA                          0.072 LAYER ME3 ;
 ANTENNAGATEAREA                          0.072 LAYER ME4 ;
 ANTENNADIFFAREA                          0.218 LAYER ME1 ;
 ANTENNADIFFAREA                          0.218 LAYER ME2 ;
 ANTENNADIFFAREA                          0.218 LAYER ME3 ;
 ANTENNADIFFAREA                          0.218 LAYER ME4 ;
 ANTENNAMAXAREACAR                       13.984 LAYER ME1 ;
 ANTENNAMAXAREACAR                       16.784 LAYER ME2 ;
 ANTENNAMAXAREACAR                       19.584 LAYER ME3 ;
 ANTENNAMAXAREACAR                       22.384 LAYER ME4 ;
END DI20
PIN DO20
  DIRECTION OUTPUT ;
 PORT
  LAYER ME4 ;
  RECT 166.788 0.000 167.068 0.720 ;
  LAYER ME3 ;
  RECT 166.788 0.000 167.068 0.720 ;
  LAYER ME2 ;
  RECT 166.788 0.000 167.068 0.720 ;
  LAYER ME1 ;
  RECT 166.788 0.000 167.068 0.720 ;
 END
 ANTENNAPARTIALMETALAREA                  2.030 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME3 ;
 ANTENNADIFFAREA                          1.293 LAYER ME4 ;
END DO20
PIN DI19
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 160.758 0.000 161.038 0.720 ;
  LAYER ME3 ;
  RECT 160.758 0.000 161.038 0.720 ;
  LAYER ME2 ;
  RECT 160.758 0.000 161.038 0.720 ;
  LAYER ME1 ;
  RECT 160.758 0.000 161.038 0.720 ;
 END
 ANTENNAPARTIALMETALAREA                  0.805 LAYER ME1 ;
 ANTENNAGATEAREA                          0.072 LAYER ME1 ;
 ANTENNAGATEAREA                          0.072 LAYER ME2 ;
 ANTENNAGATEAREA                          0.072 LAYER ME3 ;
 ANTENNAGATEAREA                          0.072 LAYER ME4 ;
 ANTENNADIFFAREA                          0.218 LAYER ME1 ;
 ANTENNADIFFAREA                          0.218 LAYER ME2 ;
 ANTENNADIFFAREA                          0.218 LAYER ME3 ;
 ANTENNADIFFAREA                          0.218 LAYER ME4 ;
 ANTENNAMAXAREACAR                       13.984 LAYER ME1 ;
 ANTENNAMAXAREACAR                       16.784 LAYER ME2 ;
 ANTENNAMAXAREACAR                       19.584 LAYER ME3 ;
 ANTENNAMAXAREACAR                       22.384 LAYER ME4 ;
END DI19
PIN DO19
  DIRECTION OUTPUT ;
 PORT
  LAYER ME4 ;
  RECT 158.780 0.000 159.060 0.720 ;
  LAYER ME3 ;
  RECT 158.780 0.000 159.060 0.720 ;
  LAYER ME2 ;
  RECT 158.780 0.000 159.060 0.720 ;
  LAYER ME1 ;
  RECT 158.780 0.000 159.060 0.720 ;
 END
 ANTENNAPARTIALMETALAREA                  2.030 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME3 ;
 ANTENNADIFFAREA                          1.293 LAYER ME4 ;
END DO19
PIN DI18
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 152.750 0.000 153.030 0.720 ;
  LAYER ME3 ;
  RECT 152.750 0.000 153.030 0.720 ;
  LAYER ME2 ;
  RECT 152.750 0.000 153.030 0.720 ;
  LAYER ME1 ;
  RECT 152.750 0.000 153.030 0.720 ;
 END
 ANTENNAPARTIALMETALAREA                  0.805 LAYER ME1 ;
 ANTENNAGATEAREA                          0.072 LAYER ME1 ;
 ANTENNAGATEAREA                          0.072 LAYER ME2 ;
 ANTENNAGATEAREA                          0.072 LAYER ME3 ;
 ANTENNAGATEAREA                          0.072 LAYER ME4 ;
 ANTENNADIFFAREA                          0.218 LAYER ME1 ;
 ANTENNADIFFAREA                          0.218 LAYER ME2 ;
 ANTENNADIFFAREA                          0.218 LAYER ME3 ;
 ANTENNADIFFAREA                          0.218 LAYER ME4 ;
 ANTENNAMAXAREACAR                       13.984 LAYER ME1 ;
 ANTENNAMAXAREACAR                       16.784 LAYER ME2 ;
 ANTENNAMAXAREACAR                       19.584 LAYER ME3 ;
 ANTENNAMAXAREACAR                       22.384 LAYER ME4 ;
END DI18
PIN DO18
  DIRECTION OUTPUT ;
 PORT
  LAYER ME4 ;
  RECT 150.772 0.000 151.052 0.720 ;
  LAYER ME3 ;
  RECT 150.772 0.000 151.052 0.720 ;
  LAYER ME2 ;
  RECT 150.772 0.000 151.052 0.720 ;
  LAYER ME1 ;
  RECT 150.772 0.000 151.052 0.720 ;
 END
 ANTENNAPARTIALMETALAREA                  2.030 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME3 ;
 ANTENNADIFFAREA                          1.293 LAYER ME4 ;
END DO18
PIN DI17
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 144.742 0.000 145.022 0.720 ;
  LAYER ME3 ;
  RECT 144.742 0.000 145.022 0.720 ;
  LAYER ME2 ;
  RECT 144.742 0.000 145.022 0.720 ;
  LAYER ME1 ;
  RECT 144.742 0.000 145.022 0.720 ;
 END
 ANTENNAPARTIALMETALAREA                  0.805 LAYER ME1 ;
 ANTENNAGATEAREA                          0.072 LAYER ME1 ;
 ANTENNAGATEAREA                          0.072 LAYER ME2 ;
 ANTENNAGATEAREA                          0.072 LAYER ME3 ;
 ANTENNAGATEAREA                          0.072 LAYER ME4 ;
 ANTENNADIFFAREA                          0.218 LAYER ME1 ;
 ANTENNADIFFAREA                          0.218 LAYER ME2 ;
 ANTENNADIFFAREA                          0.218 LAYER ME3 ;
 ANTENNADIFFAREA                          0.218 LAYER ME4 ;
 ANTENNAMAXAREACAR                       13.984 LAYER ME1 ;
 ANTENNAMAXAREACAR                       16.784 LAYER ME2 ;
 ANTENNAMAXAREACAR                       19.584 LAYER ME3 ;
 ANTENNAMAXAREACAR                       22.384 LAYER ME4 ;
END DI17
PIN DO17
  DIRECTION OUTPUT ;
 PORT
  LAYER ME4 ;
  RECT 142.764 0.000 143.044 0.720 ;
  LAYER ME3 ;
  RECT 142.764 0.000 143.044 0.720 ;
  LAYER ME2 ;
  RECT 142.764 0.000 143.044 0.720 ;
  LAYER ME1 ;
  RECT 142.764 0.000 143.044 0.720 ;
 END
 ANTENNAPARTIALMETALAREA                  2.030 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME3 ;
 ANTENNADIFFAREA                          1.293 LAYER ME4 ;
END DO17
PIN DI16
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 136.734 0.000 137.014 0.720 ;
  LAYER ME3 ;
  RECT 136.734 0.000 137.014 0.720 ;
  LAYER ME2 ;
  RECT 136.734 0.000 137.014 0.720 ;
  LAYER ME1 ;
  RECT 136.734 0.000 137.014 0.720 ;
 END
 ANTENNAPARTIALMETALAREA                  0.522 LAYER ME1 ;
 ANTENNAGATEAREA                          0.072 LAYER ME1 ;
 ANTENNAGATEAREA                          0.072 LAYER ME2 ;
 ANTENNAGATEAREA                          0.072 LAYER ME3 ;
 ANTENNAGATEAREA                          0.072 LAYER ME4 ;
 ANTENNADIFFAREA                          0.218 LAYER ME1 ;
 ANTENNADIFFAREA                          0.218 LAYER ME2 ;
 ANTENNADIFFAREA                          0.218 LAYER ME3 ;
 ANTENNADIFFAREA                          0.218 LAYER ME4 ;
 ANTENNAMAXAREACAR                       10.048 LAYER ME1 ;
 ANTENNAMAXAREACAR                       12.848 LAYER ME2 ;
 ANTENNAMAXAREACAR                       15.648 LAYER ME3 ;
 ANTENNAMAXAREACAR                       18.448 LAYER ME4 ;
END DI16
PIN DO16
  DIRECTION OUTPUT ;
 PORT
  LAYER ME4 ;
  RECT 134.676 0.000 134.956 0.720 ;
  LAYER ME3 ;
  RECT 134.676 0.000 134.956 0.720 ;
  LAYER ME2 ;
  RECT 134.676 0.000 134.956 0.720 ;
  LAYER ME1 ;
  RECT 134.676 0.000 134.956 0.720 ;
 END
 ANTENNAPARTIALMETALAREA                  2.030 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME3 ;
 ANTENNADIFFAREA                          1.293 LAYER ME4 ;
END DO16
PIN WEB2
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 135.156 0.000 135.436 0.720 ;
  LAYER ME3 ;
  RECT 135.156 0.000 135.436 0.720 ;
  LAYER ME2 ;
  RECT 135.156 0.000 135.436 0.720 ;
  LAYER ME1 ;
  RECT 135.156 0.000 135.436 0.720 ;
 END
 ANTENNAPARTIALMETALAREA                  0.436 LAYER ME2 ;
 ANTENNAGATEAREA                          0.288 LAYER ME2 ;
 ANTENNAGATEAREA                          0.288 LAYER ME3 ;
 ANTENNAGATEAREA                          0.288 LAYER ME4 ;
 ANTENNADIFFAREA                          0.218 LAYER ME2 ;
 ANTENNADIFFAREA                          0.218 LAYER ME3 ;
 ANTENNADIFFAREA                          0.218 LAYER ME4 ;
 ANTENNAMAXAREACAR                        4.602 LAYER ME2 ;
 ANTENNAMAXAREACAR                        5.302 LAYER ME3 ;
 ANTENNAMAXAREACAR                        6.002 LAYER ME4 ;
END WEB2
PIN DI15
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 128.726 0.000 129.006 0.720 ;
  LAYER ME3 ;
  RECT 128.726 0.000 129.006 0.720 ;
  LAYER ME2 ;
  RECT 128.726 0.000 129.006 0.720 ;
  LAYER ME1 ;
  RECT 128.726 0.000 129.006 0.720 ;
 END
 ANTENNAPARTIALMETALAREA                  0.805 LAYER ME1 ;
 ANTENNAGATEAREA                          0.072 LAYER ME1 ;
 ANTENNAGATEAREA                          0.072 LAYER ME2 ;
 ANTENNAGATEAREA                          0.072 LAYER ME3 ;
 ANTENNAGATEAREA                          0.072 LAYER ME4 ;
 ANTENNADIFFAREA                          0.218 LAYER ME1 ;
 ANTENNADIFFAREA                          0.218 LAYER ME2 ;
 ANTENNADIFFAREA                          0.218 LAYER ME3 ;
 ANTENNADIFFAREA                          0.218 LAYER ME4 ;
 ANTENNAMAXAREACAR                       13.984 LAYER ME1 ;
 ANTENNAMAXAREACAR                       16.784 LAYER ME2 ;
 ANTENNAMAXAREACAR                       19.584 LAYER ME3 ;
 ANTENNAMAXAREACAR                       22.384 LAYER ME4 ;
END DI15
PIN DO15
  DIRECTION OUTPUT ;
 PORT
  LAYER ME4 ;
  RECT 126.748 0.000 127.028 0.720 ;
  LAYER ME3 ;
  RECT 126.748 0.000 127.028 0.720 ;
  LAYER ME2 ;
  RECT 126.748 0.000 127.028 0.720 ;
  LAYER ME1 ;
  RECT 126.748 0.000 127.028 0.720 ;
 END
 ANTENNAPARTIALMETALAREA                  2.030 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME3 ;
 ANTENNADIFFAREA                          1.293 LAYER ME4 ;
END DO15
PIN DI14
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 120.718 0.000 120.998 0.720 ;
  LAYER ME3 ;
  RECT 120.718 0.000 120.998 0.720 ;
  LAYER ME2 ;
  RECT 120.718 0.000 120.998 0.720 ;
  LAYER ME1 ;
  RECT 120.718 0.000 120.998 0.720 ;
 END
 ANTENNAPARTIALMETALAREA                  0.805 LAYER ME1 ;
 ANTENNAGATEAREA                          0.072 LAYER ME1 ;
 ANTENNAGATEAREA                          0.072 LAYER ME2 ;
 ANTENNAGATEAREA                          0.072 LAYER ME3 ;
 ANTENNAGATEAREA                          0.072 LAYER ME4 ;
 ANTENNADIFFAREA                          0.218 LAYER ME1 ;
 ANTENNADIFFAREA                          0.218 LAYER ME2 ;
 ANTENNADIFFAREA                          0.218 LAYER ME3 ;
 ANTENNADIFFAREA                          0.218 LAYER ME4 ;
 ANTENNAMAXAREACAR                       13.984 LAYER ME1 ;
 ANTENNAMAXAREACAR                       16.784 LAYER ME2 ;
 ANTENNAMAXAREACAR                       19.584 LAYER ME3 ;
 ANTENNAMAXAREACAR                       22.384 LAYER ME4 ;
END DI14
PIN DO14
  DIRECTION OUTPUT ;
 PORT
  LAYER ME4 ;
  RECT 118.740 0.000 119.020 0.720 ;
  LAYER ME3 ;
  RECT 118.740 0.000 119.020 0.720 ;
  LAYER ME2 ;
  RECT 118.740 0.000 119.020 0.720 ;
  LAYER ME1 ;
  RECT 118.740 0.000 119.020 0.720 ;
 END
 ANTENNAPARTIALMETALAREA                  2.030 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME3 ;
 ANTENNADIFFAREA                          1.293 LAYER ME4 ;
END DO14
PIN DI13
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 112.710 0.000 112.990 0.720 ;
  LAYER ME3 ;
  RECT 112.710 0.000 112.990 0.720 ;
  LAYER ME2 ;
  RECT 112.710 0.000 112.990 0.720 ;
  LAYER ME1 ;
  RECT 112.710 0.000 112.990 0.720 ;
 END
 ANTENNAPARTIALMETALAREA                  0.805 LAYER ME1 ;
 ANTENNAGATEAREA                          0.072 LAYER ME1 ;
 ANTENNAGATEAREA                          0.072 LAYER ME2 ;
 ANTENNAGATEAREA                          0.072 LAYER ME3 ;
 ANTENNAGATEAREA                          0.072 LAYER ME4 ;
 ANTENNADIFFAREA                          0.218 LAYER ME1 ;
 ANTENNADIFFAREA                          0.218 LAYER ME2 ;
 ANTENNADIFFAREA                          0.218 LAYER ME3 ;
 ANTENNADIFFAREA                          0.218 LAYER ME4 ;
 ANTENNAMAXAREACAR                       13.984 LAYER ME1 ;
 ANTENNAMAXAREACAR                       16.784 LAYER ME2 ;
 ANTENNAMAXAREACAR                       19.584 LAYER ME3 ;
 ANTENNAMAXAREACAR                       22.384 LAYER ME4 ;
END DI13
PIN DO13
  DIRECTION OUTPUT ;
 PORT
  LAYER ME4 ;
  RECT 110.732 0.000 111.012 0.720 ;
  LAYER ME3 ;
  RECT 110.732 0.000 111.012 0.720 ;
  LAYER ME2 ;
  RECT 110.732 0.000 111.012 0.720 ;
  LAYER ME1 ;
  RECT 110.732 0.000 111.012 0.720 ;
 END
 ANTENNAPARTIALMETALAREA                  2.030 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME3 ;
 ANTENNADIFFAREA                          1.293 LAYER ME4 ;
END DO13
PIN DI12
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 104.702 0.000 104.982 0.720 ;
  LAYER ME3 ;
  RECT 104.702 0.000 104.982 0.720 ;
  LAYER ME2 ;
  RECT 104.702 0.000 104.982 0.720 ;
  LAYER ME1 ;
  RECT 104.702 0.000 104.982 0.720 ;
 END
 ANTENNAPARTIALMETALAREA                  0.805 LAYER ME1 ;
 ANTENNAGATEAREA                          0.072 LAYER ME1 ;
 ANTENNAGATEAREA                          0.072 LAYER ME2 ;
 ANTENNAGATEAREA                          0.072 LAYER ME3 ;
 ANTENNAGATEAREA                          0.072 LAYER ME4 ;
 ANTENNADIFFAREA                          0.218 LAYER ME1 ;
 ANTENNADIFFAREA                          0.218 LAYER ME2 ;
 ANTENNADIFFAREA                          0.218 LAYER ME3 ;
 ANTENNADIFFAREA                          0.218 LAYER ME4 ;
 ANTENNAMAXAREACAR                       13.984 LAYER ME1 ;
 ANTENNAMAXAREACAR                       16.784 LAYER ME2 ;
 ANTENNAMAXAREACAR                       19.584 LAYER ME3 ;
 ANTENNAMAXAREACAR                       22.384 LAYER ME4 ;
END DI12
PIN DO12
  DIRECTION OUTPUT ;
 PORT
  LAYER ME4 ;
  RECT 102.724 0.000 103.004 0.720 ;
  LAYER ME3 ;
  RECT 102.724 0.000 103.004 0.720 ;
  LAYER ME2 ;
  RECT 102.724 0.000 103.004 0.720 ;
  LAYER ME1 ;
  RECT 102.724 0.000 103.004 0.720 ;
 END
 ANTENNAPARTIALMETALAREA                  2.030 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME3 ;
 ANTENNADIFFAREA                          1.293 LAYER ME4 ;
END DO12
PIN DI11
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 96.694 0.000 96.974 0.720 ;
  LAYER ME3 ;
  RECT 96.694 0.000 96.974 0.720 ;
  LAYER ME2 ;
  RECT 96.694 0.000 96.974 0.720 ;
  LAYER ME1 ;
  RECT 96.694 0.000 96.974 0.720 ;
 END
 ANTENNAPARTIALMETALAREA                  0.805 LAYER ME1 ;
 ANTENNAGATEAREA                          0.072 LAYER ME1 ;
 ANTENNAGATEAREA                          0.072 LAYER ME2 ;
 ANTENNAGATEAREA                          0.072 LAYER ME3 ;
 ANTENNAGATEAREA                          0.072 LAYER ME4 ;
 ANTENNADIFFAREA                          0.218 LAYER ME1 ;
 ANTENNADIFFAREA                          0.218 LAYER ME2 ;
 ANTENNADIFFAREA                          0.218 LAYER ME3 ;
 ANTENNADIFFAREA                          0.218 LAYER ME4 ;
 ANTENNAMAXAREACAR                       13.984 LAYER ME1 ;
 ANTENNAMAXAREACAR                       16.784 LAYER ME2 ;
 ANTENNAMAXAREACAR                       19.584 LAYER ME3 ;
 ANTENNAMAXAREACAR                       22.384 LAYER ME4 ;
END DI11
PIN DO11
  DIRECTION OUTPUT ;
 PORT
  LAYER ME4 ;
  RECT 94.716 0.000 94.996 0.720 ;
  LAYER ME3 ;
  RECT 94.716 0.000 94.996 0.720 ;
  LAYER ME2 ;
  RECT 94.716 0.000 94.996 0.720 ;
  LAYER ME1 ;
  RECT 94.716 0.000 94.996 0.720 ;
 END
 ANTENNAPARTIALMETALAREA                  2.030 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME3 ;
 ANTENNADIFFAREA                          1.293 LAYER ME4 ;
END DO11
PIN DI10
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 88.686 0.000 88.966 0.720 ;
  LAYER ME3 ;
  RECT 88.686 0.000 88.966 0.720 ;
  LAYER ME2 ;
  RECT 88.686 0.000 88.966 0.720 ;
  LAYER ME1 ;
  RECT 88.686 0.000 88.966 0.720 ;
 END
 ANTENNAPARTIALMETALAREA                  0.805 LAYER ME1 ;
 ANTENNAGATEAREA                          0.072 LAYER ME1 ;
 ANTENNAGATEAREA                          0.072 LAYER ME2 ;
 ANTENNAGATEAREA                          0.072 LAYER ME3 ;
 ANTENNAGATEAREA                          0.072 LAYER ME4 ;
 ANTENNADIFFAREA                          0.218 LAYER ME1 ;
 ANTENNADIFFAREA                          0.218 LAYER ME2 ;
 ANTENNADIFFAREA                          0.218 LAYER ME3 ;
 ANTENNADIFFAREA                          0.218 LAYER ME4 ;
 ANTENNAMAXAREACAR                       13.984 LAYER ME1 ;
 ANTENNAMAXAREACAR                       16.784 LAYER ME2 ;
 ANTENNAMAXAREACAR                       19.584 LAYER ME3 ;
 ANTENNAMAXAREACAR                       22.384 LAYER ME4 ;
END DI10
PIN DO10
  DIRECTION OUTPUT ;
 PORT
  LAYER ME4 ;
  RECT 86.708 0.000 86.988 0.720 ;
  LAYER ME3 ;
  RECT 86.708 0.000 86.988 0.720 ;
  LAYER ME2 ;
  RECT 86.708 0.000 86.988 0.720 ;
  LAYER ME1 ;
  RECT 86.708 0.000 86.988 0.720 ;
 END
 ANTENNAPARTIALMETALAREA                  2.030 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME3 ;
 ANTENNADIFFAREA                          1.293 LAYER ME4 ;
END DO10
PIN DI9
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 80.678 0.000 80.958 0.720 ;
  LAYER ME3 ;
  RECT 80.678 0.000 80.958 0.720 ;
  LAYER ME2 ;
  RECT 80.678 0.000 80.958 0.720 ;
  LAYER ME1 ;
  RECT 80.678 0.000 80.958 0.720 ;
 END
 ANTENNAPARTIALMETALAREA                  0.805 LAYER ME1 ;
 ANTENNAGATEAREA                          0.072 LAYER ME1 ;
 ANTENNAGATEAREA                          0.072 LAYER ME2 ;
 ANTENNAGATEAREA                          0.072 LAYER ME3 ;
 ANTENNAGATEAREA                          0.072 LAYER ME4 ;
 ANTENNADIFFAREA                          0.218 LAYER ME1 ;
 ANTENNADIFFAREA                          0.218 LAYER ME2 ;
 ANTENNADIFFAREA                          0.218 LAYER ME3 ;
 ANTENNADIFFAREA                          0.218 LAYER ME4 ;
 ANTENNAMAXAREACAR                       13.984 LAYER ME1 ;
 ANTENNAMAXAREACAR                       16.784 LAYER ME2 ;
 ANTENNAMAXAREACAR                       19.584 LAYER ME3 ;
 ANTENNAMAXAREACAR                       22.384 LAYER ME4 ;
END DI9
PIN DO9
  DIRECTION OUTPUT ;
 PORT
  LAYER ME4 ;
  RECT 78.700 0.000 78.980 0.720 ;
  LAYER ME3 ;
  RECT 78.700 0.000 78.980 0.720 ;
  LAYER ME2 ;
  RECT 78.700 0.000 78.980 0.720 ;
  LAYER ME1 ;
  RECT 78.700 0.000 78.980 0.720 ;
 END
 ANTENNAPARTIALMETALAREA                  2.030 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME3 ;
 ANTENNADIFFAREA                          1.293 LAYER ME4 ;
END DO9
PIN DI8
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 72.670 0.000 72.950 0.720 ;
  LAYER ME3 ;
  RECT 72.670 0.000 72.950 0.720 ;
  LAYER ME2 ;
  RECT 72.670 0.000 72.950 0.720 ;
  LAYER ME1 ;
  RECT 72.670 0.000 72.950 0.720 ;
 END
 ANTENNAPARTIALMETALAREA                  0.522 LAYER ME1 ;
 ANTENNAGATEAREA                          0.072 LAYER ME1 ;
 ANTENNAGATEAREA                          0.072 LAYER ME2 ;
 ANTENNAGATEAREA                          0.072 LAYER ME3 ;
 ANTENNAGATEAREA                          0.072 LAYER ME4 ;
 ANTENNADIFFAREA                          0.218 LAYER ME1 ;
 ANTENNADIFFAREA                          0.218 LAYER ME2 ;
 ANTENNADIFFAREA                          0.218 LAYER ME3 ;
 ANTENNADIFFAREA                          0.218 LAYER ME4 ;
 ANTENNAMAXAREACAR                       10.048 LAYER ME1 ;
 ANTENNAMAXAREACAR                       12.848 LAYER ME2 ;
 ANTENNAMAXAREACAR                       15.648 LAYER ME3 ;
 ANTENNAMAXAREACAR                       18.448 LAYER ME4 ;
END DI8
PIN DO8
  DIRECTION OUTPUT ;
 PORT
  LAYER ME4 ;
  RECT 70.612 0.000 70.892 0.720 ;
  LAYER ME3 ;
  RECT 70.612 0.000 70.892 0.720 ;
  LAYER ME2 ;
  RECT 70.612 0.000 70.892 0.720 ;
  LAYER ME1 ;
  RECT 70.612 0.000 70.892 0.720 ;
 END
 ANTENNAPARTIALMETALAREA                  2.030 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME3 ;
 ANTENNADIFFAREA                          1.293 LAYER ME4 ;
END DO8
PIN WEB1
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 71.092 0.000 71.372 0.720 ;
  LAYER ME3 ;
  RECT 71.092 0.000 71.372 0.720 ;
  LAYER ME2 ;
  RECT 71.092 0.000 71.372 0.720 ;
  LAYER ME1 ;
  RECT 71.092 0.000 71.372 0.720 ;
 END
 ANTENNAPARTIALMETALAREA                  0.436 LAYER ME2 ;
 ANTENNAGATEAREA                          0.288 LAYER ME2 ;
 ANTENNAGATEAREA                          0.288 LAYER ME3 ;
 ANTENNAGATEAREA                          0.288 LAYER ME4 ;
 ANTENNADIFFAREA                          0.218 LAYER ME2 ;
 ANTENNADIFFAREA                          0.218 LAYER ME3 ;
 ANTENNADIFFAREA                          0.218 LAYER ME4 ;
 ANTENNAMAXAREACAR                        4.602 LAYER ME2 ;
 ANTENNAMAXAREACAR                        5.302 LAYER ME3 ;
 ANTENNAMAXAREACAR                        6.002 LAYER ME4 ;
END WEB1
PIN DI7
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 64.662 0.000 64.942 0.720 ;
  LAYER ME3 ;
  RECT 64.662 0.000 64.942 0.720 ;
  LAYER ME2 ;
  RECT 64.662 0.000 64.942 0.720 ;
  LAYER ME1 ;
  RECT 64.662 0.000 64.942 0.720 ;
 END
 ANTENNAPARTIALMETALAREA                  0.805 LAYER ME1 ;
 ANTENNAGATEAREA                          0.072 LAYER ME1 ;
 ANTENNAGATEAREA                          0.072 LAYER ME2 ;
 ANTENNAGATEAREA                          0.072 LAYER ME3 ;
 ANTENNAGATEAREA                          0.072 LAYER ME4 ;
 ANTENNADIFFAREA                          0.218 LAYER ME1 ;
 ANTENNADIFFAREA                          0.218 LAYER ME2 ;
 ANTENNADIFFAREA                          0.218 LAYER ME3 ;
 ANTENNADIFFAREA                          0.218 LAYER ME4 ;
 ANTENNAMAXAREACAR                       13.984 LAYER ME1 ;
 ANTENNAMAXAREACAR                       16.784 LAYER ME2 ;
 ANTENNAMAXAREACAR                       19.584 LAYER ME3 ;
 ANTENNAMAXAREACAR                       22.384 LAYER ME4 ;
END DI7
PIN DO7
  DIRECTION OUTPUT ;
 PORT
  LAYER ME4 ;
  RECT 62.684 0.000 62.964 0.720 ;
  LAYER ME3 ;
  RECT 62.684 0.000 62.964 0.720 ;
  LAYER ME2 ;
  RECT 62.684 0.000 62.964 0.720 ;
  LAYER ME1 ;
  RECT 62.684 0.000 62.964 0.720 ;
 END
 ANTENNAPARTIALMETALAREA                  2.030 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME3 ;
 ANTENNADIFFAREA                          1.293 LAYER ME4 ;
END DO7
PIN DI6
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 56.654 0.000 56.934 0.720 ;
  LAYER ME3 ;
  RECT 56.654 0.000 56.934 0.720 ;
  LAYER ME2 ;
  RECT 56.654 0.000 56.934 0.720 ;
  LAYER ME1 ;
  RECT 56.654 0.000 56.934 0.720 ;
 END
 ANTENNAPARTIALMETALAREA                  0.805 LAYER ME1 ;
 ANTENNAGATEAREA                          0.072 LAYER ME1 ;
 ANTENNAGATEAREA                          0.072 LAYER ME2 ;
 ANTENNAGATEAREA                          0.072 LAYER ME3 ;
 ANTENNAGATEAREA                          0.072 LAYER ME4 ;
 ANTENNADIFFAREA                          0.218 LAYER ME1 ;
 ANTENNADIFFAREA                          0.218 LAYER ME2 ;
 ANTENNADIFFAREA                          0.218 LAYER ME3 ;
 ANTENNADIFFAREA                          0.218 LAYER ME4 ;
 ANTENNAMAXAREACAR                       13.984 LAYER ME1 ;
 ANTENNAMAXAREACAR                       16.784 LAYER ME2 ;
 ANTENNAMAXAREACAR                       19.584 LAYER ME3 ;
 ANTENNAMAXAREACAR                       22.384 LAYER ME4 ;
END DI6
PIN DO6
  DIRECTION OUTPUT ;
 PORT
  LAYER ME4 ;
  RECT 54.676 0.000 54.956 0.720 ;
  LAYER ME3 ;
  RECT 54.676 0.000 54.956 0.720 ;
  LAYER ME2 ;
  RECT 54.676 0.000 54.956 0.720 ;
  LAYER ME1 ;
  RECT 54.676 0.000 54.956 0.720 ;
 END
 ANTENNAPARTIALMETALAREA                  2.030 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME3 ;
 ANTENNADIFFAREA                          1.293 LAYER ME4 ;
END DO6
PIN DI5
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 48.646 0.000 48.926 0.720 ;
  LAYER ME3 ;
  RECT 48.646 0.000 48.926 0.720 ;
  LAYER ME2 ;
  RECT 48.646 0.000 48.926 0.720 ;
  LAYER ME1 ;
  RECT 48.646 0.000 48.926 0.720 ;
 END
 ANTENNAPARTIALMETALAREA                  0.805 LAYER ME1 ;
 ANTENNAGATEAREA                          0.072 LAYER ME1 ;
 ANTENNAGATEAREA                          0.072 LAYER ME2 ;
 ANTENNAGATEAREA                          0.072 LAYER ME3 ;
 ANTENNAGATEAREA                          0.072 LAYER ME4 ;
 ANTENNADIFFAREA                          0.218 LAYER ME1 ;
 ANTENNADIFFAREA                          0.218 LAYER ME2 ;
 ANTENNADIFFAREA                          0.218 LAYER ME3 ;
 ANTENNADIFFAREA                          0.218 LAYER ME4 ;
 ANTENNAMAXAREACAR                       13.984 LAYER ME1 ;
 ANTENNAMAXAREACAR                       16.784 LAYER ME2 ;
 ANTENNAMAXAREACAR                       19.584 LAYER ME3 ;
 ANTENNAMAXAREACAR                       22.384 LAYER ME4 ;
END DI5
PIN DO5
  DIRECTION OUTPUT ;
 PORT
  LAYER ME4 ;
  RECT 46.668 0.000 46.948 0.720 ;
  LAYER ME3 ;
  RECT 46.668 0.000 46.948 0.720 ;
  LAYER ME2 ;
  RECT 46.668 0.000 46.948 0.720 ;
  LAYER ME1 ;
  RECT 46.668 0.000 46.948 0.720 ;
 END
 ANTENNAPARTIALMETALAREA                  2.030 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME3 ;
 ANTENNADIFFAREA                          1.293 LAYER ME4 ;
END DO5
PIN DI4
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 40.638 0.000 40.918 0.720 ;
  LAYER ME3 ;
  RECT 40.638 0.000 40.918 0.720 ;
  LAYER ME2 ;
  RECT 40.638 0.000 40.918 0.720 ;
  LAYER ME1 ;
  RECT 40.638 0.000 40.918 0.720 ;
 END
 ANTENNAPARTIALMETALAREA                  0.805 LAYER ME1 ;
 ANTENNAGATEAREA                          0.072 LAYER ME1 ;
 ANTENNAGATEAREA                          0.072 LAYER ME2 ;
 ANTENNAGATEAREA                          0.072 LAYER ME3 ;
 ANTENNAGATEAREA                          0.072 LAYER ME4 ;
 ANTENNADIFFAREA                          0.218 LAYER ME1 ;
 ANTENNADIFFAREA                          0.218 LAYER ME2 ;
 ANTENNADIFFAREA                          0.218 LAYER ME3 ;
 ANTENNADIFFAREA                          0.218 LAYER ME4 ;
 ANTENNAMAXAREACAR                       13.984 LAYER ME1 ;
 ANTENNAMAXAREACAR                       16.784 LAYER ME2 ;
 ANTENNAMAXAREACAR                       19.584 LAYER ME3 ;
 ANTENNAMAXAREACAR                       22.384 LAYER ME4 ;
END DI4
PIN DO4
  DIRECTION OUTPUT ;
 PORT
  LAYER ME4 ;
  RECT 38.660 0.000 38.940 0.720 ;
  LAYER ME3 ;
  RECT 38.660 0.000 38.940 0.720 ;
  LAYER ME2 ;
  RECT 38.660 0.000 38.940 0.720 ;
  LAYER ME1 ;
  RECT 38.660 0.000 38.940 0.720 ;
 END
 ANTENNAPARTIALMETALAREA                  2.030 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME3 ;
 ANTENNADIFFAREA                          1.293 LAYER ME4 ;
END DO4
PIN DI3
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 32.630 0.000 32.910 0.720 ;
  LAYER ME3 ;
  RECT 32.630 0.000 32.910 0.720 ;
  LAYER ME2 ;
  RECT 32.630 0.000 32.910 0.720 ;
  LAYER ME1 ;
  RECT 32.630 0.000 32.910 0.720 ;
 END
 ANTENNAPARTIALMETALAREA                  0.805 LAYER ME1 ;
 ANTENNAGATEAREA                          0.072 LAYER ME1 ;
 ANTENNAGATEAREA                          0.072 LAYER ME2 ;
 ANTENNAGATEAREA                          0.072 LAYER ME3 ;
 ANTENNAGATEAREA                          0.072 LAYER ME4 ;
 ANTENNADIFFAREA                          0.218 LAYER ME1 ;
 ANTENNADIFFAREA                          0.218 LAYER ME2 ;
 ANTENNADIFFAREA                          0.218 LAYER ME3 ;
 ANTENNADIFFAREA                          0.218 LAYER ME4 ;
 ANTENNAMAXAREACAR                       13.984 LAYER ME1 ;
 ANTENNAMAXAREACAR                       16.784 LAYER ME2 ;
 ANTENNAMAXAREACAR                       19.584 LAYER ME3 ;
 ANTENNAMAXAREACAR                       22.384 LAYER ME4 ;
END DI3
PIN DO3
  DIRECTION OUTPUT ;
 PORT
  LAYER ME4 ;
  RECT 30.652 0.000 30.932 0.720 ;
  LAYER ME3 ;
  RECT 30.652 0.000 30.932 0.720 ;
  LAYER ME2 ;
  RECT 30.652 0.000 30.932 0.720 ;
  LAYER ME1 ;
  RECT 30.652 0.000 30.932 0.720 ;
 END
 ANTENNAPARTIALMETALAREA                  2.030 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME3 ;
 ANTENNADIFFAREA                          1.293 LAYER ME4 ;
END DO3
PIN DI2
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 24.622 0.000 24.902 0.720 ;
  LAYER ME3 ;
  RECT 24.622 0.000 24.902 0.720 ;
  LAYER ME2 ;
  RECT 24.622 0.000 24.902 0.720 ;
  LAYER ME1 ;
  RECT 24.622 0.000 24.902 0.720 ;
 END
 ANTENNAPARTIALMETALAREA                  0.805 LAYER ME1 ;
 ANTENNAGATEAREA                          0.072 LAYER ME1 ;
 ANTENNAGATEAREA                          0.072 LAYER ME2 ;
 ANTENNAGATEAREA                          0.072 LAYER ME3 ;
 ANTENNAGATEAREA                          0.072 LAYER ME4 ;
 ANTENNADIFFAREA                          0.218 LAYER ME1 ;
 ANTENNADIFFAREA                          0.218 LAYER ME2 ;
 ANTENNADIFFAREA                          0.218 LAYER ME3 ;
 ANTENNADIFFAREA                          0.218 LAYER ME4 ;
 ANTENNAMAXAREACAR                       13.984 LAYER ME1 ;
 ANTENNAMAXAREACAR                       16.784 LAYER ME2 ;
 ANTENNAMAXAREACAR                       19.584 LAYER ME3 ;
 ANTENNAMAXAREACAR                       22.384 LAYER ME4 ;
END DI2
PIN DO2
  DIRECTION OUTPUT ;
 PORT
  LAYER ME4 ;
  RECT 22.644 0.000 22.924 0.720 ;
  LAYER ME3 ;
  RECT 22.644 0.000 22.924 0.720 ;
  LAYER ME2 ;
  RECT 22.644 0.000 22.924 0.720 ;
  LAYER ME1 ;
  RECT 22.644 0.000 22.924 0.720 ;
 END
 ANTENNAPARTIALMETALAREA                  2.030 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME3 ;
 ANTENNADIFFAREA                          1.293 LAYER ME4 ;
END DO2
PIN DI1
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 16.614 0.000 16.894 0.720 ;
  LAYER ME3 ;
  RECT 16.614 0.000 16.894 0.720 ;
  LAYER ME2 ;
  RECT 16.614 0.000 16.894 0.720 ;
  LAYER ME1 ;
  RECT 16.614 0.000 16.894 0.720 ;
 END
 ANTENNAPARTIALMETALAREA                  0.805 LAYER ME1 ;
 ANTENNAGATEAREA                          0.072 LAYER ME1 ;
 ANTENNAGATEAREA                          0.072 LAYER ME2 ;
 ANTENNAGATEAREA                          0.072 LAYER ME3 ;
 ANTENNAGATEAREA                          0.072 LAYER ME4 ;
 ANTENNADIFFAREA                          0.218 LAYER ME1 ;
 ANTENNADIFFAREA                          0.218 LAYER ME2 ;
 ANTENNADIFFAREA                          0.218 LAYER ME3 ;
 ANTENNADIFFAREA                          0.218 LAYER ME4 ;
 ANTENNAMAXAREACAR                       13.984 LAYER ME1 ;
 ANTENNAMAXAREACAR                       16.784 LAYER ME2 ;
 ANTENNAMAXAREACAR                       19.584 LAYER ME3 ;
 ANTENNAMAXAREACAR                       22.384 LAYER ME4 ;
END DI1
PIN DO1
  DIRECTION OUTPUT ;
 PORT
  LAYER ME4 ;
  RECT 14.636 0.000 14.916 0.720 ;
  LAYER ME3 ;
  RECT 14.636 0.000 14.916 0.720 ;
  LAYER ME2 ;
  RECT 14.636 0.000 14.916 0.720 ;
  LAYER ME1 ;
  RECT 14.636 0.000 14.916 0.720 ;
 END
 ANTENNAPARTIALMETALAREA                  2.030 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME3 ;
 ANTENNADIFFAREA                          1.293 LAYER ME4 ;
END DO1
PIN DI0
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 8.606 0.000 8.886 0.720 ;
  LAYER ME3 ;
  RECT 8.606 0.000 8.886 0.720 ;
  LAYER ME2 ;
  RECT 8.606 0.000 8.886 0.720 ;
  LAYER ME1 ;
  RECT 8.606 0.000 8.886 0.720 ;
 END
 ANTENNAPARTIALMETALAREA                  0.522 LAYER ME1 ;
 ANTENNAGATEAREA                          0.072 LAYER ME1 ;
 ANTENNAGATEAREA                          0.072 LAYER ME2 ;
 ANTENNAGATEAREA                          0.072 LAYER ME3 ;
 ANTENNAGATEAREA                          0.072 LAYER ME4 ;
 ANTENNADIFFAREA                          0.218 LAYER ME1 ;
 ANTENNADIFFAREA                          0.218 LAYER ME2 ;
 ANTENNADIFFAREA                          0.218 LAYER ME3 ;
 ANTENNADIFFAREA                          0.218 LAYER ME4 ;
 ANTENNAMAXAREACAR                       10.048 LAYER ME1 ;
 ANTENNAMAXAREACAR                       12.848 LAYER ME2 ;
 ANTENNAMAXAREACAR                       15.648 LAYER ME3 ;
 ANTENNAMAXAREACAR                       18.448 LAYER ME4 ;
END DI0
PIN DO0
  DIRECTION OUTPUT ;
 PORT
  LAYER ME4 ;
  RECT 6.548 0.000 6.828 0.720 ;
  LAYER ME3 ;
  RECT 6.548 0.000 6.828 0.720 ;
  LAYER ME2 ;
  RECT 6.548 0.000 6.828 0.720 ;
  LAYER ME1 ;
  RECT 6.548 0.000 6.828 0.720 ;
 END
 ANTENNAPARTIALMETALAREA                  2.030 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME3 ;
 ANTENNADIFFAREA                          1.293 LAYER ME4 ;
END DO0
PIN WEB0
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 7.028 0.000 7.308 0.720 ;
  LAYER ME3 ;
  RECT 7.028 0.000 7.308 0.720 ;
  LAYER ME2 ;
  RECT 7.028 0.000 7.308 0.720 ;
  LAYER ME1 ;
  RECT 7.028 0.000 7.308 0.720 ;
 END
 ANTENNAPARTIALMETALAREA                  0.436 LAYER ME2 ;
 ANTENNAGATEAREA                          0.288 LAYER ME2 ;
 ANTENNAGATEAREA                          0.288 LAYER ME3 ;
 ANTENNAGATEAREA                          0.288 LAYER ME4 ;
 ANTENNADIFFAREA                          0.218 LAYER ME2 ;
 ANTENNADIFFAREA                          0.218 LAYER ME3 ;
 ANTENNADIFFAREA                          0.218 LAYER ME4 ;
 ANTENNAMAXAREACAR                        4.602 LAYER ME2 ;
 ANTENNAMAXAREACAR                        5.302 LAYER ME3 ;
 ANTENNAMAXAREACAR                        6.002 LAYER ME4 ;
END WEB0
PIN A2
  DIRECTION INPUT ;
 PORT
  LAYER ME3 ;
  RECT 276.740 0.000 277.060 0.600 ;
  LAYER ME2 ;
  RECT 276.740 0.000 277.060 0.600 ;
  LAYER ME1 ;
  RECT 276.740 0.000 277.060 0.600 ;
 END
 ANTENNAPARTIALMETALAREA                  1.067 LAYER ME2 ;
 ANTENNAGATEAREA                          0.144 LAYER ME2 ;
 ANTENNAGATEAREA                          0.144 LAYER ME3 ;
 ANTENNADIFFAREA                          0.218 LAYER ME2 ;
 ANTENNADIFFAREA                          0.218 LAYER ME3 ;
 ANTENNAMAXAREACAR                        9.746 LAYER ME2 ;
 ANTENNAMAXAREACAR                       11.079 LAYER ME3 ;
END A2
PIN A3
  DIRECTION INPUT ;
 PORT
  LAYER ME3 ;
  RECT 277.327 0.000 277.647 0.600 ;
  LAYER ME2 ;
  RECT 277.327 0.000 277.647 0.600 ;
  LAYER ME1 ;
  RECT 277.327 0.000 277.647 0.600 ;
 END
 ANTENNAPARTIALMETALAREA                  1.188 LAYER ME2 ;
 ANTENNAGATEAREA                          0.144 LAYER ME2 ;
 ANTENNAGATEAREA                          0.144 LAYER ME3 ;
 ANTENNADIFFAREA                          0.218 LAYER ME2 ;
 ANTENNADIFFAREA                          0.218 LAYER ME3 ;
 ANTENNAMAXAREACAR                       10.582 LAYER ME2 ;
 ANTENNAMAXAREACAR                       11.915 LAYER ME3 ;
END A3
PIN A4
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 270.488 0.000 270.808 0.600 ;
  LAYER ME3 ;
  RECT 270.488 0.000 270.808 0.600 ;
  LAYER ME2 ;
  RECT 270.488 0.000 270.808 0.600 ;
  LAYER ME1 ;
  RECT 270.488 0.000 270.808 0.600 ;
 END
 ANTENNAPARTIALMETALAREA                  1.910 LAYER ME2 ;
 ANTENNAGATEAREA                          0.180 LAYER ME2 ;
 ANTENNAGATEAREA                          0.180 LAYER ME3 ;
 ANTENNAGATEAREA                          0.180 LAYER ME4 ;
 ANTENNADIFFAREA                          0.218 LAYER ME2 ;
 ANTENNADIFFAREA                          0.218 LAYER ME3 ;
 ANTENNADIFFAREA                          0.218 LAYER ME4 ;
 ANTENNAMAXAREACAR                       13.456 LAYER ME2 ;
 ANTENNAMAXAREACAR                       14.522 LAYER ME3 ;
 ANTENNAMAXAREACAR                       15.589 LAYER ME4 ;
END A4
PIN A5
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 269.868 0.000 270.188 0.600 ;
  LAYER ME3 ;
  RECT 269.868 0.000 270.188 0.600 ;
  LAYER ME2 ;
  RECT 269.868 0.000 270.188 0.600 ;
  LAYER ME1 ;
  RECT 269.868 0.000 270.188 0.600 ;
 END
 ANTENNAPARTIALMETALAREA                  1.447 LAYER ME2 ;
 ANTENNAGATEAREA                          0.180 LAYER ME2 ;
 ANTENNAGATEAREA                          0.180 LAYER ME3 ;
 ANTENNAGATEAREA                          0.180 LAYER ME4 ;
 ANTENNADIFFAREA                          0.218 LAYER ME2 ;
 ANTENNADIFFAREA                          0.218 LAYER ME3 ;
 ANTENNADIFFAREA                          0.218 LAYER ME4 ;
 ANTENNAMAXAREACAR                       12.818 LAYER ME2 ;
 ANTENNAMAXAREACAR                       13.884 LAYER ME3 ;
 ANTENNAMAXAREACAR                       14.951 LAYER ME4 ;
END A5
PIN A6
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 266.328 0.000 266.648 0.600 ;
  LAYER ME3 ;
  RECT 266.328 0.000 266.648 0.600 ;
  LAYER ME2 ;
  RECT 266.328 0.000 266.648 0.600 ;
  LAYER ME1 ;
  RECT 266.328 0.000 266.648 0.600 ;
 END
 ANTENNAPARTIALMETALAREA                  1.910 LAYER ME2 ;
 ANTENNAGATEAREA                          0.180 LAYER ME2 ;
 ANTENNAGATEAREA                          0.180 LAYER ME3 ;
 ANTENNAGATEAREA                          0.180 LAYER ME4 ;
 ANTENNADIFFAREA                          0.218 LAYER ME2 ;
 ANTENNADIFFAREA                          0.218 LAYER ME3 ;
 ANTENNADIFFAREA                          0.218 LAYER ME4 ;
 ANTENNAMAXAREACAR                       13.456 LAYER ME2 ;
 ANTENNAMAXAREACAR                       14.522 LAYER ME3 ;
 ANTENNAMAXAREACAR                       15.589 LAYER ME4 ;
END A6
PIN A7
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 265.708 0.000 266.028 0.600 ;
  LAYER ME3 ;
  RECT 265.708 0.000 266.028 0.600 ;
  LAYER ME2 ;
  RECT 265.708 0.000 266.028 0.600 ;
  LAYER ME1 ;
  RECT 265.708 0.000 266.028 0.600 ;
 END
 ANTENNAPARTIALMETALAREA                  1.447 LAYER ME2 ;
 ANTENNAGATEAREA                          0.180 LAYER ME2 ;
 ANTENNAGATEAREA                          0.180 LAYER ME3 ;
 ANTENNAGATEAREA                          0.180 LAYER ME4 ;
 ANTENNADIFFAREA                          0.218 LAYER ME2 ;
 ANTENNADIFFAREA                          0.218 LAYER ME3 ;
 ANTENNADIFFAREA                          0.218 LAYER ME4 ;
 ANTENNAMAXAREACAR                       12.818 LAYER ME2 ;
 ANTENNAMAXAREACAR                       13.884 LAYER ME3 ;
 ANTENNAMAXAREACAR                       14.951 LAYER ME4 ;
END A7
PIN A8
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 262.168 0.000 262.488 0.600 ;
  LAYER ME3 ;
  RECT 262.168 0.000 262.488 0.600 ;
  LAYER ME2 ;
  RECT 262.168 0.000 262.488 0.600 ;
  LAYER ME1 ;
  RECT 262.168 0.000 262.488 0.600 ;
 END
 ANTENNAPARTIALMETALAREA                  1.910 LAYER ME2 ;
 ANTENNAGATEAREA                          0.180 LAYER ME2 ;
 ANTENNAGATEAREA                          0.180 LAYER ME3 ;
 ANTENNAGATEAREA                          0.180 LAYER ME4 ;
 ANTENNADIFFAREA                          0.218 LAYER ME2 ;
 ANTENNADIFFAREA                          0.218 LAYER ME3 ;
 ANTENNADIFFAREA                          0.218 LAYER ME4 ;
 ANTENNAMAXAREACAR                       13.456 LAYER ME2 ;
 ANTENNAMAXAREACAR                       14.522 LAYER ME3 ;
 ANTENNAMAXAREACAR                       15.589 LAYER ME4 ;
END A8
PIN A9
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 261.548 0.000 261.868 0.600 ;
  LAYER ME3 ;
  RECT 261.548 0.000 261.868 0.600 ;
  LAYER ME2 ;
  RECT 261.548 0.000 261.868 0.600 ;
  LAYER ME1 ;
  RECT 261.548 0.000 261.868 0.600 ;
 END
 ANTENNAPARTIALMETALAREA                  1.447 LAYER ME2 ;
 ANTENNAGATEAREA                          0.180 LAYER ME2 ;
 ANTENNAGATEAREA                          0.180 LAYER ME3 ;
 ANTENNAGATEAREA                          0.180 LAYER ME4 ;
 ANTENNADIFFAREA                          0.218 LAYER ME2 ;
 ANTENNADIFFAREA                          0.218 LAYER ME3 ;
 ANTENNADIFFAREA                          0.218 LAYER ME4 ;
 ANTENNAMAXAREACAR                       12.818 LAYER ME2 ;
 ANTENNAMAXAREACAR                       13.884 LAYER ME3 ;
 ANTENNAMAXAREACAR                       14.951 LAYER ME4 ;
END A9
PIN A1
  DIRECTION INPUT ;
 PORT
  LAYER ME3 ;
  RECT 281.613 0.000 281.933 0.712 ;
  LAYER ME2 ;
  RECT 281.613 0.000 281.933 0.712 ;
  LAYER ME1 ;
  RECT 281.613 0.000 281.933 0.712 ;
 END
 ANTENNAPARTIALMETALAREA                  3.219 LAYER ME2 ;
 ANTENNAGATEAREA                          0.108 LAYER ME2 ;
 ANTENNAGATEAREA                          0.108 LAYER ME3 ;
 ANTENNADIFFAREA                          0.218 LAYER ME2 ;
 ANTENNADIFFAREA                          0.218 LAYER ME3 ;
 ANTENNAMAXAREACAR                       33.245 LAYER ME2 ;
 ANTENNAMAXAREACAR                       35.355 LAYER ME3 ;
END A1
PIN A0
  DIRECTION INPUT ;
 PORT
  LAYER ME3 ;
  RECT 284.842 0.000 285.162 0.712 ;
  LAYER ME2 ;
  RECT 284.842 0.000 285.162 0.712 ;
  LAYER ME1 ;
  RECT 284.842 0.000 285.162 0.712 ;
 END
 ANTENNAPARTIALMETALAREA                  3.457 LAYER ME2 ;
 ANTENNAGATEAREA                          0.108 LAYER ME2 ;
 ANTENNAGATEAREA                          0.108 LAYER ME3 ;
 ANTENNADIFFAREA                          0.218 LAYER ME2 ;
 ANTENNADIFFAREA                          0.218 LAYER ME3 ;
 ANTENNAMAXAREACAR                       35.986 LAYER ME2 ;
 ANTENNAMAXAREACAR                       38.095 LAYER ME3 ;
END A0
PIN DVSE
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 297.433 0.000 297.753 0.717 ;
  LAYER ME3 ;
  RECT 297.433 0.000 297.753 0.717 ;
  LAYER ME3 ;
  RECT 297.433 0.000 297.753 0.717 ;
  LAYER ME2 ;
  RECT 297.433 0.000 297.753 0.717 ;
  LAYER ME2 ;
  RECT 297.433 0.000 297.753 0.717 ;
  LAYER ME1 ;
  RECT 297.433 0.000 297.753 0.717 ;
  LAYER ME1 ;
  RECT 297.433 0.000 297.753 0.717 ;
 END
 ANTENNAPARTIALMETALAREA                  5.305 LAYER ME2 ;
 ANTENNAGATEAREA                          0.612 LAYER ME2 ;
 ANTENNAGATEAREA                          0.612 LAYER ME3 ;
 ANTENNAGATEAREA                          0.612 LAYER ME4 ;
 ANTENNADIFFAREA                          0.218 LAYER ME2 ;
 ANTENNADIFFAREA                          0.218 LAYER ME3 ;
 ANTENNADIFFAREA                          0.218 LAYER ME4 ;
 ANTENNAMAXAREACAR                       53.132 LAYER ME2 ;
 ANTENNAMAXAREACAR                       55.256 LAYER ME3 ;
 ANTENNAMAXAREACAR                       57.381 LAYER ME4 ;
END DVSE
PIN DVS3
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 296.913 0.000 297.233 0.717 ;
  LAYER ME3 ;
  RECT 296.913 0.000 297.233 0.717 ;
  LAYER ME3 ;
  RECT 296.913 0.000 297.233 0.717 ;
  LAYER ME2 ;
  RECT 296.913 0.000 297.233 0.717 ;
  LAYER ME2 ;
  RECT 296.913 0.000 297.233 0.717 ;
  LAYER ME1 ;
  RECT 296.913 0.000 297.233 0.717 ;
  LAYER ME1 ;
  RECT 296.913 0.000 297.233 0.717 ;
 END
 ANTENNAPARTIALMETALAREA                  3.675 LAYER ME2 ;
 ANTENNAGATEAREA                          0.108 LAYER ME2 ;
 ANTENNAGATEAREA                          0.108 LAYER ME3 ;
 ANTENNAGATEAREA                          0.108 LAYER ME4 ;
 ANTENNADIFFAREA                          0.218 LAYER ME2 ;
 ANTENNADIFFAREA                          0.218 LAYER ME3 ;
 ANTENNADIFFAREA                          0.218 LAYER ME4 ;
 ANTENNAMAXAREACAR                       45.625 LAYER ME2 ;
 ANTENNAMAXAREACAR                       47.749 LAYER ME3 ;
 ANTENNAMAXAREACAR                       49.874 LAYER ME4 ;
END DVS3
PIN DVS2
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 297.953 0.000 298.273 0.717 ;
  LAYER ME3 ;
  RECT 297.953 0.000 298.273 0.717 ;
  LAYER ME3 ;
  RECT 297.953 0.000 298.273 0.717 ;
  LAYER ME2 ;
  RECT 297.953 0.000 298.273 0.717 ;
  LAYER ME2 ;
  RECT 297.953 0.000 298.273 0.717 ;
  LAYER ME1 ;
  RECT 297.953 0.000 298.273 0.717 ;
  LAYER ME1 ;
  RECT 297.953 0.000 298.273 0.717 ;
 END
 ANTENNAPARTIALMETALAREA                  5.371 LAYER ME2 ;
 ANTENNAGATEAREA                          0.108 LAYER ME2 ;
 ANTENNAGATEAREA                          0.108 LAYER ME3 ;
 ANTENNAGATEAREA                          0.108 LAYER ME4 ;
 ANTENNADIFFAREA                          0.218 LAYER ME2 ;
 ANTENNADIFFAREA                          0.218 LAYER ME3 ;
 ANTENNADIFFAREA                          0.218 LAYER ME4 ;
 ANTENNAMAXAREACAR                       60.060 LAYER ME2 ;
 ANTENNAMAXAREACAR                       62.184 LAYER ME3 ;
 ANTENNAMAXAREACAR                       64.309 LAYER ME4 ;
END DVS2
PIN DVS1
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 296.393 0.000 296.713 0.717 ;
  LAYER ME3 ;
  RECT 296.393 0.000 296.713 0.717 ;
  LAYER ME3 ;
  RECT 296.393 0.000 296.713 0.717 ;
  LAYER ME2 ;
  RECT 296.393 0.000 296.713 0.717 ;
  LAYER ME2 ;
  RECT 296.393 0.000 296.713 0.717 ;
  LAYER ME1 ;
  RECT 296.393 0.000 296.713 0.717 ;
  LAYER ME1 ;
  RECT 296.393 0.000 296.713 0.717 ;
 END
 ANTENNAPARTIALMETALAREA                  3.307 LAYER ME2 ;
 ANTENNAGATEAREA                          0.108 LAYER ME2 ;
 ANTENNAGATEAREA                          0.108 LAYER ME3 ;
 ANTENNAGATEAREA                          0.108 LAYER ME4 ;
 ANTENNADIFFAREA                          0.218 LAYER ME2 ;
 ANTENNADIFFAREA                          0.218 LAYER ME3 ;
 ANTENNADIFFAREA                          0.218 LAYER ME4 ;
 ANTENNAMAXAREACAR                       42.063 LAYER ME2 ;
 ANTENNAMAXAREACAR                       44.188 LAYER ME3 ;
 ANTENNAMAXAREACAR                       46.312 LAYER ME4 ;
END DVS1
PIN DVS0
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 298.473 0.000 298.793 0.693 ;
  LAYER ME3 ;
  RECT 298.473 0.000 298.793 0.693 ;
  LAYER ME3 ;
  RECT 298.473 0.000 298.793 0.693 ;
  LAYER ME2 ;
  RECT 298.473 0.000 298.793 0.693 ;
  LAYER ME2 ;
  RECT 298.473 0.000 298.793 0.693 ;
  LAYER ME1 ;
  RECT 298.473 0.000 298.793 0.693 ;
  LAYER ME1 ;
  RECT 298.473 0.000 298.793 0.693 ;
 END
 ANTENNAPARTIALMETALAREA                  4.376 LAYER ME2 ;
 ANTENNAGATEAREA                          0.108 LAYER ME2 ;
 ANTENNAGATEAREA                          0.108 LAYER ME3 ;
 ANTENNAGATEAREA                          0.108 LAYER ME4 ;
 ANTENNADIFFAREA                          0.218 LAYER ME2 ;
 ANTENNADIFFAREA                          0.218 LAYER ME3 ;
 ANTENNADIFFAREA                          0.218 LAYER ME4 ;
 ANTENNAMAXAREACAR                       53.260 LAYER ME2 ;
 ANTENNAMAXAREACAR                       55.313 LAYER ME3 ;
 ANTENNAMAXAREACAR                       57.367 LAYER ME4 ;
END DVS0
PIN CK
  DIRECTION INPUT ;
 PORT
  LAYER ME3 ;
  RECT 289.909 0.000 290.229 0.713 ;
  LAYER ME2 ;
  RECT 289.909 0.000 290.229 0.713 ;
  LAYER ME1 ;
  RECT 289.909 0.000 290.229 0.713 ;
 END
 ANTENNAPARTIALMETALAREA                  2.392 LAYER ME2 ;
 ANTENNAPARTIALMETALAREA                  8.323 LAYER ME3 ;
 ANTENNAGATEAREA                          0.072 LAYER ME2 ;
 ANTENNAGATEAREA                          1.512 LAYER ME3 ;
 ANTENNADIFFAREA                          0.218 LAYER ME2 ;
 ANTENNADIFFAREA                          0.218 LAYER ME3 ;
 ANTENNAMAXAREACAR                       46.148 LAYER ME2 ;
 ANTENNAMAXAREACAR                      164.920 LAYER ME3 ;
END CK
PIN CSB
  DIRECTION INPUT ;
 PORT
  LAYER ME3 ;
  RECT 283.121 0.000 283.441 0.712 ;
  LAYER ME2 ;
  RECT 283.121 0.000 283.441 0.712 ;
  LAYER ME1 ;
  RECT 283.121 0.000 283.441 0.712 ;
 END
 ANTENNAPARTIALMETALAREA                  3.350 LAYER ME2 ;
 ANTENNAPARTIALMETALAREA                  8.195 LAYER ME3 ;
 ANTENNAGATEAREA                          2.244 LAYER ME2 ;
 ANTENNAGATEAREA                          3.468 LAYER ME3 ;
 ANTENNADIFFAREA                          0.218 LAYER ME2 ;
 ANTENNADIFFAREA                          0.218 LAYER ME3 ;
 ANTENNAMAXAREACAR                       17.231 LAYER ME2 ;
 ANTENNAMAXAREACAR                       56.228 LAYER ME3 ;
END CSB
PIN DI63
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 552.387 0.000 552.667 0.720 ;
  LAYER ME3 ;
  RECT 552.387 0.000 552.667 0.720 ;
  LAYER ME2 ;
  RECT 552.387 0.000 552.667 0.720 ;
  LAYER ME1 ;
  RECT 552.387 0.000 552.667 0.720 ;
 END
 ANTENNAPARTIALMETALAREA                  0.805 LAYER ME1 ;
 ANTENNAGATEAREA                          0.072 LAYER ME1 ;
 ANTENNAGATEAREA                          0.072 LAYER ME2 ;
 ANTENNAGATEAREA                          0.072 LAYER ME3 ;
 ANTENNAGATEAREA                          0.072 LAYER ME4 ;
 ANTENNADIFFAREA                          0.218 LAYER ME1 ;
 ANTENNADIFFAREA                          0.218 LAYER ME2 ;
 ANTENNADIFFAREA                          0.218 LAYER ME3 ;
 ANTENNADIFFAREA                          0.218 LAYER ME4 ;
 ANTENNAMAXAREACAR                       13.984 LAYER ME1 ;
 ANTENNAMAXAREACAR                       16.784 LAYER ME2 ;
 ANTENNAMAXAREACAR                       19.584 LAYER ME3 ;
 ANTENNAMAXAREACAR                       22.384 LAYER ME4 ;
END DI63
PIN DO63
  DIRECTION OUTPUT ;
 PORT
  LAYER ME4 ;
  RECT 550.409 0.000 550.689 0.720 ;
  LAYER ME3 ;
  RECT 550.409 0.000 550.689 0.720 ;
  LAYER ME2 ;
  RECT 550.409 0.000 550.689 0.720 ;
  LAYER ME1 ;
  RECT 550.409 0.000 550.689 0.720 ;
 END
 ANTENNAPARTIALMETALAREA                  2.030 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME3 ;
 ANTENNADIFFAREA                          1.293 LAYER ME4 ;
END DO63
PIN DI62
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 544.379 0.000 544.659 0.720 ;
  LAYER ME3 ;
  RECT 544.379 0.000 544.659 0.720 ;
  LAYER ME2 ;
  RECT 544.379 0.000 544.659 0.720 ;
  LAYER ME1 ;
  RECT 544.379 0.000 544.659 0.720 ;
 END
 ANTENNAPARTIALMETALAREA                  0.805 LAYER ME1 ;
 ANTENNAGATEAREA                          0.072 LAYER ME1 ;
 ANTENNAGATEAREA                          0.072 LAYER ME2 ;
 ANTENNAGATEAREA                          0.072 LAYER ME3 ;
 ANTENNAGATEAREA                          0.072 LAYER ME4 ;
 ANTENNADIFFAREA                          0.218 LAYER ME1 ;
 ANTENNADIFFAREA                          0.218 LAYER ME2 ;
 ANTENNADIFFAREA                          0.218 LAYER ME3 ;
 ANTENNADIFFAREA                          0.218 LAYER ME4 ;
 ANTENNAMAXAREACAR                       13.984 LAYER ME1 ;
 ANTENNAMAXAREACAR                       16.784 LAYER ME2 ;
 ANTENNAMAXAREACAR                       19.584 LAYER ME3 ;
 ANTENNAMAXAREACAR                       22.384 LAYER ME4 ;
END DI62
PIN DO62
  DIRECTION OUTPUT ;
 PORT
  LAYER ME4 ;
  RECT 542.401 0.000 542.681 0.720 ;
  LAYER ME3 ;
  RECT 542.401 0.000 542.681 0.720 ;
  LAYER ME2 ;
  RECT 542.401 0.000 542.681 0.720 ;
  LAYER ME1 ;
  RECT 542.401 0.000 542.681 0.720 ;
 END
 ANTENNAPARTIALMETALAREA                  2.030 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME3 ;
 ANTENNADIFFAREA                          1.293 LAYER ME4 ;
END DO62
PIN DI61
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 536.371 0.000 536.651 0.720 ;
  LAYER ME3 ;
  RECT 536.371 0.000 536.651 0.720 ;
  LAYER ME2 ;
  RECT 536.371 0.000 536.651 0.720 ;
  LAYER ME1 ;
  RECT 536.371 0.000 536.651 0.720 ;
 END
 ANTENNAPARTIALMETALAREA                  0.805 LAYER ME1 ;
 ANTENNAGATEAREA                          0.072 LAYER ME1 ;
 ANTENNAGATEAREA                          0.072 LAYER ME2 ;
 ANTENNAGATEAREA                          0.072 LAYER ME3 ;
 ANTENNAGATEAREA                          0.072 LAYER ME4 ;
 ANTENNADIFFAREA                          0.218 LAYER ME1 ;
 ANTENNADIFFAREA                          0.218 LAYER ME2 ;
 ANTENNADIFFAREA                          0.218 LAYER ME3 ;
 ANTENNADIFFAREA                          0.218 LAYER ME4 ;
 ANTENNAMAXAREACAR                       13.984 LAYER ME1 ;
 ANTENNAMAXAREACAR                       16.784 LAYER ME2 ;
 ANTENNAMAXAREACAR                       19.584 LAYER ME3 ;
 ANTENNAMAXAREACAR                       22.384 LAYER ME4 ;
END DI61
PIN DO61
  DIRECTION OUTPUT ;
 PORT
  LAYER ME4 ;
  RECT 534.393 0.000 534.673 0.720 ;
  LAYER ME3 ;
  RECT 534.393 0.000 534.673 0.720 ;
  LAYER ME2 ;
  RECT 534.393 0.000 534.673 0.720 ;
  LAYER ME1 ;
  RECT 534.393 0.000 534.673 0.720 ;
 END
 ANTENNAPARTIALMETALAREA                  2.030 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME3 ;
 ANTENNADIFFAREA                          1.293 LAYER ME4 ;
END DO61
PIN DI60
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 528.363 0.000 528.643 0.720 ;
  LAYER ME3 ;
  RECT 528.363 0.000 528.643 0.720 ;
  LAYER ME2 ;
  RECT 528.363 0.000 528.643 0.720 ;
  LAYER ME1 ;
  RECT 528.363 0.000 528.643 0.720 ;
 END
 ANTENNAPARTIALMETALAREA                  0.805 LAYER ME1 ;
 ANTENNAGATEAREA                          0.072 LAYER ME1 ;
 ANTENNAGATEAREA                          0.072 LAYER ME2 ;
 ANTENNAGATEAREA                          0.072 LAYER ME3 ;
 ANTENNAGATEAREA                          0.072 LAYER ME4 ;
 ANTENNADIFFAREA                          0.218 LAYER ME1 ;
 ANTENNADIFFAREA                          0.218 LAYER ME2 ;
 ANTENNADIFFAREA                          0.218 LAYER ME3 ;
 ANTENNADIFFAREA                          0.218 LAYER ME4 ;
 ANTENNAMAXAREACAR                       13.984 LAYER ME1 ;
 ANTENNAMAXAREACAR                       16.784 LAYER ME2 ;
 ANTENNAMAXAREACAR                       19.584 LAYER ME3 ;
 ANTENNAMAXAREACAR                       22.384 LAYER ME4 ;
END DI60
PIN DO60
  DIRECTION OUTPUT ;
 PORT
  LAYER ME4 ;
  RECT 526.385 0.000 526.665 0.720 ;
  LAYER ME3 ;
  RECT 526.385 0.000 526.665 0.720 ;
  LAYER ME2 ;
  RECT 526.385 0.000 526.665 0.720 ;
  LAYER ME1 ;
  RECT 526.385 0.000 526.665 0.720 ;
 END
 ANTENNAPARTIALMETALAREA                  2.030 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME3 ;
 ANTENNADIFFAREA                          1.293 LAYER ME4 ;
END DO60
PIN DI59
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 520.355 0.000 520.635 0.720 ;
  LAYER ME3 ;
  RECT 520.355 0.000 520.635 0.720 ;
  LAYER ME2 ;
  RECT 520.355 0.000 520.635 0.720 ;
  LAYER ME1 ;
  RECT 520.355 0.000 520.635 0.720 ;
 END
 ANTENNAPARTIALMETALAREA                  0.805 LAYER ME1 ;
 ANTENNAGATEAREA                          0.072 LAYER ME1 ;
 ANTENNAGATEAREA                          0.072 LAYER ME2 ;
 ANTENNAGATEAREA                          0.072 LAYER ME3 ;
 ANTENNAGATEAREA                          0.072 LAYER ME4 ;
 ANTENNADIFFAREA                          0.218 LAYER ME1 ;
 ANTENNADIFFAREA                          0.218 LAYER ME2 ;
 ANTENNADIFFAREA                          0.218 LAYER ME3 ;
 ANTENNADIFFAREA                          0.218 LAYER ME4 ;
 ANTENNAMAXAREACAR                       13.984 LAYER ME1 ;
 ANTENNAMAXAREACAR                       16.784 LAYER ME2 ;
 ANTENNAMAXAREACAR                       19.584 LAYER ME3 ;
 ANTENNAMAXAREACAR                       22.384 LAYER ME4 ;
END DI59
PIN DO59
  DIRECTION OUTPUT ;
 PORT
  LAYER ME4 ;
  RECT 518.377 0.000 518.657 0.720 ;
  LAYER ME3 ;
  RECT 518.377 0.000 518.657 0.720 ;
  LAYER ME2 ;
  RECT 518.377 0.000 518.657 0.720 ;
  LAYER ME1 ;
  RECT 518.377 0.000 518.657 0.720 ;
 END
 ANTENNAPARTIALMETALAREA                  2.030 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME3 ;
 ANTENNADIFFAREA                          1.293 LAYER ME4 ;
END DO59
PIN DI58
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 512.347 0.000 512.627 0.720 ;
  LAYER ME3 ;
  RECT 512.347 0.000 512.627 0.720 ;
  LAYER ME2 ;
  RECT 512.347 0.000 512.627 0.720 ;
  LAYER ME1 ;
  RECT 512.347 0.000 512.627 0.720 ;
 END
 ANTENNAPARTIALMETALAREA                  0.805 LAYER ME1 ;
 ANTENNAGATEAREA                          0.072 LAYER ME1 ;
 ANTENNAGATEAREA                          0.072 LAYER ME2 ;
 ANTENNAGATEAREA                          0.072 LAYER ME3 ;
 ANTENNAGATEAREA                          0.072 LAYER ME4 ;
 ANTENNADIFFAREA                          0.218 LAYER ME1 ;
 ANTENNADIFFAREA                          0.218 LAYER ME2 ;
 ANTENNADIFFAREA                          0.218 LAYER ME3 ;
 ANTENNADIFFAREA                          0.218 LAYER ME4 ;
 ANTENNAMAXAREACAR                       13.984 LAYER ME1 ;
 ANTENNAMAXAREACAR                       16.784 LAYER ME2 ;
 ANTENNAMAXAREACAR                       19.584 LAYER ME3 ;
 ANTENNAMAXAREACAR                       22.384 LAYER ME4 ;
END DI58
PIN DO58
  DIRECTION OUTPUT ;
 PORT
  LAYER ME4 ;
  RECT 510.369 0.000 510.649 0.720 ;
  LAYER ME3 ;
  RECT 510.369 0.000 510.649 0.720 ;
  LAYER ME2 ;
  RECT 510.369 0.000 510.649 0.720 ;
  LAYER ME1 ;
  RECT 510.369 0.000 510.649 0.720 ;
 END
 ANTENNAPARTIALMETALAREA                  2.030 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME3 ;
 ANTENNADIFFAREA                          1.293 LAYER ME4 ;
END DO58
PIN DI57
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 504.339 0.000 504.619 0.720 ;
  LAYER ME3 ;
  RECT 504.339 0.000 504.619 0.720 ;
  LAYER ME2 ;
  RECT 504.339 0.000 504.619 0.720 ;
  LAYER ME1 ;
  RECT 504.339 0.000 504.619 0.720 ;
 END
 ANTENNAPARTIALMETALAREA                  0.805 LAYER ME1 ;
 ANTENNAGATEAREA                          0.072 LAYER ME1 ;
 ANTENNAGATEAREA                          0.072 LAYER ME2 ;
 ANTENNAGATEAREA                          0.072 LAYER ME3 ;
 ANTENNAGATEAREA                          0.072 LAYER ME4 ;
 ANTENNADIFFAREA                          0.218 LAYER ME1 ;
 ANTENNADIFFAREA                          0.218 LAYER ME2 ;
 ANTENNADIFFAREA                          0.218 LAYER ME3 ;
 ANTENNADIFFAREA                          0.218 LAYER ME4 ;
 ANTENNAMAXAREACAR                       13.984 LAYER ME1 ;
 ANTENNAMAXAREACAR                       16.784 LAYER ME2 ;
 ANTENNAMAXAREACAR                       19.584 LAYER ME3 ;
 ANTENNAMAXAREACAR                       22.384 LAYER ME4 ;
END DI57
PIN DO57
  DIRECTION OUTPUT ;
 PORT
  LAYER ME4 ;
  RECT 502.361 0.000 502.641 0.720 ;
  LAYER ME3 ;
  RECT 502.361 0.000 502.641 0.720 ;
  LAYER ME2 ;
  RECT 502.361 0.000 502.641 0.720 ;
  LAYER ME1 ;
  RECT 502.361 0.000 502.641 0.720 ;
 END
 ANTENNAPARTIALMETALAREA                  2.030 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME3 ;
 ANTENNADIFFAREA                          1.293 LAYER ME4 ;
END DO57
PIN DI56
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 496.331 0.000 496.611 0.720 ;
  LAYER ME3 ;
  RECT 496.331 0.000 496.611 0.720 ;
  LAYER ME2 ;
  RECT 496.331 0.000 496.611 0.720 ;
  LAYER ME1 ;
  RECT 496.331 0.000 496.611 0.720 ;
 END
 ANTENNAPARTIALMETALAREA                  0.522 LAYER ME1 ;
 ANTENNAGATEAREA                          0.072 LAYER ME1 ;
 ANTENNAGATEAREA                          0.072 LAYER ME2 ;
 ANTENNAGATEAREA                          0.072 LAYER ME3 ;
 ANTENNAGATEAREA                          0.072 LAYER ME4 ;
 ANTENNADIFFAREA                          0.218 LAYER ME1 ;
 ANTENNADIFFAREA                          0.218 LAYER ME2 ;
 ANTENNADIFFAREA                          0.218 LAYER ME3 ;
 ANTENNADIFFAREA                          0.218 LAYER ME4 ;
 ANTENNAMAXAREACAR                       10.048 LAYER ME1 ;
 ANTENNAMAXAREACAR                       12.848 LAYER ME2 ;
 ANTENNAMAXAREACAR                       15.648 LAYER ME3 ;
 ANTENNAMAXAREACAR                       18.448 LAYER ME4 ;
END DI56
PIN DO56
  DIRECTION OUTPUT ;
 PORT
  LAYER ME4 ;
  RECT 494.273 0.000 494.553 0.720 ;
  LAYER ME3 ;
  RECT 494.273 0.000 494.553 0.720 ;
  LAYER ME2 ;
  RECT 494.273 0.000 494.553 0.720 ;
  LAYER ME1 ;
  RECT 494.273 0.000 494.553 0.720 ;
 END
 ANTENNAPARTIALMETALAREA                  2.030 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME3 ;
 ANTENNADIFFAREA                          1.293 LAYER ME4 ;
END DO56
PIN WEB7
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 494.753 0.000 495.033 0.720 ;
  LAYER ME3 ;
  RECT 494.753 0.000 495.033 0.720 ;
  LAYER ME2 ;
  RECT 494.753 0.000 495.033 0.720 ;
  LAYER ME1 ;
  RECT 494.753 0.000 495.033 0.720 ;
 END
 ANTENNAPARTIALMETALAREA                  0.436 LAYER ME2 ;
 ANTENNAGATEAREA                          0.288 LAYER ME2 ;
 ANTENNAGATEAREA                          0.288 LAYER ME3 ;
 ANTENNAGATEAREA                          0.288 LAYER ME4 ;
 ANTENNADIFFAREA                          0.218 LAYER ME2 ;
 ANTENNADIFFAREA                          0.218 LAYER ME3 ;
 ANTENNADIFFAREA                          0.218 LAYER ME4 ;
 ANTENNAMAXAREACAR                        4.602 LAYER ME2 ;
 ANTENNAMAXAREACAR                        5.302 LAYER ME3 ;
 ANTENNAMAXAREACAR                        6.002 LAYER ME4 ;
END WEB7
PIN DI55
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 488.323 0.000 488.603 0.720 ;
  LAYER ME3 ;
  RECT 488.323 0.000 488.603 0.720 ;
  LAYER ME2 ;
  RECT 488.323 0.000 488.603 0.720 ;
  LAYER ME1 ;
  RECT 488.323 0.000 488.603 0.720 ;
 END
 ANTENNAPARTIALMETALAREA                  0.805 LAYER ME1 ;
 ANTENNAGATEAREA                          0.072 LAYER ME1 ;
 ANTENNAGATEAREA                          0.072 LAYER ME2 ;
 ANTENNAGATEAREA                          0.072 LAYER ME3 ;
 ANTENNAGATEAREA                          0.072 LAYER ME4 ;
 ANTENNADIFFAREA                          0.218 LAYER ME1 ;
 ANTENNADIFFAREA                          0.218 LAYER ME2 ;
 ANTENNADIFFAREA                          0.218 LAYER ME3 ;
 ANTENNADIFFAREA                          0.218 LAYER ME4 ;
 ANTENNAMAXAREACAR                       13.984 LAYER ME1 ;
 ANTENNAMAXAREACAR                       16.784 LAYER ME2 ;
 ANTENNAMAXAREACAR                       19.584 LAYER ME3 ;
 ANTENNAMAXAREACAR                       22.384 LAYER ME4 ;
END DI55
PIN DO55
  DIRECTION OUTPUT ;
 PORT
  LAYER ME4 ;
  RECT 486.345 0.000 486.625 0.720 ;
  LAYER ME3 ;
  RECT 486.345 0.000 486.625 0.720 ;
  LAYER ME2 ;
  RECT 486.345 0.000 486.625 0.720 ;
  LAYER ME1 ;
  RECT 486.345 0.000 486.625 0.720 ;
 END
 ANTENNAPARTIALMETALAREA                  2.030 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME3 ;
 ANTENNADIFFAREA                          1.293 LAYER ME4 ;
END DO55
PIN DI54
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 480.315 0.000 480.595 0.720 ;
  LAYER ME3 ;
  RECT 480.315 0.000 480.595 0.720 ;
  LAYER ME2 ;
  RECT 480.315 0.000 480.595 0.720 ;
  LAYER ME1 ;
  RECT 480.315 0.000 480.595 0.720 ;
 END
 ANTENNAPARTIALMETALAREA                  0.805 LAYER ME1 ;
 ANTENNAGATEAREA                          0.072 LAYER ME1 ;
 ANTENNAGATEAREA                          0.072 LAYER ME2 ;
 ANTENNAGATEAREA                          0.072 LAYER ME3 ;
 ANTENNAGATEAREA                          0.072 LAYER ME4 ;
 ANTENNADIFFAREA                          0.218 LAYER ME1 ;
 ANTENNADIFFAREA                          0.218 LAYER ME2 ;
 ANTENNADIFFAREA                          0.218 LAYER ME3 ;
 ANTENNADIFFAREA                          0.218 LAYER ME4 ;
 ANTENNAMAXAREACAR                       13.984 LAYER ME1 ;
 ANTENNAMAXAREACAR                       16.784 LAYER ME2 ;
 ANTENNAMAXAREACAR                       19.584 LAYER ME3 ;
 ANTENNAMAXAREACAR                       22.384 LAYER ME4 ;
END DI54
PIN DO54
  DIRECTION OUTPUT ;
 PORT
  LAYER ME4 ;
  RECT 478.337 0.000 478.617 0.720 ;
  LAYER ME3 ;
  RECT 478.337 0.000 478.617 0.720 ;
  LAYER ME2 ;
  RECT 478.337 0.000 478.617 0.720 ;
  LAYER ME1 ;
  RECT 478.337 0.000 478.617 0.720 ;
 END
 ANTENNAPARTIALMETALAREA                  2.030 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME3 ;
 ANTENNADIFFAREA                          1.293 LAYER ME4 ;
END DO54
PIN DI53
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 472.307 0.000 472.587 0.720 ;
  LAYER ME3 ;
  RECT 472.307 0.000 472.587 0.720 ;
  LAYER ME2 ;
  RECT 472.307 0.000 472.587 0.720 ;
  LAYER ME1 ;
  RECT 472.307 0.000 472.587 0.720 ;
 END
 ANTENNAPARTIALMETALAREA                  0.805 LAYER ME1 ;
 ANTENNAGATEAREA                          0.072 LAYER ME1 ;
 ANTENNAGATEAREA                          0.072 LAYER ME2 ;
 ANTENNAGATEAREA                          0.072 LAYER ME3 ;
 ANTENNAGATEAREA                          0.072 LAYER ME4 ;
 ANTENNADIFFAREA                          0.218 LAYER ME1 ;
 ANTENNADIFFAREA                          0.218 LAYER ME2 ;
 ANTENNADIFFAREA                          0.218 LAYER ME3 ;
 ANTENNADIFFAREA                          0.218 LAYER ME4 ;
 ANTENNAMAXAREACAR                       13.984 LAYER ME1 ;
 ANTENNAMAXAREACAR                       16.784 LAYER ME2 ;
 ANTENNAMAXAREACAR                       19.584 LAYER ME3 ;
 ANTENNAMAXAREACAR                       22.384 LAYER ME4 ;
END DI53
PIN DO53
  DIRECTION OUTPUT ;
 PORT
  LAYER ME4 ;
  RECT 470.329 0.000 470.609 0.720 ;
  LAYER ME3 ;
  RECT 470.329 0.000 470.609 0.720 ;
  LAYER ME2 ;
  RECT 470.329 0.000 470.609 0.720 ;
  LAYER ME1 ;
  RECT 470.329 0.000 470.609 0.720 ;
 END
 ANTENNAPARTIALMETALAREA                  2.030 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME3 ;
 ANTENNADIFFAREA                          1.293 LAYER ME4 ;
END DO53
PIN DI52
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 464.299 0.000 464.579 0.720 ;
  LAYER ME3 ;
  RECT 464.299 0.000 464.579 0.720 ;
  LAYER ME2 ;
  RECT 464.299 0.000 464.579 0.720 ;
  LAYER ME1 ;
  RECT 464.299 0.000 464.579 0.720 ;
 END
 ANTENNAPARTIALMETALAREA                  0.805 LAYER ME1 ;
 ANTENNAGATEAREA                          0.072 LAYER ME1 ;
 ANTENNAGATEAREA                          0.072 LAYER ME2 ;
 ANTENNAGATEAREA                          0.072 LAYER ME3 ;
 ANTENNAGATEAREA                          0.072 LAYER ME4 ;
 ANTENNADIFFAREA                          0.218 LAYER ME1 ;
 ANTENNADIFFAREA                          0.218 LAYER ME2 ;
 ANTENNADIFFAREA                          0.218 LAYER ME3 ;
 ANTENNADIFFAREA                          0.218 LAYER ME4 ;
 ANTENNAMAXAREACAR                       13.984 LAYER ME1 ;
 ANTENNAMAXAREACAR                       16.784 LAYER ME2 ;
 ANTENNAMAXAREACAR                       19.584 LAYER ME3 ;
 ANTENNAMAXAREACAR                       22.384 LAYER ME4 ;
END DI52
PIN DO52
  DIRECTION OUTPUT ;
 PORT
  LAYER ME4 ;
  RECT 462.321 0.000 462.601 0.720 ;
  LAYER ME3 ;
  RECT 462.321 0.000 462.601 0.720 ;
  LAYER ME2 ;
  RECT 462.321 0.000 462.601 0.720 ;
  LAYER ME1 ;
  RECT 462.321 0.000 462.601 0.720 ;
 END
 ANTENNAPARTIALMETALAREA                  2.030 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME3 ;
 ANTENNADIFFAREA                          1.293 LAYER ME4 ;
END DO52
PIN DI51
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 456.291 0.000 456.571 0.720 ;
  LAYER ME3 ;
  RECT 456.291 0.000 456.571 0.720 ;
  LAYER ME2 ;
  RECT 456.291 0.000 456.571 0.720 ;
  LAYER ME1 ;
  RECT 456.291 0.000 456.571 0.720 ;
 END
 ANTENNAPARTIALMETALAREA                  0.805 LAYER ME1 ;
 ANTENNAGATEAREA                          0.072 LAYER ME1 ;
 ANTENNAGATEAREA                          0.072 LAYER ME2 ;
 ANTENNAGATEAREA                          0.072 LAYER ME3 ;
 ANTENNAGATEAREA                          0.072 LAYER ME4 ;
 ANTENNADIFFAREA                          0.218 LAYER ME1 ;
 ANTENNADIFFAREA                          0.218 LAYER ME2 ;
 ANTENNADIFFAREA                          0.218 LAYER ME3 ;
 ANTENNADIFFAREA                          0.218 LAYER ME4 ;
 ANTENNAMAXAREACAR                       13.984 LAYER ME1 ;
 ANTENNAMAXAREACAR                       16.784 LAYER ME2 ;
 ANTENNAMAXAREACAR                       19.584 LAYER ME3 ;
 ANTENNAMAXAREACAR                       22.384 LAYER ME4 ;
END DI51
PIN DO51
  DIRECTION OUTPUT ;
 PORT
  LAYER ME4 ;
  RECT 454.313 0.000 454.593 0.720 ;
  LAYER ME3 ;
  RECT 454.313 0.000 454.593 0.720 ;
  LAYER ME2 ;
  RECT 454.313 0.000 454.593 0.720 ;
  LAYER ME1 ;
  RECT 454.313 0.000 454.593 0.720 ;
 END
 ANTENNAPARTIALMETALAREA                  2.030 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME3 ;
 ANTENNADIFFAREA                          1.293 LAYER ME4 ;
END DO51
PIN DI50
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 448.283 0.000 448.563 0.720 ;
  LAYER ME3 ;
  RECT 448.283 0.000 448.563 0.720 ;
  LAYER ME2 ;
  RECT 448.283 0.000 448.563 0.720 ;
  LAYER ME1 ;
  RECT 448.283 0.000 448.563 0.720 ;
 END
 ANTENNAPARTIALMETALAREA                  0.805 LAYER ME1 ;
 ANTENNAGATEAREA                          0.072 LAYER ME1 ;
 ANTENNAGATEAREA                          0.072 LAYER ME2 ;
 ANTENNAGATEAREA                          0.072 LAYER ME3 ;
 ANTENNAGATEAREA                          0.072 LAYER ME4 ;
 ANTENNADIFFAREA                          0.218 LAYER ME1 ;
 ANTENNADIFFAREA                          0.218 LAYER ME2 ;
 ANTENNADIFFAREA                          0.218 LAYER ME3 ;
 ANTENNADIFFAREA                          0.218 LAYER ME4 ;
 ANTENNAMAXAREACAR                       13.984 LAYER ME1 ;
 ANTENNAMAXAREACAR                       16.784 LAYER ME2 ;
 ANTENNAMAXAREACAR                       19.584 LAYER ME3 ;
 ANTENNAMAXAREACAR                       22.384 LAYER ME4 ;
END DI50
PIN DO50
  DIRECTION OUTPUT ;
 PORT
  LAYER ME4 ;
  RECT 446.305 0.000 446.585 0.720 ;
  LAYER ME3 ;
  RECT 446.305 0.000 446.585 0.720 ;
  LAYER ME2 ;
  RECT 446.305 0.000 446.585 0.720 ;
  LAYER ME1 ;
  RECT 446.305 0.000 446.585 0.720 ;
 END
 ANTENNAPARTIALMETALAREA                  2.030 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME3 ;
 ANTENNADIFFAREA                          1.293 LAYER ME4 ;
END DO50
PIN DI49
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 440.275 0.000 440.555 0.720 ;
  LAYER ME3 ;
  RECT 440.275 0.000 440.555 0.720 ;
  LAYER ME2 ;
  RECT 440.275 0.000 440.555 0.720 ;
  LAYER ME1 ;
  RECT 440.275 0.000 440.555 0.720 ;
 END
 ANTENNAPARTIALMETALAREA                  0.805 LAYER ME1 ;
 ANTENNAGATEAREA                          0.072 LAYER ME1 ;
 ANTENNAGATEAREA                          0.072 LAYER ME2 ;
 ANTENNAGATEAREA                          0.072 LAYER ME3 ;
 ANTENNAGATEAREA                          0.072 LAYER ME4 ;
 ANTENNADIFFAREA                          0.218 LAYER ME1 ;
 ANTENNADIFFAREA                          0.218 LAYER ME2 ;
 ANTENNADIFFAREA                          0.218 LAYER ME3 ;
 ANTENNADIFFAREA                          0.218 LAYER ME4 ;
 ANTENNAMAXAREACAR                       13.984 LAYER ME1 ;
 ANTENNAMAXAREACAR                       16.784 LAYER ME2 ;
 ANTENNAMAXAREACAR                       19.584 LAYER ME3 ;
 ANTENNAMAXAREACAR                       22.384 LAYER ME4 ;
END DI49
PIN DO49
  DIRECTION OUTPUT ;
 PORT
  LAYER ME4 ;
  RECT 438.297 0.000 438.577 0.720 ;
  LAYER ME3 ;
  RECT 438.297 0.000 438.577 0.720 ;
  LAYER ME2 ;
  RECT 438.297 0.000 438.577 0.720 ;
  LAYER ME1 ;
  RECT 438.297 0.000 438.577 0.720 ;
 END
 ANTENNAPARTIALMETALAREA                  2.030 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME3 ;
 ANTENNADIFFAREA                          1.293 LAYER ME4 ;
END DO49
PIN DI48
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 432.267 0.000 432.547 0.720 ;
  LAYER ME3 ;
  RECT 432.267 0.000 432.547 0.720 ;
  LAYER ME2 ;
  RECT 432.267 0.000 432.547 0.720 ;
  LAYER ME1 ;
  RECT 432.267 0.000 432.547 0.720 ;
 END
 ANTENNAPARTIALMETALAREA                  0.522 LAYER ME1 ;
 ANTENNAGATEAREA                          0.072 LAYER ME1 ;
 ANTENNAGATEAREA                          0.072 LAYER ME2 ;
 ANTENNAGATEAREA                          0.072 LAYER ME3 ;
 ANTENNAGATEAREA                          0.072 LAYER ME4 ;
 ANTENNADIFFAREA                          0.218 LAYER ME1 ;
 ANTENNADIFFAREA                          0.218 LAYER ME2 ;
 ANTENNADIFFAREA                          0.218 LAYER ME3 ;
 ANTENNADIFFAREA                          0.218 LAYER ME4 ;
 ANTENNAMAXAREACAR                       10.048 LAYER ME1 ;
 ANTENNAMAXAREACAR                       12.848 LAYER ME2 ;
 ANTENNAMAXAREACAR                       15.648 LAYER ME3 ;
 ANTENNAMAXAREACAR                       18.448 LAYER ME4 ;
END DI48
PIN DO48
  DIRECTION OUTPUT ;
 PORT
  LAYER ME4 ;
  RECT 430.209 0.000 430.489 0.720 ;
  LAYER ME3 ;
  RECT 430.209 0.000 430.489 0.720 ;
  LAYER ME2 ;
  RECT 430.209 0.000 430.489 0.720 ;
  LAYER ME1 ;
  RECT 430.209 0.000 430.489 0.720 ;
 END
 ANTENNAPARTIALMETALAREA                  2.030 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME3 ;
 ANTENNADIFFAREA                          1.293 LAYER ME4 ;
END DO48
PIN WEB6
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 430.689 0.000 430.969 0.720 ;
  LAYER ME3 ;
  RECT 430.689 0.000 430.969 0.720 ;
  LAYER ME2 ;
  RECT 430.689 0.000 430.969 0.720 ;
  LAYER ME1 ;
  RECT 430.689 0.000 430.969 0.720 ;
 END
 ANTENNAPARTIALMETALAREA                  0.436 LAYER ME2 ;
 ANTENNAGATEAREA                          0.288 LAYER ME2 ;
 ANTENNAGATEAREA                          0.288 LAYER ME3 ;
 ANTENNAGATEAREA                          0.288 LAYER ME4 ;
 ANTENNADIFFAREA                          0.218 LAYER ME2 ;
 ANTENNADIFFAREA                          0.218 LAYER ME3 ;
 ANTENNADIFFAREA                          0.218 LAYER ME4 ;
 ANTENNAMAXAREACAR                        4.602 LAYER ME2 ;
 ANTENNAMAXAREACAR                        5.302 LAYER ME3 ;
 ANTENNAMAXAREACAR                        6.002 LAYER ME4 ;
END WEB6
PIN DI47
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 424.259 0.000 424.539 0.720 ;
  LAYER ME3 ;
  RECT 424.259 0.000 424.539 0.720 ;
  LAYER ME2 ;
  RECT 424.259 0.000 424.539 0.720 ;
  LAYER ME1 ;
  RECT 424.259 0.000 424.539 0.720 ;
 END
 ANTENNAPARTIALMETALAREA                  0.805 LAYER ME1 ;
 ANTENNAGATEAREA                          0.072 LAYER ME1 ;
 ANTENNAGATEAREA                          0.072 LAYER ME2 ;
 ANTENNAGATEAREA                          0.072 LAYER ME3 ;
 ANTENNAGATEAREA                          0.072 LAYER ME4 ;
 ANTENNADIFFAREA                          0.218 LAYER ME1 ;
 ANTENNADIFFAREA                          0.218 LAYER ME2 ;
 ANTENNADIFFAREA                          0.218 LAYER ME3 ;
 ANTENNADIFFAREA                          0.218 LAYER ME4 ;
 ANTENNAMAXAREACAR                       13.984 LAYER ME1 ;
 ANTENNAMAXAREACAR                       16.784 LAYER ME2 ;
 ANTENNAMAXAREACAR                       19.584 LAYER ME3 ;
 ANTENNAMAXAREACAR                       22.384 LAYER ME4 ;
END DI47
PIN DO47
  DIRECTION OUTPUT ;
 PORT
  LAYER ME4 ;
  RECT 422.281 0.000 422.561 0.720 ;
  LAYER ME3 ;
  RECT 422.281 0.000 422.561 0.720 ;
  LAYER ME2 ;
  RECT 422.281 0.000 422.561 0.720 ;
  LAYER ME1 ;
  RECT 422.281 0.000 422.561 0.720 ;
 END
 ANTENNAPARTIALMETALAREA                  2.030 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME3 ;
 ANTENNADIFFAREA                          1.293 LAYER ME4 ;
END DO47
PIN DI46
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 416.251 0.000 416.531 0.720 ;
  LAYER ME3 ;
  RECT 416.251 0.000 416.531 0.720 ;
  LAYER ME2 ;
  RECT 416.251 0.000 416.531 0.720 ;
  LAYER ME1 ;
  RECT 416.251 0.000 416.531 0.720 ;
 END
 ANTENNAPARTIALMETALAREA                  0.805 LAYER ME1 ;
 ANTENNAGATEAREA                          0.072 LAYER ME1 ;
 ANTENNAGATEAREA                          0.072 LAYER ME2 ;
 ANTENNAGATEAREA                          0.072 LAYER ME3 ;
 ANTENNAGATEAREA                          0.072 LAYER ME4 ;
 ANTENNADIFFAREA                          0.218 LAYER ME1 ;
 ANTENNADIFFAREA                          0.218 LAYER ME2 ;
 ANTENNADIFFAREA                          0.218 LAYER ME3 ;
 ANTENNADIFFAREA                          0.218 LAYER ME4 ;
 ANTENNAMAXAREACAR                       13.984 LAYER ME1 ;
 ANTENNAMAXAREACAR                       16.784 LAYER ME2 ;
 ANTENNAMAXAREACAR                       19.584 LAYER ME3 ;
 ANTENNAMAXAREACAR                       22.384 LAYER ME4 ;
END DI46
PIN DO46
  DIRECTION OUTPUT ;
 PORT
  LAYER ME4 ;
  RECT 414.273 0.000 414.553 0.720 ;
  LAYER ME3 ;
  RECT 414.273 0.000 414.553 0.720 ;
  LAYER ME2 ;
  RECT 414.273 0.000 414.553 0.720 ;
  LAYER ME1 ;
  RECT 414.273 0.000 414.553 0.720 ;
 END
 ANTENNAPARTIALMETALAREA                  2.030 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME3 ;
 ANTENNADIFFAREA                          1.293 LAYER ME4 ;
END DO46
PIN DI45
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 408.243 0.000 408.523 0.720 ;
  LAYER ME3 ;
  RECT 408.243 0.000 408.523 0.720 ;
  LAYER ME2 ;
  RECT 408.243 0.000 408.523 0.720 ;
  LAYER ME1 ;
  RECT 408.243 0.000 408.523 0.720 ;
 END
 ANTENNAPARTIALMETALAREA                  0.805 LAYER ME1 ;
 ANTENNAGATEAREA                          0.072 LAYER ME1 ;
 ANTENNAGATEAREA                          0.072 LAYER ME2 ;
 ANTENNAGATEAREA                          0.072 LAYER ME3 ;
 ANTENNAGATEAREA                          0.072 LAYER ME4 ;
 ANTENNADIFFAREA                          0.218 LAYER ME1 ;
 ANTENNADIFFAREA                          0.218 LAYER ME2 ;
 ANTENNADIFFAREA                          0.218 LAYER ME3 ;
 ANTENNADIFFAREA                          0.218 LAYER ME4 ;
 ANTENNAMAXAREACAR                       13.984 LAYER ME1 ;
 ANTENNAMAXAREACAR                       16.784 LAYER ME2 ;
 ANTENNAMAXAREACAR                       19.584 LAYER ME3 ;
 ANTENNAMAXAREACAR                       22.384 LAYER ME4 ;
END DI45
PIN DO45
  DIRECTION OUTPUT ;
 PORT
  LAYER ME4 ;
  RECT 406.265 0.000 406.545 0.720 ;
  LAYER ME3 ;
  RECT 406.265 0.000 406.545 0.720 ;
  LAYER ME2 ;
  RECT 406.265 0.000 406.545 0.720 ;
  LAYER ME1 ;
  RECT 406.265 0.000 406.545 0.720 ;
 END
 ANTENNAPARTIALMETALAREA                  2.030 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME3 ;
 ANTENNADIFFAREA                          1.293 LAYER ME4 ;
END DO45
PIN DI44
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 400.235 0.000 400.515 0.720 ;
  LAYER ME3 ;
  RECT 400.235 0.000 400.515 0.720 ;
  LAYER ME2 ;
  RECT 400.235 0.000 400.515 0.720 ;
  LAYER ME1 ;
  RECT 400.235 0.000 400.515 0.720 ;
 END
 ANTENNAPARTIALMETALAREA                  0.805 LAYER ME1 ;
 ANTENNAGATEAREA                          0.072 LAYER ME1 ;
 ANTENNAGATEAREA                          0.072 LAYER ME2 ;
 ANTENNAGATEAREA                          0.072 LAYER ME3 ;
 ANTENNAGATEAREA                          0.072 LAYER ME4 ;
 ANTENNADIFFAREA                          0.218 LAYER ME1 ;
 ANTENNADIFFAREA                          0.218 LAYER ME2 ;
 ANTENNADIFFAREA                          0.218 LAYER ME3 ;
 ANTENNADIFFAREA                          0.218 LAYER ME4 ;
 ANTENNAMAXAREACAR                       13.984 LAYER ME1 ;
 ANTENNAMAXAREACAR                       16.784 LAYER ME2 ;
 ANTENNAMAXAREACAR                       19.584 LAYER ME3 ;
 ANTENNAMAXAREACAR                       22.384 LAYER ME4 ;
END DI44
PIN DO44
  DIRECTION OUTPUT ;
 PORT
  LAYER ME4 ;
  RECT 398.257 0.000 398.537 0.720 ;
  LAYER ME3 ;
  RECT 398.257 0.000 398.537 0.720 ;
  LAYER ME2 ;
  RECT 398.257 0.000 398.537 0.720 ;
  LAYER ME1 ;
  RECT 398.257 0.000 398.537 0.720 ;
 END
 ANTENNAPARTIALMETALAREA                  2.030 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME3 ;
 ANTENNADIFFAREA                          1.293 LAYER ME4 ;
END DO44
PIN DI43
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 392.227 0.000 392.507 0.720 ;
  LAYER ME3 ;
  RECT 392.227 0.000 392.507 0.720 ;
  LAYER ME2 ;
  RECT 392.227 0.000 392.507 0.720 ;
  LAYER ME1 ;
  RECT 392.227 0.000 392.507 0.720 ;
 END
 ANTENNAPARTIALMETALAREA                  0.805 LAYER ME1 ;
 ANTENNAGATEAREA                          0.072 LAYER ME1 ;
 ANTENNAGATEAREA                          0.072 LAYER ME2 ;
 ANTENNAGATEAREA                          0.072 LAYER ME3 ;
 ANTENNAGATEAREA                          0.072 LAYER ME4 ;
 ANTENNADIFFAREA                          0.218 LAYER ME1 ;
 ANTENNADIFFAREA                          0.218 LAYER ME2 ;
 ANTENNADIFFAREA                          0.218 LAYER ME3 ;
 ANTENNADIFFAREA                          0.218 LAYER ME4 ;
 ANTENNAMAXAREACAR                       13.984 LAYER ME1 ;
 ANTENNAMAXAREACAR                       16.784 LAYER ME2 ;
 ANTENNAMAXAREACAR                       19.584 LAYER ME3 ;
 ANTENNAMAXAREACAR                       22.384 LAYER ME4 ;
END DI43
PIN DO43
  DIRECTION OUTPUT ;
 PORT
  LAYER ME4 ;
  RECT 390.249 0.000 390.529 0.720 ;
  LAYER ME3 ;
  RECT 390.249 0.000 390.529 0.720 ;
  LAYER ME2 ;
  RECT 390.249 0.000 390.529 0.720 ;
  LAYER ME1 ;
  RECT 390.249 0.000 390.529 0.720 ;
 END
 ANTENNAPARTIALMETALAREA                  2.030 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME3 ;
 ANTENNADIFFAREA                          1.293 LAYER ME4 ;
END DO43
PIN DI42
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 384.219 0.000 384.499 0.720 ;
  LAYER ME3 ;
  RECT 384.219 0.000 384.499 0.720 ;
  LAYER ME2 ;
  RECT 384.219 0.000 384.499 0.720 ;
  LAYER ME1 ;
  RECT 384.219 0.000 384.499 0.720 ;
 END
 ANTENNAPARTIALMETALAREA                  0.805 LAYER ME1 ;
 ANTENNAGATEAREA                          0.072 LAYER ME1 ;
 ANTENNAGATEAREA                          0.072 LAYER ME2 ;
 ANTENNAGATEAREA                          0.072 LAYER ME3 ;
 ANTENNAGATEAREA                          0.072 LAYER ME4 ;
 ANTENNADIFFAREA                          0.218 LAYER ME1 ;
 ANTENNADIFFAREA                          0.218 LAYER ME2 ;
 ANTENNADIFFAREA                          0.218 LAYER ME3 ;
 ANTENNADIFFAREA                          0.218 LAYER ME4 ;
 ANTENNAMAXAREACAR                       13.984 LAYER ME1 ;
 ANTENNAMAXAREACAR                       16.784 LAYER ME2 ;
 ANTENNAMAXAREACAR                       19.584 LAYER ME3 ;
 ANTENNAMAXAREACAR                       22.384 LAYER ME4 ;
END DI42
PIN DO42
  DIRECTION OUTPUT ;
 PORT
  LAYER ME4 ;
  RECT 382.241 0.000 382.521 0.720 ;
  LAYER ME3 ;
  RECT 382.241 0.000 382.521 0.720 ;
  LAYER ME2 ;
  RECT 382.241 0.000 382.521 0.720 ;
  LAYER ME1 ;
  RECT 382.241 0.000 382.521 0.720 ;
 END
 ANTENNAPARTIALMETALAREA                  2.030 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME3 ;
 ANTENNADIFFAREA                          1.293 LAYER ME4 ;
END DO42
PIN DI41
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 376.211 0.000 376.491 0.720 ;
  LAYER ME3 ;
  RECT 376.211 0.000 376.491 0.720 ;
  LAYER ME2 ;
  RECT 376.211 0.000 376.491 0.720 ;
  LAYER ME1 ;
  RECT 376.211 0.000 376.491 0.720 ;
 END
 ANTENNAPARTIALMETALAREA                  0.805 LAYER ME1 ;
 ANTENNAGATEAREA                          0.072 LAYER ME1 ;
 ANTENNAGATEAREA                          0.072 LAYER ME2 ;
 ANTENNAGATEAREA                          0.072 LAYER ME3 ;
 ANTENNAGATEAREA                          0.072 LAYER ME4 ;
 ANTENNADIFFAREA                          0.218 LAYER ME1 ;
 ANTENNADIFFAREA                          0.218 LAYER ME2 ;
 ANTENNADIFFAREA                          0.218 LAYER ME3 ;
 ANTENNADIFFAREA                          0.218 LAYER ME4 ;
 ANTENNAMAXAREACAR                       13.984 LAYER ME1 ;
 ANTENNAMAXAREACAR                       16.784 LAYER ME2 ;
 ANTENNAMAXAREACAR                       19.584 LAYER ME3 ;
 ANTENNAMAXAREACAR                       22.384 LAYER ME4 ;
END DI41
PIN DO41
  DIRECTION OUTPUT ;
 PORT
  LAYER ME4 ;
  RECT 374.233 0.000 374.513 0.720 ;
  LAYER ME3 ;
  RECT 374.233 0.000 374.513 0.720 ;
  LAYER ME2 ;
  RECT 374.233 0.000 374.513 0.720 ;
  LAYER ME1 ;
  RECT 374.233 0.000 374.513 0.720 ;
 END
 ANTENNAPARTIALMETALAREA                  2.030 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME3 ;
 ANTENNADIFFAREA                          1.293 LAYER ME4 ;
END DO41
PIN DI40
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 368.203 0.000 368.483 0.720 ;
  LAYER ME3 ;
  RECT 368.203 0.000 368.483 0.720 ;
  LAYER ME2 ;
  RECT 368.203 0.000 368.483 0.720 ;
  LAYER ME1 ;
  RECT 368.203 0.000 368.483 0.720 ;
 END
 ANTENNAPARTIALMETALAREA                  0.522 LAYER ME1 ;
 ANTENNAGATEAREA                          0.072 LAYER ME1 ;
 ANTENNAGATEAREA                          0.072 LAYER ME2 ;
 ANTENNAGATEAREA                          0.072 LAYER ME3 ;
 ANTENNAGATEAREA                          0.072 LAYER ME4 ;
 ANTENNADIFFAREA                          0.218 LAYER ME1 ;
 ANTENNADIFFAREA                          0.218 LAYER ME2 ;
 ANTENNADIFFAREA                          0.218 LAYER ME3 ;
 ANTENNADIFFAREA                          0.218 LAYER ME4 ;
 ANTENNAMAXAREACAR                       10.048 LAYER ME1 ;
 ANTENNAMAXAREACAR                       12.848 LAYER ME2 ;
 ANTENNAMAXAREACAR                       15.648 LAYER ME3 ;
 ANTENNAMAXAREACAR                       18.448 LAYER ME4 ;
END DI40
PIN DO40
  DIRECTION OUTPUT ;
 PORT
  LAYER ME4 ;
  RECT 366.145 0.000 366.425 0.720 ;
  LAYER ME3 ;
  RECT 366.145 0.000 366.425 0.720 ;
  LAYER ME2 ;
  RECT 366.145 0.000 366.425 0.720 ;
  LAYER ME1 ;
  RECT 366.145 0.000 366.425 0.720 ;
 END
 ANTENNAPARTIALMETALAREA                  2.030 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME3 ;
 ANTENNADIFFAREA                          1.293 LAYER ME4 ;
END DO40
PIN WEB5
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 366.625 0.000 366.905 0.720 ;
  LAYER ME3 ;
  RECT 366.625 0.000 366.905 0.720 ;
  LAYER ME2 ;
  RECT 366.625 0.000 366.905 0.720 ;
  LAYER ME1 ;
  RECT 366.625 0.000 366.905 0.720 ;
 END
 ANTENNAPARTIALMETALAREA                  0.436 LAYER ME2 ;
 ANTENNAGATEAREA                          0.288 LAYER ME2 ;
 ANTENNAGATEAREA                          0.288 LAYER ME3 ;
 ANTENNAGATEAREA                          0.288 LAYER ME4 ;
 ANTENNADIFFAREA                          0.218 LAYER ME2 ;
 ANTENNADIFFAREA                          0.218 LAYER ME3 ;
 ANTENNADIFFAREA                          0.218 LAYER ME4 ;
 ANTENNAMAXAREACAR                        4.602 LAYER ME2 ;
 ANTENNAMAXAREACAR                        5.302 LAYER ME3 ;
 ANTENNAMAXAREACAR                        6.002 LAYER ME4 ;
END WEB5
PIN DI39
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 360.195 0.000 360.475 0.720 ;
  LAYER ME3 ;
  RECT 360.195 0.000 360.475 0.720 ;
  LAYER ME2 ;
  RECT 360.195 0.000 360.475 0.720 ;
  LAYER ME1 ;
  RECT 360.195 0.000 360.475 0.720 ;
 END
 ANTENNAPARTIALMETALAREA                  0.805 LAYER ME1 ;
 ANTENNAGATEAREA                          0.072 LAYER ME1 ;
 ANTENNAGATEAREA                          0.072 LAYER ME2 ;
 ANTENNAGATEAREA                          0.072 LAYER ME3 ;
 ANTENNAGATEAREA                          0.072 LAYER ME4 ;
 ANTENNADIFFAREA                          0.218 LAYER ME1 ;
 ANTENNADIFFAREA                          0.218 LAYER ME2 ;
 ANTENNADIFFAREA                          0.218 LAYER ME3 ;
 ANTENNADIFFAREA                          0.218 LAYER ME4 ;
 ANTENNAMAXAREACAR                       13.984 LAYER ME1 ;
 ANTENNAMAXAREACAR                       16.784 LAYER ME2 ;
 ANTENNAMAXAREACAR                       19.584 LAYER ME3 ;
 ANTENNAMAXAREACAR                       22.384 LAYER ME4 ;
END DI39
PIN DO39
  DIRECTION OUTPUT ;
 PORT
  LAYER ME4 ;
  RECT 358.217 0.000 358.497 0.720 ;
  LAYER ME3 ;
  RECT 358.217 0.000 358.497 0.720 ;
  LAYER ME2 ;
  RECT 358.217 0.000 358.497 0.720 ;
  LAYER ME1 ;
  RECT 358.217 0.000 358.497 0.720 ;
 END
 ANTENNAPARTIALMETALAREA                  2.030 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME3 ;
 ANTENNADIFFAREA                          1.293 LAYER ME4 ;
END DO39
PIN DI38
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 352.187 0.000 352.467 0.720 ;
  LAYER ME3 ;
  RECT 352.187 0.000 352.467 0.720 ;
  LAYER ME2 ;
  RECT 352.187 0.000 352.467 0.720 ;
  LAYER ME1 ;
  RECT 352.187 0.000 352.467 0.720 ;
 END
 ANTENNAPARTIALMETALAREA                  0.805 LAYER ME1 ;
 ANTENNAGATEAREA                          0.072 LAYER ME1 ;
 ANTENNAGATEAREA                          0.072 LAYER ME2 ;
 ANTENNAGATEAREA                          0.072 LAYER ME3 ;
 ANTENNAGATEAREA                          0.072 LAYER ME4 ;
 ANTENNADIFFAREA                          0.218 LAYER ME1 ;
 ANTENNADIFFAREA                          0.218 LAYER ME2 ;
 ANTENNADIFFAREA                          0.218 LAYER ME3 ;
 ANTENNADIFFAREA                          0.218 LAYER ME4 ;
 ANTENNAMAXAREACAR                       13.984 LAYER ME1 ;
 ANTENNAMAXAREACAR                       16.784 LAYER ME2 ;
 ANTENNAMAXAREACAR                       19.584 LAYER ME3 ;
 ANTENNAMAXAREACAR                       22.384 LAYER ME4 ;
END DI38
PIN DO38
  DIRECTION OUTPUT ;
 PORT
  LAYER ME4 ;
  RECT 350.209 0.000 350.489 0.720 ;
  LAYER ME3 ;
  RECT 350.209 0.000 350.489 0.720 ;
  LAYER ME2 ;
  RECT 350.209 0.000 350.489 0.720 ;
  LAYER ME1 ;
  RECT 350.209 0.000 350.489 0.720 ;
 END
 ANTENNAPARTIALMETALAREA                  2.030 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME3 ;
 ANTENNADIFFAREA                          1.293 LAYER ME4 ;
END DO38
PIN DI37
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 344.179 0.000 344.459 0.720 ;
  LAYER ME3 ;
  RECT 344.179 0.000 344.459 0.720 ;
  LAYER ME2 ;
  RECT 344.179 0.000 344.459 0.720 ;
  LAYER ME1 ;
  RECT 344.179 0.000 344.459 0.720 ;
 END
 ANTENNAPARTIALMETALAREA                  0.805 LAYER ME1 ;
 ANTENNAGATEAREA                          0.072 LAYER ME1 ;
 ANTENNAGATEAREA                          0.072 LAYER ME2 ;
 ANTENNAGATEAREA                          0.072 LAYER ME3 ;
 ANTENNAGATEAREA                          0.072 LAYER ME4 ;
 ANTENNADIFFAREA                          0.218 LAYER ME1 ;
 ANTENNADIFFAREA                          0.218 LAYER ME2 ;
 ANTENNADIFFAREA                          0.218 LAYER ME3 ;
 ANTENNADIFFAREA                          0.218 LAYER ME4 ;
 ANTENNAMAXAREACAR                       13.984 LAYER ME1 ;
 ANTENNAMAXAREACAR                       16.784 LAYER ME2 ;
 ANTENNAMAXAREACAR                       19.584 LAYER ME3 ;
 ANTENNAMAXAREACAR                       22.384 LAYER ME4 ;
END DI37
PIN DO37
  DIRECTION OUTPUT ;
 PORT
  LAYER ME4 ;
  RECT 342.201 0.000 342.481 0.720 ;
  LAYER ME3 ;
  RECT 342.201 0.000 342.481 0.720 ;
  LAYER ME2 ;
  RECT 342.201 0.000 342.481 0.720 ;
  LAYER ME1 ;
  RECT 342.201 0.000 342.481 0.720 ;
 END
 ANTENNAPARTIALMETALAREA                  2.030 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME3 ;
 ANTENNADIFFAREA                          1.293 LAYER ME4 ;
END DO37
PIN DI36
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 336.171 0.000 336.451 0.720 ;
  LAYER ME3 ;
  RECT 336.171 0.000 336.451 0.720 ;
  LAYER ME2 ;
  RECT 336.171 0.000 336.451 0.720 ;
  LAYER ME1 ;
  RECT 336.171 0.000 336.451 0.720 ;
 END
 ANTENNAPARTIALMETALAREA                  0.805 LAYER ME1 ;
 ANTENNAGATEAREA                          0.072 LAYER ME1 ;
 ANTENNAGATEAREA                          0.072 LAYER ME2 ;
 ANTENNAGATEAREA                          0.072 LAYER ME3 ;
 ANTENNAGATEAREA                          0.072 LAYER ME4 ;
 ANTENNADIFFAREA                          0.218 LAYER ME1 ;
 ANTENNADIFFAREA                          0.218 LAYER ME2 ;
 ANTENNADIFFAREA                          0.218 LAYER ME3 ;
 ANTENNADIFFAREA                          0.218 LAYER ME4 ;
 ANTENNAMAXAREACAR                       13.984 LAYER ME1 ;
 ANTENNAMAXAREACAR                       16.784 LAYER ME2 ;
 ANTENNAMAXAREACAR                       19.584 LAYER ME3 ;
 ANTENNAMAXAREACAR                       22.384 LAYER ME4 ;
END DI36
PIN DO36
  DIRECTION OUTPUT ;
 PORT
  LAYER ME4 ;
  RECT 334.193 0.000 334.473 0.720 ;
  LAYER ME3 ;
  RECT 334.193 0.000 334.473 0.720 ;
  LAYER ME2 ;
  RECT 334.193 0.000 334.473 0.720 ;
  LAYER ME1 ;
  RECT 334.193 0.000 334.473 0.720 ;
 END
 ANTENNAPARTIALMETALAREA                  2.030 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME3 ;
 ANTENNADIFFAREA                          1.293 LAYER ME4 ;
END DO36
PIN DI35
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 328.163 0.000 328.443 0.720 ;
  LAYER ME3 ;
  RECT 328.163 0.000 328.443 0.720 ;
  LAYER ME2 ;
  RECT 328.163 0.000 328.443 0.720 ;
  LAYER ME1 ;
  RECT 328.163 0.000 328.443 0.720 ;
 END
 ANTENNAPARTIALMETALAREA                  0.805 LAYER ME1 ;
 ANTENNAGATEAREA                          0.072 LAYER ME1 ;
 ANTENNAGATEAREA                          0.072 LAYER ME2 ;
 ANTENNAGATEAREA                          0.072 LAYER ME3 ;
 ANTENNAGATEAREA                          0.072 LAYER ME4 ;
 ANTENNADIFFAREA                          0.218 LAYER ME1 ;
 ANTENNADIFFAREA                          0.218 LAYER ME2 ;
 ANTENNADIFFAREA                          0.218 LAYER ME3 ;
 ANTENNADIFFAREA                          0.218 LAYER ME4 ;
 ANTENNAMAXAREACAR                       13.984 LAYER ME1 ;
 ANTENNAMAXAREACAR                       16.784 LAYER ME2 ;
 ANTENNAMAXAREACAR                       19.584 LAYER ME3 ;
 ANTENNAMAXAREACAR                       22.384 LAYER ME4 ;
END DI35
PIN DO35
  DIRECTION OUTPUT ;
 PORT
  LAYER ME4 ;
  RECT 326.185 0.000 326.465 0.720 ;
  LAYER ME3 ;
  RECT 326.185 0.000 326.465 0.720 ;
  LAYER ME2 ;
  RECT 326.185 0.000 326.465 0.720 ;
  LAYER ME1 ;
  RECT 326.185 0.000 326.465 0.720 ;
 END
 ANTENNAPARTIALMETALAREA                  2.030 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME3 ;
 ANTENNADIFFAREA                          1.293 LAYER ME4 ;
END DO35
PIN DI34
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 320.155 0.000 320.435 0.720 ;
  LAYER ME3 ;
  RECT 320.155 0.000 320.435 0.720 ;
  LAYER ME2 ;
  RECT 320.155 0.000 320.435 0.720 ;
  LAYER ME1 ;
  RECT 320.155 0.000 320.435 0.720 ;
 END
 ANTENNAPARTIALMETALAREA                  0.805 LAYER ME1 ;
 ANTENNAGATEAREA                          0.072 LAYER ME1 ;
 ANTENNAGATEAREA                          0.072 LAYER ME2 ;
 ANTENNAGATEAREA                          0.072 LAYER ME3 ;
 ANTENNAGATEAREA                          0.072 LAYER ME4 ;
 ANTENNADIFFAREA                          0.218 LAYER ME1 ;
 ANTENNADIFFAREA                          0.218 LAYER ME2 ;
 ANTENNADIFFAREA                          0.218 LAYER ME3 ;
 ANTENNADIFFAREA                          0.218 LAYER ME4 ;
 ANTENNAMAXAREACAR                       13.984 LAYER ME1 ;
 ANTENNAMAXAREACAR                       16.784 LAYER ME2 ;
 ANTENNAMAXAREACAR                       19.584 LAYER ME3 ;
 ANTENNAMAXAREACAR                       22.384 LAYER ME4 ;
END DI34
PIN DO34
  DIRECTION OUTPUT ;
 PORT
  LAYER ME4 ;
  RECT 318.177 0.000 318.457 0.720 ;
  LAYER ME3 ;
  RECT 318.177 0.000 318.457 0.720 ;
  LAYER ME2 ;
  RECT 318.177 0.000 318.457 0.720 ;
  LAYER ME1 ;
  RECT 318.177 0.000 318.457 0.720 ;
 END
 ANTENNAPARTIALMETALAREA                  2.030 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME3 ;
 ANTENNADIFFAREA                          1.293 LAYER ME4 ;
END DO34
PIN DI33
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 312.147 0.000 312.427 0.720 ;
  LAYER ME3 ;
  RECT 312.147 0.000 312.427 0.720 ;
  LAYER ME2 ;
  RECT 312.147 0.000 312.427 0.720 ;
  LAYER ME1 ;
  RECT 312.147 0.000 312.427 0.720 ;
 END
 ANTENNAPARTIALMETALAREA                  0.805 LAYER ME1 ;
 ANTENNAGATEAREA                          0.072 LAYER ME1 ;
 ANTENNAGATEAREA                          0.072 LAYER ME2 ;
 ANTENNAGATEAREA                          0.072 LAYER ME3 ;
 ANTENNAGATEAREA                          0.072 LAYER ME4 ;
 ANTENNADIFFAREA                          0.218 LAYER ME1 ;
 ANTENNADIFFAREA                          0.218 LAYER ME2 ;
 ANTENNADIFFAREA                          0.218 LAYER ME3 ;
 ANTENNADIFFAREA                          0.218 LAYER ME4 ;
 ANTENNAMAXAREACAR                       13.984 LAYER ME1 ;
 ANTENNAMAXAREACAR                       16.784 LAYER ME2 ;
 ANTENNAMAXAREACAR                       19.584 LAYER ME3 ;
 ANTENNAMAXAREACAR                       22.384 LAYER ME4 ;
END DI33
PIN DO33
  DIRECTION OUTPUT ;
 PORT
  LAYER ME4 ;
  RECT 310.169 0.000 310.449 0.720 ;
  LAYER ME3 ;
  RECT 310.169 0.000 310.449 0.720 ;
  LAYER ME2 ;
  RECT 310.169 0.000 310.449 0.720 ;
  LAYER ME1 ;
  RECT 310.169 0.000 310.449 0.720 ;
 END
 ANTENNAPARTIALMETALAREA                  2.030 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME3 ;
 ANTENNADIFFAREA                          1.293 LAYER ME4 ;
END DO33
PIN DI32
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 304.139 0.000 304.419 0.720 ;
  LAYER ME3 ;
  RECT 304.139 0.000 304.419 0.720 ;
  LAYER ME2 ;
  RECT 304.139 0.000 304.419 0.720 ;
  LAYER ME1 ;
  RECT 304.139 0.000 304.419 0.720 ;
 END
 ANTENNAPARTIALMETALAREA                  0.522 LAYER ME1 ;
 ANTENNAGATEAREA                          0.072 LAYER ME1 ;
 ANTENNAGATEAREA                          0.072 LAYER ME2 ;
 ANTENNAGATEAREA                          0.072 LAYER ME3 ;
 ANTENNAGATEAREA                          0.072 LAYER ME4 ;
 ANTENNADIFFAREA                          0.218 LAYER ME1 ;
 ANTENNADIFFAREA                          0.218 LAYER ME2 ;
 ANTENNADIFFAREA                          0.218 LAYER ME3 ;
 ANTENNADIFFAREA                          0.218 LAYER ME4 ;
 ANTENNAMAXAREACAR                       10.048 LAYER ME1 ;
 ANTENNAMAXAREACAR                       12.848 LAYER ME2 ;
 ANTENNAMAXAREACAR                       15.648 LAYER ME3 ;
 ANTENNAMAXAREACAR                       18.448 LAYER ME4 ;
END DI32
PIN DO32
  DIRECTION OUTPUT ;
 PORT
  LAYER ME4 ;
  RECT 302.081 0.000 302.361 0.720 ;
  LAYER ME3 ;
  RECT 302.081 0.000 302.361 0.720 ;
  LAYER ME2 ;
  RECT 302.081 0.000 302.361 0.720 ;
  LAYER ME1 ;
  RECT 302.081 0.000 302.361 0.720 ;
 END
 ANTENNAPARTIALMETALAREA                  2.030 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME3 ;
 ANTENNADIFFAREA                          1.293 LAYER ME4 ;
END DO32
PIN WEB4
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 302.561 0.000 302.841 0.720 ;
  LAYER ME3 ;
  RECT 302.561 0.000 302.841 0.720 ;
  LAYER ME2 ;
  RECT 302.561 0.000 302.841 0.720 ;
  LAYER ME1 ;
  RECT 302.561 0.000 302.841 0.720 ;
 END
 ANTENNAPARTIALMETALAREA                  0.436 LAYER ME2 ;
 ANTENNAGATEAREA                          0.288 LAYER ME2 ;
 ANTENNAGATEAREA                          0.288 LAYER ME3 ;
 ANTENNAGATEAREA                          0.288 LAYER ME4 ;
 ANTENNADIFFAREA                          0.218 LAYER ME2 ;
 ANTENNADIFFAREA                          0.218 LAYER ME3 ;
 ANTENNADIFFAREA                          0.218 LAYER ME4 ;
 ANTENNAMAXAREACAR                        4.602 LAYER ME2 ;
 ANTENNAMAXAREACAR                        5.302 LAYER ME3 ;
 ANTENNAMAXAREACAR                        6.002 LAYER ME4 ;
END WEB4
OBS
  LAYER ME3 ;
  RECT 0.000 0.000 557.611 280.651 ;
  LAYER ME2 ;
  RECT 0.000 0.000 557.611 280.651 ;
  LAYER ME1 ;
  RECT 0.000 0.000 557.611 280.651 ;
  LAYER ME4 ;
  RECT 0.000 0.000 273.598 280.651 ;
  LAYER ME4 ;
  RECT 275.252 0.000 276.372 280.651 ;
  LAYER ME4 ;
  RECT 277.967 0.000 278.687 280.651 ;
  LAYER ME4 ;
  RECT 279.417 0.000 280.137 280.651 ;
  LAYER ME4 ;
  RECT 282.197 0.000 282.797 280.651 ;
  LAYER ME4 ;
  RECT 285.411 0.000 287.097 280.651 ;
  LAYER ME4 ;
  RECT 288.487 0.000 289.607 280.651 ;
  LAYER ME4 ;
  RECT 290.882 0.000 291.602 280.651 ;
  LAYER ME4 ;
  RECT 292.597 0.000 293.317 280.651 ;
  LAYER ME4 ;
  RECT 294.517 0.000 557.611 280.651 ;
END
END SYKB110_1024X8X8CM4
END LIBRARY





