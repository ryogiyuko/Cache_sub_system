`timescale 1ns / 1ps
//======================================================
// Project: mmu_asic
// Module:  cLastFifo1_mmu
// Author:  Yang Yuyuan
// Date:    2024/11/7
// Description: 
//======================================================

module cLastFifo1_mmu (
    input  i_drive,
    input  rstn,
    output o_free,
    output o_driveNext,
    output o_fire_1
);

    wire [1:0] w_outRRelay_2, w_outARelay_2;
    wire w_driveNext;

    (* dont_touch="true" *) sender sender (
        .i_drive(i_drive),
        .o_free (o_free),
        .outR   (w_outRRelay_2[0]),
        .i_free (o_driveNext),
        .rstn   (rstn)
    );
    (* dont_touch="true" *) relay relay (
        .inR (w_outRRelay_2[0]),
        .inA (w_outARelay_2[0]),
        .outR(w_outRRelay_2[1]),
        .outA(w_outRRelay_2[1]),
        .fire(o_fire_1),
        .rstn(rstn)
    );

    (* dont_touch="true" *) delay_mmu #(1) outdelay (
        .inR (o_fire_1),
        .outR(o_driveNext),
        .rstn(rstn)
    );

endmodule

