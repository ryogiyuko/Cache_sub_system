# ________________________________________________________________________________________________
# 
# 
#             Synchronous One-Port Register File Compiler
# 
#                 UMC 0.11um LL AE Logic Process
# 
# ________________________________________________________________________________________________
# 
#               
#         Copyright (C) 2024 Faraday Technology Corporation. All Rights Reserved.       
#                
#         This source code is an unpublished work belongs to Faraday Technology Corporation       
#         It is considered a trade secret and is not to be divulged or       
#         used by parties who have not received written authorization from       
#         Faraday Technology Corporation       
#                
#         Faraday's home page can be found at: http://www.faraday-tech.com/       
#                
# ________________________________________________________________________________________________
# 
#        IP Name            :  FSR0K_B_SY                
#        IP Version         :  1.4.0                     
#        IP Release Status  :  Active                    
#        Word               :  128                       
#        Bit                :  11                        
#        Byte               :  4                         
#        Mux                :  2                         
#        Output Loading     :  0.01                      
#        Clock Input Slew   :  0.016                     
#        Data Input Slew    :  0.016                     
#        Ring Type          :  Ringless Model            
#        Ring Width         :  0                         
#        Bus Format         :  0                         
#        Memaker Path       :  /home/mem/Desktop/memlib  
#        GUI Version        :  m20230904                 
#        Date               :  2024/09/07 15:31:53       
# ________________________________________________________________________________________________
# 

VERSION 5.5 ;
NAMESCASESENSITIVE ON ;
MACRO SYKB110_128X11X4CM2
CLASS BLOCK ;
FOREIGN SYKB110_128X11X4CM2 0.000 0.000 ;
ORIGIN 0.000 0.000 ;
SIZE 219.675 BY 111.491 ;
SYMMETRY x y r90 ;
SITE core ;
PIN GND
  DIRECTION INOUT ;
  USE GROUND ;
 PORT
  LAYER ME4 ;
  RECT 132.510 1.781 132.850 111.491 ;
 END
 PORT
  LAYER ME4 ;
  RECT 128.506 1.781 128.846 111.491 ;
 END
 PORT
  LAYER ME4 ;
  RECT 130.508 1.781 130.848 111.491 ;
 END
 PORT
  LAYER ME4 ;
  RECT 131.319 0.000 132.039 44.094 ;
 END
 PORT
  LAYER ME4 ;
  RECT 136.514 1.781 136.854 111.491 ;
 END
 PORT
  LAYER ME4 ;
  RECT 134.512 1.781 134.852 111.491 ;
 END
 PORT
  LAYER ME4 ;
  RECT 135.323 0.000 136.043 44.094 ;
 END
 PORT
  LAYER ME4 ;
  RECT 140.518 1.781 140.858 111.491 ;
 END
 PORT
  LAYER ME4 ;
  RECT 138.516 1.781 138.856 111.491 ;
 END
 PORT
  LAYER ME4 ;
  RECT 139.327 0.000 140.047 44.094 ;
 END
 PORT
  LAYER ME4 ;
  RECT 144.522 1.781 144.862 111.491 ;
 END
 PORT
  LAYER ME4 ;
  RECT 142.520 1.781 142.860 111.491 ;
 END
 PORT
  LAYER ME4 ;
  RECT 143.331 0.000 144.051 44.094 ;
 END
 PORT
  LAYER ME4 ;
  RECT 148.526 1.781 148.866 111.491 ;
 END
 PORT
  LAYER ME4 ;
  RECT 146.524 1.781 146.864 111.491 ;
 END
 PORT
  LAYER ME4 ;
  RECT 147.335 0.000 148.055 44.094 ;
 END
 PORT
  LAYER ME4 ;
  RECT 152.530 1.781 152.870 111.491 ;
 END
 PORT
  LAYER ME4 ;
  RECT 150.528 1.781 150.868 111.491 ;
 END
 PORT
  LAYER ME4 ;
  RECT 151.339 0.000 152.059 44.094 ;
 END
 PORT
  LAYER ME4 ;
  RECT 156.534 1.781 156.874 111.491 ;
 END
 PORT
  LAYER ME4 ;
  RECT 154.532 1.781 154.872 111.491 ;
 END
 PORT
  LAYER ME4 ;
  RECT 155.343 0.000 156.063 44.094 ;
 END
 PORT
  LAYER ME4 ;
  RECT 160.538 1.781 160.878 111.491 ;
 END
 PORT
  LAYER ME4 ;
  RECT 158.536 1.781 158.876 111.491 ;
 END
 PORT
  LAYER ME4 ;
  RECT 159.347 0.000 160.067 44.094 ;
 END
 PORT
  LAYER ME4 ;
  RECT 164.542 1.781 164.882 111.491 ;
 END
 PORT
  LAYER ME4 ;
  RECT 162.540 1.781 162.880 111.491 ;
 END
 PORT
  LAYER ME4 ;
  RECT 163.351 0.000 164.071 44.094 ;
 END
 PORT
  LAYER ME4 ;
  RECT 168.546 1.781 168.886 111.491 ;
 END
 PORT
  LAYER ME4 ;
  RECT 166.544 1.781 166.884 111.491 ;
 END
 PORT
  LAYER ME4 ;
  RECT 167.355 0.000 168.075 44.094 ;
 END
 PORT
  LAYER ME4 ;
  RECT 172.550 1.781 172.890 111.491 ;
 END
 PORT
  LAYER ME4 ;
  RECT 170.548 1.781 170.888 111.491 ;
 END
 PORT
  LAYER ME4 ;
  RECT 171.359 0.000 172.079 44.094 ;
 END
 PORT
  LAYER ME4 ;
  RECT 176.554 1.781 176.894 111.491 ;
 END
 PORT
  LAYER ME4 ;
  RECT 174.552 1.781 174.892 111.491 ;
 END
 PORT
  LAYER ME4 ;
  RECT 175.363 0.000 176.083 44.094 ;
 END
 PORT
  LAYER ME4 ;
  RECT 180.558 1.781 180.898 111.491 ;
 END
 PORT
  LAYER ME4 ;
  RECT 178.556 1.781 178.896 111.491 ;
 END
 PORT
  LAYER ME4 ;
  RECT 179.367 0.000 180.087 44.094 ;
 END
 PORT
  LAYER ME4 ;
  RECT 184.562 1.781 184.902 111.491 ;
 END
 PORT
  LAYER ME4 ;
  RECT 182.560 1.781 182.900 111.491 ;
 END
 PORT
  LAYER ME4 ;
  RECT 183.371 0.000 184.091 44.094 ;
 END
 PORT
  LAYER ME4 ;
  RECT 188.566 1.781 188.906 111.491 ;
 END
 PORT
  LAYER ME4 ;
  RECT 186.564 1.781 186.904 111.491 ;
 END
 PORT
  LAYER ME4 ;
  RECT 187.375 0.000 188.095 44.094 ;
 END
 PORT
  LAYER ME4 ;
  RECT 192.570 1.781 192.910 111.491 ;
 END
 PORT
  LAYER ME4 ;
  RECT 190.568 1.781 190.908 111.491 ;
 END
 PORT
  LAYER ME4 ;
  RECT 191.379 0.000 192.099 44.094 ;
 END
 PORT
  LAYER ME4 ;
  RECT 196.574 1.781 196.914 111.491 ;
 END
 PORT
  LAYER ME4 ;
  RECT 194.572 1.781 194.912 111.491 ;
 END
 PORT
  LAYER ME4 ;
  RECT 195.383 0.000 196.103 44.094 ;
 END
 PORT
  LAYER ME4 ;
  RECT 200.578 1.781 200.918 111.491 ;
 END
 PORT
  LAYER ME4 ;
  RECT 198.576 1.781 198.916 111.491 ;
 END
 PORT
  LAYER ME4 ;
  RECT 199.387 0.000 200.107 44.094 ;
 END
 PORT
  LAYER ME4 ;
  RECT 204.582 1.781 204.922 111.491 ;
 END
 PORT
  LAYER ME4 ;
  RECT 202.580 1.781 202.920 111.491 ;
 END
 PORT
  LAYER ME4 ;
  RECT 203.391 0.000 204.111 44.094 ;
 END
 PORT
  LAYER ME4 ;
  RECT 208.586 1.781 208.926 111.491 ;
 END
 PORT
  LAYER ME4 ;
  RECT 206.584 1.781 206.924 111.491 ;
 END
 PORT
  LAYER ME4 ;
  RECT 207.395 0.000 208.115 44.094 ;
 END
 PORT
  LAYER ME4 ;
  RECT 212.590 1.781 212.930 111.491 ;
 END
 PORT
  LAYER ME4 ;
  RECT 210.588 1.781 210.928 111.491 ;
 END
 PORT
  LAYER ME4 ;
  RECT 211.399 0.000 212.119 44.094 ;
 END
 PORT
  LAYER ME4 ;
  RECT 216.594 1.781 216.934 111.491 ;
 END
 PORT
  LAYER ME4 ;
  RECT 214.592 1.781 214.932 111.491 ;
 END
 PORT
  LAYER ME4 ;
  RECT 215.403 0.000 216.123 44.094 ;
 END
 PORT
  LAYER ME4 ;
  RECT 217.595 0.000 217.935 111.491 ;
 END
 PORT
  LAYER ME4 ;
  RECT 109.649 0.000 110.369 111.491 ;
 END
 PORT
  LAYER ME4 ;
  RECT 115.643 0.000 116.363 111.491 ;
 END
 PORT
  LAYER ME4 ;
  RECT 121.114 0.000 121.834 111.491 ;
 END
 PORT
  LAYER ME4 ;
  RECT 122.829 0.000 123.549 111.491 ;
 END
 PORT
  LAYER ME4 ;
  RECT 125.825 0.000 126.425 111.491 ;
 END
 PORT
  LAYER ME4 ;
  RECT 127.505 1.781 127.845 111.491 ;
 END
 PORT
  LAYER ME4 ;
  RECT 102.090 0.000 102.810 111.491 ;
 END
 PORT
  LAYER ME4 ;
  RECT 100.050 1.781 100.770 110.732 ;
 END
 PORT
  LAYER ME4 ;
  RECT 97.930 0.000 98.650 111.491 ;
 END
 PORT
  LAYER ME4 ;
  RECT 95.890 1.781 96.610 111.491 ;
 END
 PORT
  LAYER ME4 ;
  RECT 1.740 0.000 2.080 111.491 ;
 END
 PORT
  LAYER ME4 ;
  RECT 6.745 1.781 7.085 111.491 ;
 END
 PORT
  LAYER ME4 ;
  RECT 2.741 1.781 3.081 111.491 ;
 END
 PORT
  LAYER ME4 ;
  RECT 4.743 1.781 5.083 111.491 ;
 END
 PORT
  LAYER ME4 ;
  RECT 5.554 0.000 6.274 44.094 ;
 END
 PORT
  LAYER ME4 ;
  RECT 10.749 1.781 11.089 111.491 ;
 END
 PORT
  LAYER ME4 ;
  RECT 8.747 1.781 9.087 111.491 ;
 END
 PORT
  LAYER ME4 ;
  RECT 9.558 0.000 10.278 44.094 ;
 END
 PORT
  LAYER ME4 ;
  RECT 14.753 1.781 15.093 111.491 ;
 END
 PORT
  LAYER ME4 ;
  RECT 12.751 1.781 13.091 111.491 ;
 END
 PORT
  LAYER ME4 ;
  RECT 13.562 0.000 14.282 44.094 ;
 END
 PORT
  LAYER ME4 ;
  RECT 18.757 1.781 19.097 111.491 ;
 END
 PORT
  LAYER ME4 ;
  RECT 16.755 1.781 17.095 111.491 ;
 END
 PORT
  LAYER ME4 ;
  RECT 17.566 0.000 18.286 44.094 ;
 END
 PORT
  LAYER ME4 ;
  RECT 22.761 1.781 23.101 111.491 ;
 END
 PORT
  LAYER ME4 ;
  RECT 20.759 1.781 21.099 111.491 ;
 END
 PORT
  LAYER ME4 ;
  RECT 21.570 0.000 22.290 44.094 ;
 END
 PORT
  LAYER ME4 ;
  RECT 26.765 1.781 27.105 111.491 ;
 END
 PORT
  LAYER ME4 ;
  RECT 24.763 1.781 25.103 111.491 ;
 END
 PORT
  LAYER ME4 ;
  RECT 25.574 0.000 26.294 44.094 ;
 END
 PORT
  LAYER ME4 ;
  RECT 30.769 1.781 31.109 111.491 ;
 END
 PORT
  LAYER ME4 ;
  RECT 28.767 1.781 29.107 111.491 ;
 END
 PORT
  LAYER ME4 ;
  RECT 29.578 0.000 30.298 44.094 ;
 END
 PORT
  LAYER ME4 ;
  RECT 34.773 1.781 35.113 111.491 ;
 END
 PORT
  LAYER ME4 ;
  RECT 32.771 1.781 33.111 111.491 ;
 END
 PORT
  LAYER ME4 ;
  RECT 33.582 0.000 34.302 44.094 ;
 END
 PORT
  LAYER ME4 ;
  RECT 38.777 1.781 39.117 111.491 ;
 END
 PORT
  LAYER ME4 ;
  RECT 36.775 1.781 37.115 111.491 ;
 END
 PORT
  LAYER ME4 ;
  RECT 37.586 0.000 38.306 44.094 ;
 END
 PORT
  LAYER ME4 ;
  RECT 42.781 1.781 43.121 111.491 ;
 END
 PORT
  LAYER ME4 ;
  RECT 40.779 1.781 41.119 111.491 ;
 END
 PORT
  LAYER ME4 ;
  RECT 41.590 0.000 42.310 44.094 ;
 END
 PORT
  LAYER ME4 ;
  RECT 46.785 1.781 47.125 111.491 ;
 END
 PORT
  LAYER ME4 ;
  RECT 44.783 1.781 45.123 111.491 ;
 END
 PORT
  LAYER ME4 ;
  RECT 45.594 0.000 46.314 44.094 ;
 END
 PORT
  LAYER ME4 ;
  RECT 50.789 1.781 51.129 111.491 ;
 END
 PORT
  LAYER ME4 ;
  RECT 48.787 1.781 49.127 111.491 ;
 END
 PORT
  LAYER ME4 ;
  RECT 49.598 0.000 50.318 44.094 ;
 END
 PORT
  LAYER ME4 ;
  RECT 54.793 1.781 55.133 111.491 ;
 END
 PORT
  LAYER ME4 ;
  RECT 52.791 1.781 53.131 111.491 ;
 END
 PORT
  LAYER ME4 ;
  RECT 53.602 0.000 54.322 44.094 ;
 END
 PORT
  LAYER ME4 ;
  RECT 58.797 1.781 59.137 111.491 ;
 END
 PORT
  LAYER ME4 ;
  RECT 56.795 1.781 57.135 111.491 ;
 END
 PORT
  LAYER ME4 ;
  RECT 57.606 0.000 58.326 44.094 ;
 END
 PORT
  LAYER ME4 ;
  RECT 62.801 1.781 63.141 111.491 ;
 END
 PORT
  LAYER ME4 ;
  RECT 60.799 1.781 61.139 111.491 ;
 END
 PORT
  LAYER ME4 ;
  RECT 61.610 0.000 62.330 44.094 ;
 END
 PORT
  LAYER ME4 ;
  RECT 66.805 1.781 67.145 111.491 ;
 END
 PORT
  LAYER ME4 ;
  RECT 64.803 1.781 65.143 111.491 ;
 END
 PORT
  LAYER ME4 ;
  RECT 65.614 0.000 66.334 44.094 ;
 END
 PORT
  LAYER ME4 ;
  RECT 70.809 1.781 71.149 111.491 ;
 END
 PORT
  LAYER ME4 ;
  RECT 68.807 1.781 69.147 111.491 ;
 END
 PORT
  LAYER ME4 ;
  RECT 69.618 0.000 70.338 44.094 ;
 END
 PORT
  LAYER ME4 ;
  RECT 74.813 1.781 75.153 111.491 ;
 END
 PORT
  LAYER ME4 ;
  RECT 72.811 1.781 73.151 111.491 ;
 END
 PORT
  LAYER ME4 ;
  RECT 73.622 0.000 74.342 44.094 ;
 END
 PORT
  LAYER ME4 ;
  RECT 78.817 1.781 79.157 111.491 ;
 END
 PORT
  LAYER ME4 ;
  RECT 76.815 1.781 77.155 111.491 ;
 END
 PORT
  LAYER ME4 ;
  RECT 77.626 0.000 78.346 44.094 ;
 END
 PORT
  LAYER ME4 ;
  RECT 82.821 1.781 83.161 111.491 ;
 END
 PORT
  LAYER ME4 ;
  RECT 80.819 1.781 81.159 111.491 ;
 END
 PORT
  LAYER ME4 ;
  RECT 81.630 0.000 82.350 44.094 ;
 END
 PORT
  LAYER ME4 ;
  RECT 86.825 1.781 87.165 111.491 ;
 END
 PORT
  LAYER ME4 ;
  RECT 84.823 1.781 85.163 111.491 ;
 END
 PORT
  LAYER ME4 ;
  RECT 85.634 0.000 86.354 44.094 ;
 END
 PORT
  LAYER ME4 ;
  RECT 90.829 1.781 91.169 111.491 ;
 END
 PORT
  LAYER ME4 ;
  RECT 88.827 1.781 89.167 111.491 ;
 END
 PORT
  LAYER ME4 ;
  RECT 89.638 0.000 90.358 44.094 ;
 END
 PORT
  LAYER ME4 ;
  RECT 93.770 0.000 94.490 111.491 ;
 END
 PORT
  LAYER ME4 ;
  RECT 91.830 0.000 92.170 111.491 ;
 END
END GND
PIN VCC
  DIRECTION INOUT ;
  USE POWER ;
 PORT
  LAYER ME4 ;
  RECT 131.509 45.394 131.849 111.491 ;
 END
 PORT
  LAYER ME4 ;
  RECT 129.317 0.000 130.037 46.394 ;
 END
 PORT
  LAYER ME4 ;
  RECT 135.513 45.394 135.853 111.491 ;
 END
 PORT
  LAYER ME4 ;
  RECT 133.321 0.000 134.041 46.394 ;
 END
 PORT
  LAYER ME4 ;
  RECT 139.517 45.394 139.857 111.491 ;
 END
 PORT
  LAYER ME4 ;
  RECT 137.325 0.000 138.045 46.394 ;
 END
 PORT
  LAYER ME4 ;
  RECT 143.521 45.394 143.861 111.491 ;
 END
 PORT
  LAYER ME4 ;
  RECT 141.329 0.000 142.049 46.394 ;
 END
 PORT
  LAYER ME4 ;
  RECT 147.525 45.394 147.865 111.491 ;
 END
 PORT
  LAYER ME4 ;
  RECT 145.333 0.000 146.053 46.394 ;
 END
 PORT
  LAYER ME4 ;
  RECT 151.529 45.394 151.869 111.491 ;
 END
 PORT
  LAYER ME4 ;
  RECT 149.337 0.000 150.057 46.394 ;
 END
 PORT
  LAYER ME4 ;
  RECT 155.533 45.394 155.873 111.491 ;
 END
 PORT
  LAYER ME4 ;
  RECT 153.341 0.000 154.061 46.394 ;
 END
 PORT
  LAYER ME4 ;
  RECT 159.537 45.394 159.877 111.491 ;
 END
 PORT
  LAYER ME4 ;
  RECT 157.345 0.000 158.065 46.394 ;
 END
 PORT
  LAYER ME4 ;
  RECT 163.541 45.394 163.881 111.491 ;
 END
 PORT
  LAYER ME4 ;
  RECT 161.349 0.000 162.069 46.394 ;
 END
 PORT
  LAYER ME4 ;
  RECT 167.545 45.394 167.885 111.491 ;
 END
 PORT
  LAYER ME4 ;
  RECT 165.353 0.000 166.073 46.394 ;
 END
 PORT
  LAYER ME4 ;
  RECT 171.549 45.394 171.889 111.491 ;
 END
 PORT
  LAYER ME4 ;
  RECT 169.357 0.000 170.077 46.394 ;
 END
 PORT
  LAYER ME4 ;
  RECT 175.553 45.394 175.893 111.491 ;
 END
 PORT
  LAYER ME4 ;
  RECT 173.361 0.000 174.081 46.394 ;
 END
 PORT
  LAYER ME4 ;
  RECT 179.557 45.394 179.897 111.491 ;
 END
 PORT
  LAYER ME4 ;
  RECT 177.365 0.000 178.085 46.394 ;
 END
 PORT
  LAYER ME4 ;
  RECT 183.561 45.394 183.901 111.491 ;
 END
 PORT
  LAYER ME4 ;
  RECT 181.369 0.000 182.089 46.394 ;
 END
 PORT
  LAYER ME4 ;
  RECT 187.565 45.394 187.905 111.491 ;
 END
 PORT
  LAYER ME4 ;
  RECT 185.373 0.000 186.093 46.394 ;
 END
 PORT
  LAYER ME4 ;
  RECT 191.569 45.394 191.909 111.491 ;
 END
 PORT
  LAYER ME4 ;
  RECT 189.377 0.000 190.097 46.394 ;
 END
 PORT
  LAYER ME4 ;
  RECT 195.573 45.394 195.913 111.491 ;
 END
 PORT
  LAYER ME4 ;
  RECT 193.381 0.000 194.101 46.394 ;
 END
 PORT
  LAYER ME4 ;
  RECT 199.577 45.394 199.917 111.491 ;
 END
 PORT
  LAYER ME4 ;
  RECT 197.385 0.000 198.105 46.394 ;
 END
 PORT
  LAYER ME4 ;
  RECT 203.581 45.394 203.921 111.491 ;
 END
 PORT
  LAYER ME4 ;
  RECT 201.389 0.000 202.109 46.394 ;
 END
 PORT
  LAYER ME4 ;
  RECT 207.585 45.394 207.925 111.491 ;
 END
 PORT
  LAYER ME4 ;
  RECT 205.393 0.000 206.113 46.394 ;
 END
 PORT
  LAYER ME4 ;
  RECT 211.589 45.394 211.929 111.491 ;
 END
 PORT
  LAYER ME4 ;
  RECT 209.397 0.000 210.117 46.394 ;
 END
 PORT
  LAYER ME4 ;
  RECT 215.593 45.394 215.933 111.491 ;
 END
 PORT
  LAYER ME4 ;
  RECT 213.401 0.000 214.121 46.394 ;
 END
 PORT
  LAYER ME4 ;
  RECT 218.375 0.000 218.755 111.491 ;
 END
 PORT
  LAYER ME4 ;
  RECT 112.429 0.000 113.029 111.491 ;
 END
 PORT
  LAYER ME4 ;
  RECT 116.609 0.000 117.329 111.491 ;
 END
 PORT
  LAYER ME4 ;
  RECT 118.719 0.000 119.839 111.491 ;
 END
 PORT
  LAYER ME4 ;
  RECT 124.749 0.000 125.469 111.491 ;
 END
 PORT
  LAYER ME4 ;
  RECT 126.685 1.781 127.065 111.491 ;
 END
 PORT
  LAYER ME4 ;
  RECT 108.199 0.000 108.919 111.491 ;
 END
 PORT
  LAYER ME4 ;
  RECT 105.484 0.000 106.604 111.491 ;
 END
 PORT
  LAYER ME4 ;
  RECT 103.110 0.000 103.830 110.732 ;
 END
 PORT
  LAYER ME4 ;
  RECT 101.070 1.781 101.790 111.491 ;
 END
 PORT
  LAYER ME4 ;
  RECT 98.950 0.000 99.670 111.491 ;
 END
 PORT
  LAYER ME4 ;
  RECT 96.910 1.781 97.630 111.491 ;
 END
 PORT
  LAYER ME4 ;
  RECT 0.920 0.000 1.300 111.491 ;
 END
 PORT
  LAYER ME4 ;
  RECT 5.744 45.394 6.084 111.491 ;
 END
 PORT
  LAYER ME4 ;
  RECT 3.552 0.000 4.272 46.394 ;
 END
 PORT
  LAYER ME4 ;
  RECT 9.748 45.394 10.088 111.491 ;
 END
 PORT
  LAYER ME4 ;
  RECT 7.556 0.000 8.276 46.394 ;
 END
 PORT
  LAYER ME4 ;
  RECT 13.752 45.394 14.092 111.491 ;
 END
 PORT
  LAYER ME4 ;
  RECT 11.560 0.000 12.280 46.394 ;
 END
 PORT
  LAYER ME4 ;
  RECT 17.756 45.394 18.096 111.491 ;
 END
 PORT
  LAYER ME4 ;
  RECT 15.564 0.000 16.284 46.394 ;
 END
 PORT
  LAYER ME4 ;
  RECT 21.760 45.394 22.100 111.491 ;
 END
 PORT
  LAYER ME4 ;
  RECT 19.568 0.000 20.288 46.394 ;
 END
 PORT
  LAYER ME4 ;
  RECT 25.764 45.394 26.104 111.491 ;
 END
 PORT
  LAYER ME4 ;
  RECT 23.572 0.000 24.292 46.394 ;
 END
 PORT
  LAYER ME4 ;
  RECT 29.768 45.394 30.108 111.491 ;
 END
 PORT
  LAYER ME4 ;
  RECT 27.576 0.000 28.296 46.394 ;
 END
 PORT
  LAYER ME4 ;
  RECT 33.772 45.394 34.112 111.491 ;
 END
 PORT
  LAYER ME4 ;
  RECT 31.580 0.000 32.300 46.394 ;
 END
 PORT
  LAYER ME4 ;
  RECT 37.776 45.394 38.116 111.491 ;
 END
 PORT
  LAYER ME4 ;
  RECT 35.584 0.000 36.304 46.394 ;
 END
 PORT
  LAYER ME4 ;
  RECT 41.780 45.394 42.120 111.491 ;
 END
 PORT
  LAYER ME4 ;
  RECT 39.588 0.000 40.308 46.394 ;
 END
 PORT
  LAYER ME4 ;
  RECT 45.784 45.394 46.124 111.491 ;
 END
 PORT
  LAYER ME4 ;
  RECT 43.592 0.000 44.312 46.394 ;
 END
 PORT
  LAYER ME4 ;
  RECT 49.788 45.394 50.128 111.491 ;
 END
 PORT
  LAYER ME4 ;
  RECT 47.596 0.000 48.316 46.394 ;
 END
 PORT
  LAYER ME4 ;
  RECT 53.792 45.394 54.132 111.491 ;
 END
 PORT
  LAYER ME4 ;
  RECT 51.600 0.000 52.320 46.394 ;
 END
 PORT
  LAYER ME4 ;
  RECT 57.796 45.394 58.136 111.491 ;
 END
 PORT
  LAYER ME4 ;
  RECT 55.604 0.000 56.324 46.394 ;
 END
 PORT
  LAYER ME4 ;
  RECT 61.800 45.394 62.140 111.491 ;
 END
 PORT
  LAYER ME4 ;
  RECT 59.608 0.000 60.328 46.394 ;
 END
 PORT
  LAYER ME4 ;
  RECT 65.804 45.394 66.144 111.491 ;
 END
 PORT
  LAYER ME4 ;
  RECT 63.612 0.000 64.332 46.394 ;
 END
 PORT
  LAYER ME4 ;
  RECT 69.808 45.394 70.148 111.491 ;
 END
 PORT
  LAYER ME4 ;
  RECT 67.616 0.000 68.336 46.394 ;
 END
 PORT
  LAYER ME4 ;
  RECT 73.812 45.394 74.152 111.491 ;
 END
 PORT
  LAYER ME4 ;
  RECT 71.620 0.000 72.340 46.394 ;
 END
 PORT
  LAYER ME4 ;
  RECT 77.816 45.394 78.156 111.491 ;
 END
 PORT
  LAYER ME4 ;
  RECT 75.624 0.000 76.344 46.394 ;
 END
 PORT
  LAYER ME4 ;
  RECT 81.820 45.394 82.160 111.491 ;
 END
 PORT
  LAYER ME4 ;
  RECT 79.628 0.000 80.348 46.394 ;
 END
 PORT
  LAYER ME4 ;
  RECT 85.824 45.394 86.164 111.491 ;
 END
 PORT
  LAYER ME4 ;
  RECT 83.632 0.000 84.352 46.394 ;
 END
 PORT
  LAYER ME4 ;
  RECT 89.828 45.394 90.168 111.491 ;
 END
 PORT
  LAYER ME4 ;
  RECT 87.636 0.000 88.356 46.394 ;
 END
 PORT
  LAYER ME4 ;
  RECT 94.790 0.000 95.510 111.491 ;
 END
 PORT
  LAYER ME4 ;
  RECT 92.610 0.000 92.990 111.491 ;
 END
 PORT
  LAYER ME4 ;
  RECT 129.507 47.744 129.847 111.491 ;
 END
 PORT
  LAYER ME4 ;
  RECT 133.511 47.744 133.851 111.491 ;
 END
 PORT
  LAYER ME4 ;
  RECT 137.515 47.744 137.855 111.491 ;
 END
 PORT
  LAYER ME4 ;
  RECT 141.519 47.744 141.859 111.491 ;
 END
 PORT
  LAYER ME4 ;
  RECT 145.523 47.744 145.863 111.491 ;
 END
 PORT
  LAYER ME4 ;
  RECT 149.527 47.744 149.867 111.491 ;
 END
 PORT
  LAYER ME4 ;
  RECT 153.531 47.744 153.871 111.491 ;
 END
 PORT
  LAYER ME4 ;
  RECT 157.535 47.744 157.875 111.491 ;
 END
 PORT
  LAYER ME4 ;
  RECT 161.539 47.744 161.879 111.491 ;
 END
 PORT
  LAYER ME4 ;
  RECT 165.543 47.744 165.883 111.491 ;
 END
 PORT
  LAYER ME4 ;
  RECT 169.547 47.744 169.887 111.491 ;
 END
 PORT
  LAYER ME4 ;
  RECT 173.551 47.744 173.891 111.491 ;
 END
 PORT
  LAYER ME4 ;
  RECT 177.555 47.744 177.895 111.491 ;
 END
 PORT
  LAYER ME4 ;
  RECT 181.559 47.744 181.899 111.491 ;
 END
 PORT
  LAYER ME4 ;
  RECT 185.563 47.744 185.903 111.491 ;
 END
 PORT
  LAYER ME4 ;
  RECT 189.567 47.744 189.907 111.491 ;
 END
 PORT
  LAYER ME4 ;
  RECT 193.571 47.744 193.911 111.491 ;
 END
 PORT
  LAYER ME4 ;
  RECT 197.575 47.744 197.915 111.491 ;
 END
 PORT
  LAYER ME4 ;
  RECT 201.579 47.744 201.919 111.491 ;
 END
 PORT
  LAYER ME4 ;
  RECT 205.583 47.744 205.923 111.491 ;
 END
 PORT
  LAYER ME4 ;
  RECT 209.587 47.744 209.927 111.491 ;
 END
 PORT
  LAYER ME4 ;
  RECT 213.591 47.744 213.931 111.491 ;
 END
 PORT
  LAYER ME4 ;
  RECT 3.742 47.744 4.082 111.491 ;
 END
 PORT
  LAYER ME4 ;
  RECT 7.746 47.744 8.086 111.491 ;
 END
 PORT
  LAYER ME4 ;
  RECT 11.750 47.744 12.090 111.491 ;
 END
 PORT
  LAYER ME4 ;
  RECT 15.754 47.744 16.094 111.491 ;
 END
 PORT
  LAYER ME4 ;
  RECT 19.758 47.744 20.098 111.491 ;
 END
 PORT
  LAYER ME4 ;
  RECT 23.762 47.744 24.102 111.491 ;
 END
 PORT
  LAYER ME4 ;
  RECT 27.766 47.744 28.106 111.491 ;
 END
 PORT
  LAYER ME4 ;
  RECT 31.770 47.744 32.110 111.491 ;
 END
 PORT
  LAYER ME4 ;
  RECT 35.774 47.744 36.114 111.491 ;
 END
 PORT
  LAYER ME4 ;
  RECT 39.778 47.744 40.118 111.491 ;
 END
 PORT
  LAYER ME4 ;
  RECT 43.782 47.744 44.122 111.491 ;
 END
 PORT
  LAYER ME4 ;
  RECT 47.786 47.744 48.126 111.491 ;
 END
 PORT
  LAYER ME4 ;
  RECT 51.790 47.744 52.130 111.491 ;
 END
 PORT
  LAYER ME4 ;
  RECT 55.794 47.744 56.134 111.491 ;
 END
 PORT
  LAYER ME4 ;
  RECT 59.798 47.744 60.138 111.491 ;
 END
 PORT
  LAYER ME4 ;
  RECT 63.802 47.744 64.142 111.491 ;
 END
 PORT
  LAYER ME4 ;
  RECT 67.806 47.744 68.146 111.491 ;
 END
 PORT
  LAYER ME4 ;
  RECT 71.810 47.744 72.150 111.491 ;
 END
 PORT
  LAYER ME4 ;
  RECT 75.814 47.744 76.154 111.491 ;
 END
 PORT
  LAYER ME4 ;
  RECT 79.818 47.744 80.158 111.491 ;
 END
 PORT
  LAYER ME4 ;
  RECT 83.822 47.744 84.162 111.491 ;
 END
 PORT
  LAYER ME4 ;
  RECT 87.826 47.744 88.166 111.491 ;
 END
END VCC
PIN DI21
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 89.118 0.000 89.438 0.600 ;
  LAYER ME3 ;
  RECT 89.118 0.000 89.438 0.600 ;
  LAYER ME2 ;
  RECT 89.118 0.000 89.438 0.600 ;
  LAYER ME1 ;
  RECT 89.118 0.000 89.438 0.600 ;
 END
 ANTENNAPARTIALMETALAREA                  1.058 LAYER ME2 ;
 ANTENNAGATEAREA                          0.072 LAYER ME2 ;
 ANTENNAGATEAREA                          0.072 LAYER ME3 ;
 ANTENNAGATEAREA                          0.072 LAYER ME4 ;
 ANTENNADIFFAREA                          0.160 LAYER ME2 ;
 ANTENNADIFFAREA                          0.160 LAYER ME3 ;
 ANTENNADIFFAREA                          0.160 LAYER ME4 ;
 ANTENNAMAXAREACAR                       21.782 LAYER ME2 ;
 ANTENNAMAXAREACAR                       24.449 LAYER ME3 ;
 ANTENNAMAXAREACAR                       27.116 LAYER ME4 ;
END DI21
PIN DO21
  DIRECTION OUTPUT ;
 PORT
  LAYER ME4 ;
  RECT 88.556 0.000 88.876 0.600 ;
  LAYER ME3 ;
  RECT 88.556 0.000 88.876 0.600 ;
  LAYER ME2 ;
  RECT 88.556 0.000 88.876 0.600 ;
  LAYER ME1 ;
  RECT 88.556 0.000 88.876 0.600 ;
 END
 ANTENNAPARTIALMETALAREA                  5.273 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME3 ;
 ANTENNADIFFAREA                          1.293 LAYER ME4 ;
END DO21
PIN DI20
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 85.114 0.000 85.434 0.600 ;
  LAYER ME3 ;
  RECT 85.114 0.000 85.434 0.600 ;
  LAYER ME2 ;
  RECT 85.114 0.000 85.434 0.600 ;
  LAYER ME1 ;
  RECT 85.114 0.000 85.434 0.600 ;
 END
 ANTENNAPARTIALMETALAREA                  1.058 LAYER ME2 ;
 ANTENNAGATEAREA                          0.072 LAYER ME2 ;
 ANTENNAGATEAREA                          0.072 LAYER ME3 ;
 ANTENNAGATEAREA                          0.072 LAYER ME4 ;
 ANTENNADIFFAREA                          0.160 LAYER ME2 ;
 ANTENNADIFFAREA                          0.160 LAYER ME3 ;
 ANTENNADIFFAREA                          0.160 LAYER ME4 ;
 ANTENNAMAXAREACAR                       21.782 LAYER ME2 ;
 ANTENNAMAXAREACAR                       24.449 LAYER ME3 ;
 ANTENNAMAXAREACAR                       27.116 LAYER ME4 ;
END DI20
PIN DO20
  DIRECTION OUTPUT ;
 PORT
  LAYER ME4 ;
  RECT 84.552 0.000 84.872 0.600 ;
  LAYER ME3 ;
  RECT 84.552 0.000 84.872 0.600 ;
  LAYER ME2 ;
  RECT 84.552 0.000 84.872 0.600 ;
  LAYER ME1 ;
  RECT 84.552 0.000 84.872 0.600 ;
 END
 ANTENNAPARTIALMETALAREA                  5.273 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME3 ;
 ANTENNADIFFAREA                          1.293 LAYER ME4 ;
END DO20
PIN DI19
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 81.110 0.000 81.430 0.600 ;
  LAYER ME3 ;
  RECT 81.110 0.000 81.430 0.600 ;
  LAYER ME2 ;
  RECT 81.110 0.000 81.430 0.600 ;
  LAYER ME1 ;
  RECT 81.110 0.000 81.430 0.600 ;
 END
 ANTENNAPARTIALMETALAREA                  1.058 LAYER ME2 ;
 ANTENNAGATEAREA                          0.072 LAYER ME2 ;
 ANTENNAGATEAREA                          0.072 LAYER ME3 ;
 ANTENNAGATEAREA                          0.072 LAYER ME4 ;
 ANTENNADIFFAREA                          0.160 LAYER ME2 ;
 ANTENNADIFFAREA                          0.160 LAYER ME3 ;
 ANTENNADIFFAREA                          0.160 LAYER ME4 ;
 ANTENNAMAXAREACAR                       21.782 LAYER ME2 ;
 ANTENNAMAXAREACAR                       24.449 LAYER ME3 ;
 ANTENNAMAXAREACAR                       27.116 LAYER ME4 ;
END DI19
PIN DO19
  DIRECTION OUTPUT ;
 PORT
  LAYER ME4 ;
  RECT 80.548 0.000 80.868 0.600 ;
  LAYER ME3 ;
  RECT 80.548 0.000 80.868 0.600 ;
  LAYER ME2 ;
  RECT 80.548 0.000 80.868 0.600 ;
  LAYER ME1 ;
  RECT 80.548 0.000 80.868 0.600 ;
 END
 ANTENNAPARTIALMETALAREA                  5.273 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME3 ;
 ANTENNADIFFAREA                          1.293 LAYER ME4 ;
END DO19
PIN DI18
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 77.106 0.000 77.426 0.600 ;
  LAYER ME3 ;
  RECT 77.106 0.000 77.426 0.600 ;
  LAYER ME2 ;
  RECT 77.106 0.000 77.426 0.600 ;
  LAYER ME1 ;
  RECT 77.106 0.000 77.426 0.600 ;
 END
 ANTENNAPARTIALMETALAREA                  1.058 LAYER ME2 ;
 ANTENNAGATEAREA                          0.072 LAYER ME2 ;
 ANTENNAGATEAREA                          0.072 LAYER ME3 ;
 ANTENNAGATEAREA                          0.072 LAYER ME4 ;
 ANTENNADIFFAREA                          0.160 LAYER ME2 ;
 ANTENNADIFFAREA                          0.160 LAYER ME3 ;
 ANTENNADIFFAREA                          0.160 LAYER ME4 ;
 ANTENNAMAXAREACAR                       21.782 LAYER ME2 ;
 ANTENNAMAXAREACAR                       24.449 LAYER ME3 ;
 ANTENNAMAXAREACAR                       27.116 LAYER ME4 ;
END DI18
PIN DO18
  DIRECTION OUTPUT ;
 PORT
  LAYER ME4 ;
  RECT 76.544 0.000 76.864 0.600 ;
  LAYER ME3 ;
  RECT 76.544 0.000 76.864 0.600 ;
  LAYER ME2 ;
  RECT 76.544 0.000 76.864 0.600 ;
  LAYER ME1 ;
  RECT 76.544 0.000 76.864 0.600 ;
 END
 ANTENNAPARTIALMETALAREA                  5.273 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME3 ;
 ANTENNADIFFAREA                          1.293 LAYER ME4 ;
END DO18
PIN DI17
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 73.102 0.000 73.422 0.600 ;
  LAYER ME3 ;
  RECT 73.102 0.000 73.422 0.600 ;
  LAYER ME2 ;
  RECT 73.102 0.000 73.422 0.600 ;
  LAYER ME1 ;
  RECT 73.102 0.000 73.422 0.600 ;
 END
 ANTENNAPARTIALMETALAREA                  1.058 LAYER ME2 ;
 ANTENNAGATEAREA                          0.072 LAYER ME2 ;
 ANTENNAGATEAREA                          0.072 LAYER ME3 ;
 ANTENNAGATEAREA                          0.072 LAYER ME4 ;
 ANTENNADIFFAREA                          0.160 LAYER ME2 ;
 ANTENNADIFFAREA                          0.160 LAYER ME3 ;
 ANTENNADIFFAREA                          0.160 LAYER ME4 ;
 ANTENNAMAXAREACAR                       21.782 LAYER ME2 ;
 ANTENNAMAXAREACAR                       24.449 LAYER ME3 ;
 ANTENNAMAXAREACAR                       27.116 LAYER ME4 ;
END DI17
PIN DO17
  DIRECTION OUTPUT ;
 PORT
  LAYER ME4 ;
  RECT 72.540 0.000 72.860 0.600 ;
  LAYER ME3 ;
  RECT 72.540 0.000 72.860 0.600 ;
  LAYER ME2 ;
  RECT 72.540 0.000 72.860 0.600 ;
  LAYER ME1 ;
  RECT 72.540 0.000 72.860 0.600 ;
 END
 ANTENNAPARTIALMETALAREA                  5.273 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME3 ;
 ANTENNADIFFAREA                          1.293 LAYER ME4 ;
END DO17
PIN DI16
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 69.098 0.000 69.418 0.600 ;
  LAYER ME3 ;
  RECT 69.098 0.000 69.418 0.600 ;
  LAYER ME2 ;
  RECT 69.098 0.000 69.418 0.600 ;
  LAYER ME1 ;
  RECT 69.098 0.000 69.418 0.600 ;
 END
 ANTENNAPARTIALMETALAREA                  1.058 LAYER ME2 ;
 ANTENNAGATEAREA                          0.072 LAYER ME2 ;
 ANTENNAGATEAREA                          0.072 LAYER ME3 ;
 ANTENNAGATEAREA                          0.072 LAYER ME4 ;
 ANTENNADIFFAREA                          0.160 LAYER ME2 ;
 ANTENNADIFFAREA                          0.160 LAYER ME3 ;
 ANTENNADIFFAREA                          0.160 LAYER ME4 ;
 ANTENNAMAXAREACAR                       21.782 LAYER ME2 ;
 ANTENNAMAXAREACAR                       24.449 LAYER ME3 ;
 ANTENNAMAXAREACAR                       27.116 LAYER ME4 ;
END DI16
PIN DO16
  DIRECTION OUTPUT ;
 PORT
  LAYER ME4 ;
  RECT 68.536 0.000 68.856 0.600 ;
  LAYER ME3 ;
  RECT 68.536 0.000 68.856 0.600 ;
  LAYER ME2 ;
  RECT 68.536 0.000 68.856 0.600 ;
  LAYER ME1 ;
  RECT 68.536 0.000 68.856 0.600 ;
 END
 ANTENNAPARTIALMETALAREA                  5.273 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME3 ;
 ANTENNADIFFAREA                          1.293 LAYER ME4 ;
END DO16
PIN DI15
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 65.094 0.000 65.414 0.600 ;
  LAYER ME3 ;
  RECT 65.094 0.000 65.414 0.600 ;
  LAYER ME2 ;
  RECT 65.094 0.000 65.414 0.600 ;
  LAYER ME1 ;
  RECT 65.094 0.000 65.414 0.600 ;
 END
 ANTENNAPARTIALMETALAREA                  1.058 LAYER ME2 ;
 ANTENNAGATEAREA                          0.072 LAYER ME2 ;
 ANTENNAGATEAREA                          0.072 LAYER ME3 ;
 ANTENNAGATEAREA                          0.072 LAYER ME4 ;
 ANTENNADIFFAREA                          0.160 LAYER ME2 ;
 ANTENNADIFFAREA                          0.160 LAYER ME3 ;
 ANTENNADIFFAREA                          0.160 LAYER ME4 ;
 ANTENNAMAXAREACAR                       21.782 LAYER ME2 ;
 ANTENNAMAXAREACAR                       24.449 LAYER ME3 ;
 ANTENNAMAXAREACAR                       27.116 LAYER ME4 ;
END DI15
PIN DO15
  DIRECTION OUTPUT ;
 PORT
  LAYER ME4 ;
  RECT 64.532 0.000 64.852 0.600 ;
  LAYER ME3 ;
  RECT 64.532 0.000 64.852 0.600 ;
  LAYER ME2 ;
  RECT 64.532 0.000 64.852 0.600 ;
  LAYER ME1 ;
  RECT 64.532 0.000 64.852 0.600 ;
 END
 ANTENNAPARTIALMETALAREA                  5.273 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME3 ;
 ANTENNADIFFAREA                          1.293 LAYER ME4 ;
END DO15
PIN DI14
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 61.090 0.000 61.410 0.600 ;
  LAYER ME3 ;
  RECT 61.090 0.000 61.410 0.600 ;
  LAYER ME2 ;
  RECT 61.090 0.000 61.410 0.600 ;
  LAYER ME1 ;
  RECT 61.090 0.000 61.410 0.600 ;
 END
 ANTENNAPARTIALMETALAREA                  1.058 LAYER ME2 ;
 ANTENNAGATEAREA                          0.072 LAYER ME2 ;
 ANTENNAGATEAREA                          0.072 LAYER ME3 ;
 ANTENNAGATEAREA                          0.072 LAYER ME4 ;
 ANTENNADIFFAREA                          0.160 LAYER ME2 ;
 ANTENNADIFFAREA                          0.160 LAYER ME3 ;
 ANTENNADIFFAREA                          0.160 LAYER ME4 ;
 ANTENNAMAXAREACAR                       21.782 LAYER ME2 ;
 ANTENNAMAXAREACAR                       24.449 LAYER ME3 ;
 ANTENNAMAXAREACAR                       27.116 LAYER ME4 ;
END DI14
PIN DO14
  DIRECTION OUTPUT ;
 PORT
  LAYER ME4 ;
  RECT 60.528 0.000 60.848 0.600 ;
  LAYER ME3 ;
  RECT 60.528 0.000 60.848 0.600 ;
  LAYER ME2 ;
  RECT 60.528 0.000 60.848 0.600 ;
  LAYER ME1 ;
  RECT 60.528 0.000 60.848 0.600 ;
 END
 ANTENNAPARTIALMETALAREA                  5.273 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME3 ;
 ANTENNADIFFAREA                          1.293 LAYER ME4 ;
END DO14
PIN DI13
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 57.086 0.000 57.406 0.600 ;
  LAYER ME3 ;
  RECT 57.086 0.000 57.406 0.600 ;
  LAYER ME2 ;
  RECT 57.086 0.000 57.406 0.600 ;
  LAYER ME1 ;
  RECT 57.086 0.000 57.406 0.600 ;
 END
 ANTENNAPARTIALMETALAREA                  1.058 LAYER ME2 ;
 ANTENNAGATEAREA                          0.072 LAYER ME2 ;
 ANTENNAGATEAREA                          0.072 LAYER ME3 ;
 ANTENNAGATEAREA                          0.072 LAYER ME4 ;
 ANTENNADIFFAREA                          0.160 LAYER ME2 ;
 ANTENNADIFFAREA                          0.160 LAYER ME3 ;
 ANTENNADIFFAREA                          0.160 LAYER ME4 ;
 ANTENNAMAXAREACAR                       21.782 LAYER ME2 ;
 ANTENNAMAXAREACAR                       24.449 LAYER ME3 ;
 ANTENNAMAXAREACAR                       27.116 LAYER ME4 ;
END DI13
PIN DO13
  DIRECTION OUTPUT ;
 PORT
  LAYER ME4 ;
  RECT 56.524 0.000 56.844 0.600 ;
  LAYER ME3 ;
  RECT 56.524 0.000 56.844 0.600 ;
  LAYER ME2 ;
  RECT 56.524 0.000 56.844 0.600 ;
  LAYER ME1 ;
  RECT 56.524 0.000 56.844 0.600 ;
 END
 ANTENNAPARTIALMETALAREA                  5.273 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME3 ;
 ANTENNADIFFAREA                          1.293 LAYER ME4 ;
END DO13
PIN DI12
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 53.082 0.000 53.402 0.600 ;
  LAYER ME3 ;
  RECT 53.082 0.000 53.402 0.600 ;
  LAYER ME2 ;
  RECT 53.082 0.000 53.402 0.600 ;
  LAYER ME1 ;
  RECT 53.082 0.000 53.402 0.600 ;
 END
 ANTENNAPARTIALMETALAREA                  1.058 LAYER ME2 ;
 ANTENNAGATEAREA                          0.072 LAYER ME2 ;
 ANTENNAGATEAREA                          0.072 LAYER ME3 ;
 ANTENNAGATEAREA                          0.072 LAYER ME4 ;
 ANTENNADIFFAREA                          0.160 LAYER ME2 ;
 ANTENNADIFFAREA                          0.160 LAYER ME3 ;
 ANTENNADIFFAREA                          0.160 LAYER ME4 ;
 ANTENNAMAXAREACAR                       21.782 LAYER ME2 ;
 ANTENNAMAXAREACAR                       24.449 LAYER ME3 ;
 ANTENNAMAXAREACAR                       27.116 LAYER ME4 ;
END DI12
PIN DO12
  DIRECTION OUTPUT ;
 PORT
  LAYER ME4 ;
  RECT 52.520 0.000 52.840 0.600 ;
  LAYER ME3 ;
  RECT 52.520 0.000 52.840 0.600 ;
  LAYER ME2 ;
  RECT 52.520 0.000 52.840 0.600 ;
  LAYER ME1 ;
  RECT 52.520 0.000 52.840 0.600 ;
 END
 ANTENNAPARTIALMETALAREA                  5.273 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME3 ;
 ANTENNADIFFAREA                          1.293 LAYER ME4 ;
END DO12
PIN DI11
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 48.516 0.000 48.836 0.600 ;
  LAYER ME3 ;
  RECT 48.516 0.000 48.836 0.600 ;
  LAYER ME2 ;
  RECT 48.516 0.000 48.836 0.600 ;
  LAYER ME1 ;
  RECT 48.516 0.000 48.836 0.600 ;
 END
 ANTENNAPARTIALMETALAREA                  0.346 LAYER ME1 ;
 ANTENNAPARTIALMETALAREA                  1.466 LAYER ME2 ;
 ANTENNAPARTIALMETALAREA                  0.508 LAYER ME3 ;
 ANTENNAGATEAREA                          0.072 LAYER ME3 ;
 ANTENNAGATEAREA                          0.072 LAYER ME4 ;
 ANTENNADIFFAREA                          0.218 LAYER ME1 ;
 ANTENNADIFFAREA                          0.218 LAYER ME2 ;
 ANTENNADIFFAREA                          0.218 LAYER ME3 ;
 ANTENNADIFFAREA                          0.218 LAYER ME4 ;
 ANTENNAMAXAREACAR                       17.267 LAYER ME3 ;
 ANTENNAMAXAREACAR                       19.933 LAYER ME4 ;
END DI11
PIN DO11
  DIRECTION OUTPUT ;
 PORT
  LAYER ME4 ;
  RECT 49.078 0.000 49.398 0.600 ;
  LAYER ME3 ;
  RECT 49.078 0.000 49.398 0.600 ;
  LAYER ME2 ;
  RECT 49.078 0.000 49.398 0.600 ;
  LAYER ME1 ;
  RECT 49.078 0.000 49.398 0.600 ;
 END
 ANTENNAPARTIALMETALAREA                  5.602 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME3 ;
 ANTENNADIFFAREA                          1.293 LAYER ME4 ;
END DO11
PIN WEB1
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 47.076 0.000 47.396 0.600 ;
  LAYER ME3 ;
  RECT 47.076 0.000 47.396 0.600 ;
  LAYER ME2 ;
  RECT 47.076 0.000 47.396 0.600 ;
  LAYER ME1 ;
  RECT 47.076 0.000 47.396 0.600 ;
 END
 ANTENNAPARTIALMETALAREA                  1.036 LAYER ME2 ;
 ANTENNAGATEAREA                          0.288 LAYER ME2 ;
 ANTENNAGATEAREA                          0.288 LAYER ME3 ;
 ANTENNAGATEAREA                          0.288 LAYER ME4 ;
 ANTENNADIFFAREA                          0.206 LAYER ME2 ;
 ANTENNADIFFAREA                          0.206 LAYER ME3 ;
 ANTENNADIFFAREA                          0.206 LAYER ME4 ;
 ANTENNAMAXAREACAR                        5.844 LAYER ME2 ;
 ANTENNAMAXAREACAR                        6.511 LAYER ME3 ;
 ANTENNAMAXAREACAR                        7.178 LAYER ME4 ;
END WEB1
PIN DI10
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 45.074 0.000 45.394 0.600 ;
  LAYER ME3 ;
  RECT 45.074 0.000 45.394 0.600 ;
  LAYER ME2 ;
  RECT 45.074 0.000 45.394 0.600 ;
  LAYER ME1 ;
  RECT 45.074 0.000 45.394 0.600 ;
 END
 ANTENNAPARTIALMETALAREA                  1.058 LAYER ME2 ;
 ANTENNAGATEAREA                          0.072 LAYER ME2 ;
 ANTENNAGATEAREA                          0.072 LAYER ME3 ;
 ANTENNAGATEAREA                          0.072 LAYER ME4 ;
 ANTENNADIFFAREA                          0.160 LAYER ME2 ;
 ANTENNADIFFAREA                          0.160 LAYER ME3 ;
 ANTENNADIFFAREA                          0.160 LAYER ME4 ;
 ANTENNAMAXAREACAR                       21.782 LAYER ME2 ;
 ANTENNAMAXAREACAR                       24.449 LAYER ME3 ;
 ANTENNAMAXAREACAR                       27.116 LAYER ME4 ;
END DI10
PIN DO10
  DIRECTION OUTPUT ;
 PORT
  LAYER ME4 ;
  RECT 44.512 0.000 44.832 0.600 ;
  LAYER ME3 ;
  RECT 44.512 0.000 44.832 0.600 ;
  LAYER ME2 ;
  RECT 44.512 0.000 44.832 0.600 ;
  LAYER ME1 ;
  RECT 44.512 0.000 44.832 0.600 ;
 END
 ANTENNAPARTIALMETALAREA                  5.273 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME3 ;
 ANTENNADIFFAREA                          1.293 LAYER ME4 ;
END DO10
PIN DI9
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 41.070 0.000 41.390 0.600 ;
  LAYER ME3 ;
  RECT 41.070 0.000 41.390 0.600 ;
  LAYER ME2 ;
  RECT 41.070 0.000 41.390 0.600 ;
  LAYER ME1 ;
  RECT 41.070 0.000 41.390 0.600 ;
 END
 ANTENNAPARTIALMETALAREA                  1.058 LAYER ME2 ;
 ANTENNAGATEAREA                          0.072 LAYER ME2 ;
 ANTENNAGATEAREA                          0.072 LAYER ME3 ;
 ANTENNAGATEAREA                          0.072 LAYER ME4 ;
 ANTENNADIFFAREA                          0.160 LAYER ME2 ;
 ANTENNADIFFAREA                          0.160 LAYER ME3 ;
 ANTENNADIFFAREA                          0.160 LAYER ME4 ;
 ANTENNAMAXAREACAR                       21.782 LAYER ME2 ;
 ANTENNAMAXAREACAR                       24.449 LAYER ME3 ;
 ANTENNAMAXAREACAR                       27.116 LAYER ME4 ;
END DI9
PIN DO9
  DIRECTION OUTPUT ;
 PORT
  LAYER ME4 ;
  RECT 40.508 0.000 40.828 0.600 ;
  LAYER ME3 ;
  RECT 40.508 0.000 40.828 0.600 ;
  LAYER ME2 ;
  RECT 40.508 0.000 40.828 0.600 ;
  LAYER ME1 ;
  RECT 40.508 0.000 40.828 0.600 ;
 END
 ANTENNAPARTIALMETALAREA                  5.273 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME3 ;
 ANTENNADIFFAREA                          1.293 LAYER ME4 ;
END DO9
PIN DI8
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 37.066 0.000 37.386 0.600 ;
  LAYER ME3 ;
  RECT 37.066 0.000 37.386 0.600 ;
  LAYER ME2 ;
  RECT 37.066 0.000 37.386 0.600 ;
  LAYER ME1 ;
  RECT 37.066 0.000 37.386 0.600 ;
 END
 ANTENNAPARTIALMETALAREA                  1.058 LAYER ME2 ;
 ANTENNAGATEAREA                          0.072 LAYER ME2 ;
 ANTENNAGATEAREA                          0.072 LAYER ME3 ;
 ANTENNAGATEAREA                          0.072 LAYER ME4 ;
 ANTENNADIFFAREA                          0.160 LAYER ME2 ;
 ANTENNADIFFAREA                          0.160 LAYER ME3 ;
 ANTENNADIFFAREA                          0.160 LAYER ME4 ;
 ANTENNAMAXAREACAR                       21.782 LAYER ME2 ;
 ANTENNAMAXAREACAR                       24.449 LAYER ME3 ;
 ANTENNAMAXAREACAR                       27.116 LAYER ME4 ;
END DI8
PIN DO8
  DIRECTION OUTPUT ;
 PORT
  LAYER ME4 ;
  RECT 36.504 0.000 36.824 0.600 ;
  LAYER ME3 ;
  RECT 36.504 0.000 36.824 0.600 ;
  LAYER ME2 ;
  RECT 36.504 0.000 36.824 0.600 ;
  LAYER ME1 ;
  RECT 36.504 0.000 36.824 0.600 ;
 END
 ANTENNAPARTIALMETALAREA                  5.273 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME3 ;
 ANTENNADIFFAREA                          1.293 LAYER ME4 ;
END DO8
PIN DI7
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 33.062 0.000 33.382 0.600 ;
  LAYER ME3 ;
  RECT 33.062 0.000 33.382 0.600 ;
  LAYER ME2 ;
  RECT 33.062 0.000 33.382 0.600 ;
  LAYER ME1 ;
  RECT 33.062 0.000 33.382 0.600 ;
 END
 ANTENNAPARTIALMETALAREA                  1.058 LAYER ME2 ;
 ANTENNAGATEAREA                          0.072 LAYER ME2 ;
 ANTENNAGATEAREA                          0.072 LAYER ME3 ;
 ANTENNAGATEAREA                          0.072 LAYER ME4 ;
 ANTENNADIFFAREA                          0.160 LAYER ME2 ;
 ANTENNADIFFAREA                          0.160 LAYER ME3 ;
 ANTENNADIFFAREA                          0.160 LAYER ME4 ;
 ANTENNAMAXAREACAR                       21.782 LAYER ME2 ;
 ANTENNAMAXAREACAR                       24.449 LAYER ME3 ;
 ANTENNAMAXAREACAR                       27.116 LAYER ME4 ;
END DI7
PIN DO7
  DIRECTION OUTPUT ;
 PORT
  LAYER ME4 ;
  RECT 32.500 0.000 32.820 0.600 ;
  LAYER ME3 ;
  RECT 32.500 0.000 32.820 0.600 ;
  LAYER ME2 ;
  RECT 32.500 0.000 32.820 0.600 ;
  LAYER ME1 ;
  RECT 32.500 0.000 32.820 0.600 ;
 END
 ANTENNAPARTIALMETALAREA                  5.273 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME3 ;
 ANTENNADIFFAREA                          1.293 LAYER ME4 ;
END DO7
PIN DI6
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 29.058 0.000 29.378 0.600 ;
  LAYER ME3 ;
  RECT 29.058 0.000 29.378 0.600 ;
  LAYER ME2 ;
  RECT 29.058 0.000 29.378 0.600 ;
  LAYER ME1 ;
  RECT 29.058 0.000 29.378 0.600 ;
 END
 ANTENNAPARTIALMETALAREA                  1.058 LAYER ME2 ;
 ANTENNAGATEAREA                          0.072 LAYER ME2 ;
 ANTENNAGATEAREA                          0.072 LAYER ME3 ;
 ANTENNAGATEAREA                          0.072 LAYER ME4 ;
 ANTENNADIFFAREA                          0.160 LAYER ME2 ;
 ANTENNADIFFAREA                          0.160 LAYER ME3 ;
 ANTENNADIFFAREA                          0.160 LAYER ME4 ;
 ANTENNAMAXAREACAR                       21.782 LAYER ME2 ;
 ANTENNAMAXAREACAR                       24.449 LAYER ME3 ;
 ANTENNAMAXAREACAR                       27.116 LAYER ME4 ;
END DI6
PIN DO6
  DIRECTION OUTPUT ;
 PORT
  LAYER ME4 ;
  RECT 28.496 0.000 28.816 0.600 ;
  LAYER ME3 ;
  RECT 28.496 0.000 28.816 0.600 ;
  LAYER ME2 ;
  RECT 28.496 0.000 28.816 0.600 ;
  LAYER ME1 ;
  RECT 28.496 0.000 28.816 0.600 ;
 END
 ANTENNAPARTIALMETALAREA                  5.273 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME3 ;
 ANTENNADIFFAREA                          1.293 LAYER ME4 ;
END DO6
PIN DI5
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 25.054 0.000 25.374 0.600 ;
  LAYER ME3 ;
  RECT 25.054 0.000 25.374 0.600 ;
  LAYER ME2 ;
  RECT 25.054 0.000 25.374 0.600 ;
  LAYER ME1 ;
  RECT 25.054 0.000 25.374 0.600 ;
 END
 ANTENNAPARTIALMETALAREA                  1.058 LAYER ME2 ;
 ANTENNAGATEAREA                          0.072 LAYER ME2 ;
 ANTENNAGATEAREA                          0.072 LAYER ME3 ;
 ANTENNAGATEAREA                          0.072 LAYER ME4 ;
 ANTENNADIFFAREA                          0.160 LAYER ME2 ;
 ANTENNADIFFAREA                          0.160 LAYER ME3 ;
 ANTENNADIFFAREA                          0.160 LAYER ME4 ;
 ANTENNAMAXAREACAR                       21.782 LAYER ME2 ;
 ANTENNAMAXAREACAR                       24.449 LAYER ME3 ;
 ANTENNAMAXAREACAR                       27.116 LAYER ME4 ;
END DI5
PIN DO5
  DIRECTION OUTPUT ;
 PORT
  LAYER ME4 ;
  RECT 24.492 0.000 24.812 0.600 ;
  LAYER ME3 ;
  RECT 24.492 0.000 24.812 0.600 ;
  LAYER ME2 ;
  RECT 24.492 0.000 24.812 0.600 ;
  LAYER ME1 ;
  RECT 24.492 0.000 24.812 0.600 ;
 END
 ANTENNAPARTIALMETALAREA                  5.273 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME3 ;
 ANTENNADIFFAREA                          1.293 LAYER ME4 ;
END DO5
PIN DI4
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 21.050 0.000 21.370 0.600 ;
  LAYER ME3 ;
  RECT 21.050 0.000 21.370 0.600 ;
  LAYER ME2 ;
  RECT 21.050 0.000 21.370 0.600 ;
  LAYER ME1 ;
  RECT 21.050 0.000 21.370 0.600 ;
 END
 ANTENNAPARTIALMETALAREA                  1.058 LAYER ME2 ;
 ANTENNAGATEAREA                          0.072 LAYER ME2 ;
 ANTENNAGATEAREA                          0.072 LAYER ME3 ;
 ANTENNAGATEAREA                          0.072 LAYER ME4 ;
 ANTENNADIFFAREA                          0.160 LAYER ME2 ;
 ANTENNADIFFAREA                          0.160 LAYER ME3 ;
 ANTENNADIFFAREA                          0.160 LAYER ME4 ;
 ANTENNAMAXAREACAR                       21.782 LAYER ME2 ;
 ANTENNAMAXAREACAR                       24.449 LAYER ME3 ;
 ANTENNAMAXAREACAR                       27.116 LAYER ME4 ;
END DI4
PIN DO4
  DIRECTION OUTPUT ;
 PORT
  LAYER ME4 ;
  RECT 20.488 0.000 20.808 0.600 ;
  LAYER ME3 ;
  RECT 20.488 0.000 20.808 0.600 ;
  LAYER ME2 ;
  RECT 20.488 0.000 20.808 0.600 ;
  LAYER ME1 ;
  RECT 20.488 0.000 20.808 0.600 ;
 END
 ANTENNAPARTIALMETALAREA                  5.273 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME3 ;
 ANTENNADIFFAREA                          1.293 LAYER ME4 ;
END DO4
PIN DI3
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 17.046 0.000 17.366 0.600 ;
  LAYER ME3 ;
  RECT 17.046 0.000 17.366 0.600 ;
  LAYER ME2 ;
  RECT 17.046 0.000 17.366 0.600 ;
  LAYER ME1 ;
  RECT 17.046 0.000 17.366 0.600 ;
 END
 ANTENNAPARTIALMETALAREA                  1.058 LAYER ME2 ;
 ANTENNAGATEAREA                          0.072 LAYER ME2 ;
 ANTENNAGATEAREA                          0.072 LAYER ME3 ;
 ANTENNAGATEAREA                          0.072 LAYER ME4 ;
 ANTENNADIFFAREA                          0.160 LAYER ME2 ;
 ANTENNADIFFAREA                          0.160 LAYER ME3 ;
 ANTENNADIFFAREA                          0.160 LAYER ME4 ;
 ANTENNAMAXAREACAR                       21.782 LAYER ME2 ;
 ANTENNAMAXAREACAR                       24.449 LAYER ME3 ;
 ANTENNAMAXAREACAR                       27.116 LAYER ME4 ;
END DI3
PIN DO3
  DIRECTION OUTPUT ;
 PORT
  LAYER ME4 ;
  RECT 16.484 0.000 16.804 0.600 ;
  LAYER ME3 ;
  RECT 16.484 0.000 16.804 0.600 ;
  LAYER ME2 ;
  RECT 16.484 0.000 16.804 0.600 ;
  LAYER ME1 ;
  RECT 16.484 0.000 16.804 0.600 ;
 END
 ANTENNAPARTIALMETALAREA                  5.273 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME3 ;
 ANTENNADIFFAREA                          1.293 LAYER ME4 ;
END DO3
PIN DI2
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 13.042 0.000 13.362 0.600 ;
  LAYER ME3 ;
  RECT 13.042 0.000 13.362 0.600 ;
  LAYER ME2 ;
  RECT 13.042 0.000 13.362 0.600 ;
  LAYER ME1 ;
  RECT 13.042 0.000 13.362 0.600 ;
 END
 ANTENNAPARTIALMETALAREA                  1.058 LAYER ME2 ;
 ANTENNAGATEAREA                          0.072 LAYER ME2 ;
 ANTENNAGATEAREA                          0.072 LAYER ME3 ;
 ANTENNAGATEAREA                          0.072 LAYER ME4 ;
 ANTENNADIFFAREA                          0.160 LAYER ME2 ;
 ANTENNADIFFAREA                          0.160 LAYER ME3 ;
 ANTENNADIFFAREA                          0.160 LAYER ME4 ;
 ANTENNAMAXAREACAR                       21.782 LAYER ME2 ;
 ANTENNAMAXAREACAR                       24.449 LAYER ME3 ;
 ANTENNAMAXAREACAR                       27.116 LAYER ME4 ;
END DI2
PIN DO2
  DIRECTION OUTPUT ;
 PORT
  LAYER ME4 ;
  RECT 12.480 0.000 12.800 0.600 ;
  LAYER ME3 ;
  RECT 12.480 0.000 12.800 0.600 ;
  LAYER ME2 ;
  RECT 12.480 0.000 12.800 0.600 ;
  LAYER ME1 ;
  RECT 12.480 0.000 12.800 0.600 ;
 END
 ANTENNAPARTIALMETALAREA                  5.273 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME3 ;
 ANTENNADIFFAREA                          1.293 LAYER ME4 ;
END DO2
PIN DI1
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 9.038 0.000 9.358 0.600 ;
  LAYER ME3 ;
  RECT 9.038 0.000 9.358 0.600 ;
  LAYER ME2 ;
  RECT 9.038 0.000 9.358 0.600 ;
  LAYER ME1 ;
  RECT 9.038 0.000 9.358 0.600 ;
 END
 ANTENNAPARTIALMETALAREA                  1.058 LAYER ME2 ;
 ANTENNAGATEAREA                          0.072 LAYER ME2 ;
 ANTENNAGATEAREA                          0.072 LAYER ME3 ;
 ANTENNAGATEAREA                          0.072 LAYER ME4 ;
 ANTENNADIFFAREA                          0.160 LAYER ME2 ;
 ANTENNADIFFAREA                          0.160 LAYER ME3 ;
 ANTENNADIFFAREA                          0.160 LAYER ME4 ;
 ANTENNAMAXAREACAR                       21.782 LAYER ME2 ;
 ANTENNAMAXAREACAR                       24.449 LAYER ME3 ;
 ANTENNAMAXAREACAR                       27.116 LAYER ME4 ;
END DI1
PIN DO1
  DIRECTION OUTPUT ;
 PORT
  LAYER ME4 ;
  RECT 8.476 0.000 8.796 0.600 ;
  LAYER ME3 ;
  RECT 8.476 0.000 8.796 0.600 ;
  LAYER ME2 ;
  RECT 8.476 0.000 8.796 0.600 ;
  LAYER ME1 ;
  RECT 8.476 0.000 8.796 0.600 ;
 END
 ANTENNAPARTIALMETALAREA                  5.273 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME3 ;
 ANTENNADIFFAREA                          1.293 LAYER ME4 ;
END DO1
PIN DI0
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 4.472 0.000 4.792 0.600 ;
  LAYER ME3 ;
  RECT 4.472 0.000 4.792 0.600 ;
  LAYER ME2 ;
  RECT 4.472 0.000 4.792 0.600 ;
  LAYER ME1 ;
  RECT 4.472 0.000 4.792 0.600 ;
 END
 ANTENNAPARTIALMETALAREA                  0.346 LAYER ME1 ;
 ANTENNAPARTIALMETALAREA                  1.466 LAYER ME2 ;
 ANTENNAPARTIALMETALAREA                  0.508 LAYER ME3 ;
 ANTENNAGATEAREA                          0.072 LAYER ME3 ;
 ANTENNAGATEAREA                          0.072 LAYER ME4 ;
 ANTENNADIFFAREA                          0.218 LAYER ME1 ;
 ANTENNADIFFAREA                          0.218 LAYER ME2 ;
 ANTENNADIFFAREA                          0.218 LAYER ME3 ;
 ANTENNADIFFAREA                          0.218 LAYER ME4 ;
 ANTENNAMAXAREACAR                       17.267 LAYER ME3 ;
 ANTENNAMAXAREACAR                       19.933 LAYER ME4 ;
END DI0
PIN DO0
  DIRECTION OUTPUT ;
 PORT
  LAYER ME4 ;
  RECT 5.034 0.000 5.354 0.600 ;
  LAYER ME3 ;
  RECT 5.034 0.000 5.354 0.600 ;
  LAYER ME2 ;
  RECT 5.034 0.000 5.354 0.600 ;
  LAYER ME1 ;
  RECT 5.034 0.000 5.354 0.600 ;
 END
 ANTENNAPARTIALMETALAREA                  5.602 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME3 ;
 ANTENNADIFFAREA                          1.293 LAYER ME4 ;
END DO0
PIN WEB0
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 3.032 0.000 3.352 0.600 ;
  LAYER ME3 ;
  RECT 3.032 0.000 3.352 0.600 ;
  LAYER ME2 ;
  RECT 3.032 0.000 3.352 0.600 ;
  LAYER ME1 ;
  RECT 3.032 0.000 3.352 0.600 ;
 END
 ANTENNAPARTIALMETALAREA                  1.036 LAYER ME2 ;
 ANTENNAGATEAREA                          0.288 LAYER ME2 ;
 ANTENNAGATEAREA                          0.288 LAYER ME3 ;
 ANTENNAGATEAREA                          0.288 LAYER ME4 ;
 ANTENNADIFFAREA                          0.206 LAYER ME2 ;
 ANTENNADIFFAREA                          0.206 LAYER ME3 ;
 ANTENNADIFFAREA                          0.206 LAYER ME4 ;
 ANTENNAMAXAREACAR                        5.844 LAYER ME2 ;
 ANTENNAMAXAREACAR                        6.511 LAYER ME3 ;
 ANTENNAMAXAREACAR                        7.178 LAYER ME4 ;
END WEB0
PIN A1
  DIRECTION INPUT ;
 PORT
  LAYER ME3 ;
  RECT 106.968 0.000 107.288 0.720 ;
  LAYER ME2 ;
  RECT 106.968 0.000 107.288 0.720 ;
  LAYER ME1 ;
  RECT 106.968 0.000 107.288 0.720 ;
 END
 ANTENNAPARTIALMETALAREA                  3.547 LAYER ME2 ;
 ANTENNAGATEAREA                          0.144 LAYER ME2 ;
 ANTENNAGATEAREA                          0.144 LAYER ME3 ;
 ANTENNADIFFAREA                          0.218 LAYER ME2 ;
 ANTENNADIFFAREA                          0.218 LAYER ME3 ;
 ANTENNAMAXAREACAR                       27.235 LAYER ME2 ;
 ANTENNAMAXAREACAR                       28.835 LAYER ME3 ;
END A1
PIN A2
  DIRECTION INPUT ;
 PORT
  LAYER ME3 ;
  RECT 107.538 0.000 107.858 0.720 ;
  LAYER ME2 ;
  RECT 107.538 0.000 107.858 0.720 ;
  LAYER ME1 ;
  RECT 107.538 0.000 107.858 0.720 ;
 END
 ANTENNAPARTIALMETALAREA                  3.688 LAYER ME2 ;
 ANTENNAGATEAREA                          0.144 LAYER ME2 ;
 ANTENNAGATEAREA                          0.144 LAYER ME3 ;
 ANTENNADIFFAREA                          0.218 LAYER ME2 ;
 ANTENNADIFFAREA                          0.218 LAYER ME3 ;
 ANTENNAMAXAREACAR                       28.214 LAYER ME2 ;
 ANTENNAMAXAREACAR                       29.814 LAYER ME3 ;
END A2
PIN A3
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 100.720 0.000 101.040 0.720 ;
  LAYER ME3 ;
  RECT 100.720 0.000 101.040 0.720 ;
  LAYER ME2 ;
  RECT 100.720 0.000 101.040 0.720 ;
  LAYER ME1 ;
  RECT 100.720 0.000 101.040 0.720 ;
 END
 ANTENNAPARTIALMETALAREA                  4.391 LAYER ME2 ;
 ANTENNAGATEAREA                          0.180 LAYER ME2 ;
 ANTENNAGATEAREA                          0.180 LAYER ME3 ;
 ANTENNAGATEAREA                          0.180 LAYER ME4 ;
 ANTENNADIFFAREA                          0.218 LAYER ME2 ;
 ANTENNADIFFAREA                          0.218 LAYER ME3 ;
 ANTENNADIFFAREA                          0.218 LAYER ME4 ;
 ANTENNAMAXAREACAR                       27.451 LAYER ME2 ;
 ANTENNAMAXAREACAR                       28.731 LAYER ME3 ;
 ANTENNAMAXAREACAR                       30.011 LAYER ME4 ;
END A3
PIN A4
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 100.040 0.000 100.360 0.720 ;
  LAYER ME3 ;
  RECT 100.040 0.000 100.360 0.720 ;
  LAYER ME2 ;
  RECT 100.040 0.000 100.360 0.720 ;
  LAYER ME1 ;
  RECT 100.040 0.000 100.360 0.720 ;
 END
 ANTENNAPARTIALMETALAREA                  3.928 LAYER ME2 ;
 ANTENNAGATEAREA                          0.180 LAYER ME2 ;
 ANTENNAGATEAREA                          0.180 LAYER ME3 ;
 ANTENNAGATEAREA                          0.180 LAYER ME4 ;
 ANTENNADIFFAREA                          0.218 LAYER ME2 ;
 ANTENNADIFFAREA                          0.218 LAYER ME3 ;
 ANTENNADIFFAREA                          0.218 LAYER ME4 ;
 ANTENNAMAXAREACAR                       26.813 LAYER ME2 ;
 ANTENNAMAXAREACAR                       28.093 LAYER ME3 ;
 ANTENNAMAXAREACAR                       29.373 LAYER ME4 ;
END A4
PIN A5
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 96.560 0.000 96.880 0.720 ;
  LAYER ME3 ;
  RECT 96.560 0.000 96.880 0.720 ;
  LAYER ME2 ;
  RECT 96.560 0.000 96.880 0.720 ;
  LAYER ME1 ;
  RECT 96.560 0.000 96.880 0.720 ;
 END
 ANTENNAPARTIALMETALAREA                  4.391 LAYER ME2 ;
 ANTENNAGATEAREA                          0.180 LAYER ME2 ;
 ANTENNAGATEAREA                          0.180 LAYER ME3 ;
 ANTENNAGATEAREA                          0.180 LAYER ME4 ;
 ANTENNADIFFAREA                          0.218 LAYER ME2 ;
 ANTENNADIFFAREA                          0.218 LAYER ME3 ;
 ANTENNADIFFAREA                          0.218 LAYER ME4 ;
 ANTENNAMAXAREACAR                       27.451 LAYER ME2 ;
 ANTENNAMAXAREACAR                       28.731 LAYER ME3 ;
 ANTENNAMAXAREACAR                       30.011 LAYER ME4 ;
END A5
PIN A6
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 95.880 0.000 96.200 0.720 ;
  LAYER ME3 ;
  RECT 95.880 0.000 96.200 0.720 ;
  LAYER ME2 ;
  RECT 95.880 0.000 96.200 0.720 ;
  LAYER ME1 ;
  RECT 95.880 0.000 96.200 0.720 ;
 END
 ANTENNAPARTIALMETALAREA                  3.928 LAYER ME2 ;
 ANTENNAGATEAREA                          0.180 LAYER ME2 ;
 ANTENNAGATEAREA                          0.180 LAYER ME3 ;
 ANTENNAGATEAREA                          0.180 LAYER ME4 ;
 ANTENNADIFFAREA                          0.218 LAYER ME2 ;
 ANTENNADIFFAREA                          0.218 LAYER ME3 ;
 ANTENNADIFFAREA                          0.218 LAYER ME4 ;
 ANTENNAMAXAREACAR                       26.813 LAYER ME2 ;
 ANTENNAMAXAREACAR                       28.093 LAYER ME3 ;
 ANTENNAMAXAREACAR                       29.373 LAYER ME4 ;
END A6
PIN A0
  DIRECTION INPUT ;
 PORT
  LAYER ME3 ;
  RECT 117.554 0.000 117.874 0.662 ;
  LAYER ME2 ;
  RECT 117.554 0.000 117.874 0.662 ;
  LAYER ME1 ;
  RECT 117.554 0.000 117.874 0.662 ;
 END
 ANTENNAPARTIALMETALAREA                  5.907 LAYER ME2 ;
 ANTENNAGATEAREA                          0.108 LAYER ME2 ;
 ANTENNAGATEAREA                          0.108 LAYER ME3 ;
 ANTENNADIFFAREA                          0.218 LAYER ME2 ;
 ANTENNADIFFAREA                          0.218 LAYER ME3 ;
 ANTENNAMAXAREACAR                       58.521 LAYER ME2 ;
 ANTENNAMAXAREACAR                       60.482 LAYER ME3 ;
END A0
PIN DVSE
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 127.145 0.000 127.465 0.720 ;
  LAYER ME3 ;
  RECT 127.145 0.000 127.465 0.720 ;
  LAYER ME3 ;
  RECT 127.145 0.000 127.465 0.720 ;
  LAYER ME2 ;
  RECT 127.145 0.000 127.465 0.720 ;
  LAYER ME2 ;
  RECT 127.145 0.000 127.465 0.720 ;
  LAYER ME1 ;
  RECT 127.145 0.000 127.465 0.720 ;
  LAYER ME1 ;
  RECT 127.145 0.000 127.465 0.720 ;
 END
 ANTENNAPARTIALMETALAREA                  7.809 LAYER ME2 ;
 ANTENNAGATEAREA                          0.612 LAYER ME2 ;
 ANTENNAGATEAREA                          0.612 LAYER ME3 ;
 ANTENNAGATEAREA                          0.612 LAYER ME4 ;
 ANTENNADIFFAREA                          0.218 LAYER ME2 ;
 ANTENNADIFFAREA                          0.218 LAYER ME3 ;
 ANTENNADIFFAREA                          0.218 LAYER ME4 ;
 ANTENNAMAXAREACAR                       76.330 LAYER ME2 ;
 ANTENNAMAXAREACAR                       78.463 LAYER ME3 ;
 ANTENNAMAXAREACAR                       80.596 LAYER ME4 ;
END DVSE
PIN DVS3
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 126.625 0.000 126.945 0.720 ;
  LAYER ME3 ;
  RECT 126.625 0.000 126.945 0.720 ;
  LAYER ME3 ;
  RECT 126.625 0.000 126.945 0.720 ;
  LAYER ME2 ;
  RECT 126.625 0.000 126.945 0.720 ;
  LAYER ME2 ;
  RECT 126.625 0.000 126.945 0.720 ;
  LAYER ME1 ;
  RECT 126.625 0.000 126.945 0.720 ;
  LAYER ME1 ;
  RECT 126.625 0.000 126.945 0.720 ;
 END
 ANTENNAPARTIALMETALAREA                  6.179 LAYER ME2 ;
 ANTENNAGATEAREA                          0.108 LAYER ME2 ;
 ANTENNAGATEAREA                          0.108 LAYER ME3 ;
 ANTENNAGATEAREA                          0.108 LAYER ME4 ;
 ANTENNADIFFAREA                          0.218 LAYER ME2 ;
 ANTENNADIFFAREA                          0.218 LAYER ME3 ;
 ANTENNADIFFAREA                          0.218 LAYER ME4 ;
 ANTENNAMAXAREACAR                       68.823 LAYER ME2 ;
 ANTENNAMAXAREACAR                       70.956 LAYER ME3 ;
 ANTENNAMAXAREACAR                       73.089 LAYER ME4 ;
END DVS3
PIN DVS2
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 127.665 0.000 127.985 0.720 ;
  LAYER ME3 ;
  RECT 127.665 0.000 127.985 0.720 ;
  LAYER ME3 ;
  RECT 127.665 0.000 127.985 0.720 ;
  LAYER ME2 ;
  RECT 127.665 0.000 127.985 0.720 ;
  LAYER ME2 ;
  RECT 127.665 0.000 127.985 0.720 ;
  LAYER ME1 ;
  RECT 127.665 0.000 127.985 0.720 ;
  LAYER ME1 ;
  RECT 127.665 0.000 127.985 0.720 ;
 END
 ANTENNAPARTIALMETALAREA                  7.876 LAYER ME2 ;
 ANTENNAGATEAREA                          0.108 LAYER ME2 ;
 ANTENNAGATEAREA                          0.108 LAYER ME3 ;
 ANTENNAGATEAREA                          0.108 LAYER ME4 ;
 ANTENNADIFFAREA                          0.218 LAYER ME2 ;
 ANTENNADIFFAREA                          0.218 LAYER ME3 ;
 ANTENNADIFFAREA                          0.218 LAYER ME4 ;
 ANTENNAMAXAREACAR                       83.257 LAYER ME2 ;
 ANTENNAMAXAREACAR                       85.391 LAYER ME3 ;
 ANTENNAMAXAREACAR                       87.524 LAYER ME4 ;
END DVS2
PIN DVS1
  DIRECTION INPUT ;
 PORT
  LAYER ME3 ;
  RECT 124.009 0.000 124.329 0.720 ;
  LAYER ME2 ;
  RECT 124.009 0.000 124.329 0.720 ;
  LAYER ME1 ;
  RECT 124.009 0.000 124.329 0.720 ;
 END
 ANTENNAPARTIALMETALAREA                  6.247 LAYER ME2 ;
 ANTENNAGATEAREA                          0.108 LAYER ME2 ;
 ANTENNAGATEAREA                          0.108 LAYER ME3 ;
 ANTENNADIFFAREA                          0.218 LAYER ME2 ;
 ANTENNADIFFAREA                          0.218 LAYER ME3 ;
 ANTENNAMAXAREACAR                       69.294 LAYER ME2 ;
 ANTENNAMAXAREACAR                       71.427 LAYER ME3 ;
END DVS1
PIN DVS0
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 128.185 0.000 128.505 0.720 ;
  LAYER ME3 ;
  RECT 128.185 0.000 128.505 0.720 ;
  LAYER ME3 ;
  RECT 128.185 0.000 128.505 0.720 ;
  LAYER ME2 ;
  RECT 128.185 0.000 128.505 0.720 ;
  LAYER ME2 ;
  RECT 128.185 0.000 128.505 0.720 ;
  LAYER ME1 ;
  RECT 128.185 0.000 128.505 0.720 ;
  LAYER ME1 ;
  RECT 128.185 0.000 128.505 0.720 ;
 END
 ANTENNAPARTIALMETALAREA                  7.119 LAYER ME2 ;
 ANTENNAGATEAREA                          0.108 LAYER ME2 ;
 ANTENNAGATEAREA                          0.108 LAYER ME3 ;
 ANTENNAGATEAREA                          0.108 LAYER ME4 ;
 ANTENNADIFFAREA                          0.218 LAYER ME2 ;
 ANTENNADIFFAREA                          0.218 LAYER ME3 ;
 ANTENNADIFFAREA                          0.218 LAYER ME4 ;
 ANTENNAMAXAREACAR                       77.987 LAYER ME2 ;
 ANTENNAMAXAREACAR                       80.120 LAYER ME3 ;
 ANTENNAMAXAREACAR                       82.254 LAYER ME4 ;
END DVS0
PIN CK
  DIRECTION INPUT ;
 PORT
  LAYER ME3 ;
  RECT 120.093 0.000 120.413 0.720 ;
  LAYER ME2 ;
  RECT 120.093 0.000 120.413 0.720 ;
  LAYER ME1 ;
  RECT 120.093 0.000 120.413 0.720 ;
 END
 ANTENNAPARTIALMETALAREA                  5.257 LAYER ME2 ;
 ANTENNAPARTIALMETALAREA                  7.044 LAYER ME3 ;
 ANTENNAGATEAREA                          0.072 LAYER ME2 ;
 ANTENNAGATEAREA                          1.044 LAYER ME3 ;
 ANTENNADIFFAREA                          0.218 LAYER ME2 ;
 ANTENNADIFFAREA                          0.218 LAYER ME3 ;
 ANTENNAMAXAREACAR                       86.308 LAYER ME2 ;
 ANTENNAMAXAREACAR                      187.347 LAYER ME3 ;
END CK
PIN CSB
  DIRECTION INPUT ;
 PORT
  LAYER ME3 ;
  RECT 111.479 0.000 111.799 0.720 ;
  LAYER ME2 ;
  RECT 111.479 0.000 111.799 0.720 ;
  LAYER ME1 ;
  RECT 111.479 0.000 111.799 0.720 ;
 END
 ANTENNAPARTIALMETALAREA                  5.788 LAYER ME2 ;
 ANTENNAPARTIALMETALAREA                  7.100 LAYER ME3 ;
 ANTENNAGATEAREA                          2.508 LAYER ME2 ;
 ANTENNAGATEAREA                          3.480 LAYER ME3 ;
 ANTENNADIFFAREA                          0.218 LAYER ME2 ;
 ANTENNADIFFAREA                          0.218 LAYER ME3 ;
 ANTENNAMAXAREACAR                        3.046 LAYER ME2 ;
 ANTENNAMAXAREACAR                       36.487 LAYER ME3 ;
END CSB
PIN DI43
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 214.883 0.000 215.203 0.600 ;
  LAYER ME3 ;
  RECT 214.883 0.000 215.203 0.600 ;
  LAYER ME2 ;
  RECT 214.883 0.000 215.203 0.600 ;
  LAYER ME1 ;
  RECT 214.883 0.000 215.203 0.600 ;
 END
 ANTENNAPARTIALMETALAREA                  1.058 LAYER ME2 ;
 ANTENNAGATEAREA                          0.072 LAYER ME2 ;
 ANTENNAGATEAREA                          0.072 LAYER ME3 ;
 ANTENNAGATEAREA                          0.072 LAYER ME4 ;
 ANTENNADIFFAREA                          0.160 LAYER ME2 ;
 ANTENNADIFFAREA                          0.160 LAYER ME3 ;
 ANTENNADIFFAREA                          0.160 LAYER ME4 ;
 ANTENNAMAXAREACAR                       21.782 LAYER ME2 ;
 ANTENNAMAXAREACAR                       24.449 LAYER ME3 ;
 ANTENNAMAXAREACAR                       27.116 LAYER ME4 ;
END DI43
PIN DO43
  DIRECTION OUTPUT ;
 PORT
  LAYER ME4 ;
  RECT 214.321 0.000 214.641 0.600 ;
  LAYER ME3 ;
  RECT 214.321 0.000 214.641 0.600 ;
  LAYER ME2 ;
  RECT 214.321 0.000 214.641 0.600 ;
  LAYER ME1 ;
  RECT 214.321 0.000 214.641 0.600 ;
 END
 ANTENNAPARTIALMETALAREA                  5.273 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME3 ;
 ANTENNADIFFAREA                          1.293 LAYER ME4 ;
END DO43
PIN DI42
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 210.879 0.000 211.199 0.600 ;
  LAYER ME3 ;
  RECT 210.879 0.000 211.199 0.600 ;
  LAYER ME2 ;
  RECT 210.879 0.000 211.199 0.600 ;
  LAYER ME1 ;
  RECT 210.879 0.000 211.199 0.600 ;
 END
 ANTENNAPARTIALMETALAREA                  1.058 LAYER ME2 ;
 ANTENNAGATEAREA                          0.072 LAYER ME2 ;
 ANTENNAGATEAREA                          0.072 LAYER ME3 ;
 ANTENNAGATEAREA                          0.072 LAYER ME4 ;
 ANTENNADIFFAREA                          0.160 LAYER ME2 ;
 ANTENNADIFFAREA                          0.160 LAYER ME3 ;
 ANTENNADIFFAREA                          0.160 LAYER ME4 ;
 ANTENNAMAXAREACAR                       21.782 LAYER ME2 ;
 ANTENNAMAXAREACAR                       24.449 LAYER ME3 ;
 ANTENNAMAXAREACAR                       27.116 LAYER ME4 ;
END DI42
PIN DO42
  DIRECTION OUTPUT ;
 PORT
  LAYER ME4 ;
  RECT 210.317 0.000 210.637 0.600 ;
  LAYER ME3 ;
  RECT 210.317 0.000 210.637 0.600 ;
  LAYER ME2 ;
  RECT 210.317 0.000 210.637 0.600 ;
  LAYER ME1 ;
  RECT 210.317 0.000 210.637 0.600 ;
 END
 ANTENNAPARTIALMETALAREA                  5.273 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME3 ;
 ANTENNADIFFAREA                          1.293 LAYER ME4 ;
END DO42
PIN DI41
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 206.875 0.000 207.195 0.600 ;
  LAYER ME3 ;
  RECT 206.875 0.000 207.195 0.600 ;
  LAYER ME2 ;
  RECT 206.875 0.000 207.195 0.600 ;
  LAYER ME1 ;
  RECT 206.875 0.000 207.195 0.600 ;
 END
 ANTENNAPARTIALMETALAREA                  1.058 LAYER ME2 ;
 ANTENNAGATEAREA                          0.072 LAYER ME2 ;
 ANTENNAGATEAREA                          0.072 LAYER ME3 ;
 ANTENNAGATEAREA                          0.072 LAYER ME4 ;
 ANTENNADIFFAREA                          0.160 LAYER ME2 ;
 ANTENNADIFFAREA                          0.160 LAYER ME3 ;
 ANTENNADIFFAREA                          0.160 LAYER ME4 ;
 ANTENNAMAXAREACAR                       21.782 LAYER ME2 ;
 ANTENNAMAXAREACAR                       24.449 LAYER ME3 ;
 ANTENNAMAXAREACAR                       27.116 LAYER ME4 ;
END DI41
PIN DO41
  DIRECTION OUTPUT ;
 PORT
  LAYER ME4 ;
  RECT 206.313 0.000 206.633 0.600 ;
  LAYER ME3 ;
  RECT 206.313 0.000 206.633 0.600 ;
  LAYER ME2 ;
  RECT 206.313 0.000 206.633 0.600 ;
  LAYER ME1 ;
  RECT 206.313 0.000 206.633 0.600 ;
 END
 ANTENNAPARTIALMETALAREA                  5.273 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME3 ;
 ANTENNADIFFAREA                          1.293 LAYER ME4 ;
END DO41
PIN DI40
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 202.871 0.000 203.191 0.600 ;
  LAYER ME3 ;
  RECT 202.871 0.000 203.191 0.600 ;
  LAYER ME2 ;
  RECT 202.871 0.000 203.191 0.600 ;
  LAYER ME1 ;
  RECT 202.871 0.000 203.191 0.600 ;
 END
 ANTENNAPARTIALMETALAREA                  1.058 LAYER ME2 ;
 ANTENNAGATEAREA                          0.072 LAYER ME2 ;
 ANTENNAGATEAREA                          0.072 LAYER ME3 ;
 ANTENNAGATEAREA                          0.072 LAYER ME4 ;
 ANTENNADIFFAREA                          0.160 LAYER ME2 ;
 ANTENNADIFFAREA                          0.160 LAYER ME3 ;
 ANTENNADIFFAREA                          0.160 LAYER ME4 ;
 ANTENNAMAXAREACAR                       21.782 LAYER ME2 ;
 ANTENNAMAXAREACAR                       24.449 LAYER ME3 ;
 ANTENNAMAXAREACAR                       27.116 LAYER ME4 ;
END DI40
PIN DO40
  DIRECTION OUTPUT ;
 PORT
  LAYER ME4 ;
  RECT 202.309 0.000 202.629 0.600 ;
  LAYER ME3 ;
  RECT 202.309 0.000 202.629 0.600 ;
  LAYER ME2 ;
  RECT 202.309 0.000 202.629 0.600 ;
  LAYER ME1 ;
  RECT 202.309 0.000 202.629 0.600 ;
 END
 ANTENNAPARTIALMETALAREA                  5.273 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME3 ;
 ANTENNADIFFAREA                          1.293 LAYER ME4 ;
END DO40
PIN DI39
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 198.867 0.000 199.187 0.600 ;
  LAYER ME3 ;
  RECT 198.867 0.000 199.187 0.600 ;
  LAYER ME2 ;
  RECT 198.867 0.000 199.187 0.600 ;
  LAYER ME1 ;
  RECT 198.867 0.000 199.187 0.600 ;
 END
 ANTENNAPARTIALMETALAREA                  1.058 LAYER ME2 ;
 ANTENNAGATEAREA                          0.072 LAYER ME2 ;
 ANTENNAGATEAREA                          0.072 LAYER ME3 ;
 ANTENNAGATEAREA                          0.072 LAYER ME4 ;
 ANTENNADIFFAREA                          0.160 LAYER ME2 ;
 ANTENNADIFFAREA                          0.160 LAYER ME3 ;
 ANTENNADIFFAREA                          0.160 LAYER ME4 ;
 ANTENNAMAXAREACAR                       21.782 LAYER ME2 ;
 ANTENNAMAXAREACAR                       24.449 LAYER ME3 ;
 ANTENNAMAXAREACAR                       27.116 LAYER ME4 ;
END DI39
PIN DO39
  DIRECTION OUTPUT ;
 PORT
  LAYER ME4 ;
  RECT 198.305 0.000 198.625 0.600 ;
  LAYER ME3 ;
  RECT 198.305 0.000 198.625 0.600 ;
  LAYER ME2 ;
  RECT 198.305 0.000 198.625 0.600 ;
  LAYER ME1 ;
  RECT 198.305 0.000 198.625 0.600 ;
 END
 ANTENNAPARTIALMETALAREA                  5.273 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME3 ;
 ANTENNADIFFAREA                          1.293 LAYER ME4 ;
END DO39
PIN DI38
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 194.863 0.000 195.183 0.600 ;
  LAYER ME3 ;
  RECT 194.863 0.000 195.183 0.600 ;
  LAYER ME2 ;
  RECT 194.863 0.000 195.183 0.600 ;
  LAYER ME1 ;
  RECT 194.863 0.000 195.183 0.600 ;
 END
 ANTENNAPARTIALMETALAREA                  1.058 LAYER ME2 ;
 ANTENNAGATEAREA                          0.072 LAYER ME2 ;
 ANTENNAGATEAREA                          0.072 LAYER ME3 ;
 ANTENNAGATEAREA                          0.072 LAYER ME4 ;
 ANTENNADIFFAREA                          0.160 LAYER ME2 ;
 ANTENNADIFFAREA                          0.160 LAYER ME3 ;
 ANTENNADIFFAREA                          0.160 LAYER ME4 ;
 ANTENNAMAXAREACAR                       21.782 LAYER ME2 ;
 ANTENNAMAXAREACAR                       24.449 LAYER ME3 ;
 ANTENNAMAXAREACAR                       27.116 LAYER ME4 ;
END DI38
PIN DO38
  DIRECTION OUTPUT ;
 PORT
  LAYER ME4 ;
  RECT 194.301 0.000 194.621 0.600 ;
  LAYER ME3 ;
  RECT 194.301 0.000 194.621 0.600 ;
  LAYER ME2 ;
  RECT 194.301 0.000 194.621 0.600 ;
  LAYER ME1 ;
  RECT 194.301 0.000 194.621 0.600 ;
 END
 ANTENNAPARTIALMETALAREA                  5.273 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME3 ;
 ANTENNADIFFAREA                          1.293 LAYER ME4 ;
END DO38
PIN DI37
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 190.859 0.000 191.179 0.600 ;
  LAYER ME3 ;
  RECT 190.859 0.000 191.179 0.600 ;
  LAYER ME2 ;
  RECT 190.859 0.000 191.179 0.600 ;
  LAYER ME1 ;
  RECT 190.859 0.000 191.179 0.600 ;
 END
 ANTENNAPARTIALMETALAREA                  1.058 LAYER ME2 ;
 ANTENNAGATEAREA                          0.072 LAYER ME2 ;
 ANTENNAGATEAREA                          0.072 LAYER ME3 ;
 ANTENNAGATEAREA                          0.072 LAYER ME4 ;
 ANTENNADIFFAREA                          0.160 LAYER ME2 ;
 ANTENNADIFFAREA                          0.160 LAYER ME3 ;
 ANTENNADIFFAREA                          0.160 LAYER ME4 ;
 ANTENNAMAXAREACAR                       21.782 LAYER ME2 ;
 ANTENNAMAXAREACAR                       24.449 LAYER ME3 ;
 ANTENNAMAXAREACAR                       27.116 LAYER ME4 ;
END DI37
PIN DO37
  DIRECTION OUTPUT ;
 PORT
  LAYER ME4 ;
  RECT 190.297 0.000 190.617 0.600 ;
  LAYER ME3 ;
  RECT 190.297 0.000 190.617 0.600 ;
  LAYER ME2 ;
  RECT 190.297 0.000 190.617 0.600 ;
  LAYER ME1 ;
  RECT 190.297 0.000 190.617 0.600 ;
 END
 ANTENNAPARTIALMETALAREA                  5.273 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME3 ;
 ANTENNADIFFAREA                          1.293 LAYER ME4 ;
END DO37
PIN DI36
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 186.855 0.000 187.175 0.600 ;
  LAYER ME3 ;
  RECT 186.855 0.000 187.175 0.600 ;
  LAYER ME2 ;
  RECT 186.855 0.000 187.175 0.600 ;
  LAYER ME1 ;
  RECT 186.855 0.000 187.175 0.600 ;
 END
 ANTENNAPARTIALMETALAREA                  1.058 LAYER ME2 ;
 ANTENNAGATEAREA                          0.072 LAYER ME2 ;
 ANTENNAGATEAREA                          0.072 LAYER ME3 ;
 ANTENNAGATEAREA                          0.072 LAYER ME4 ;
 ANTENNADIFFAREA                          0.160 LAYER ME2 ;
 ANTENNADIFFAREA                          0.160 LAYER ME3 ;
 ANTENNADIFFAREA                          0.160 LAYER ME4 ;
 ANTENNAMAXAREACAR                       21.782 LAYER ME2 ;
 ANTENNAMAXAREACAR                       24.449 LAYER ME3 ;
 ANTENNAMAXAREACAR                       27.116 LAYER ME4 ;
END DI36
PIN DO36
  DIRECTION OUTPUT ;
 PORT
  LAYER ME4 ;
  RECT 186.293 0.000 186.613 0.600 ;
  LAYER ME3 ;
  RECT 186.293 0.000 186.613 0.600 ;
  LAYER ME2 ;
  RECT 186.293 0.000 186.613 0.600 ;
  LAYER ME1 ;
  RECT 186.293 0.000 186.613 0.600 ;
 END
 ANTENNAPARTIALMETALAREA                  5.273 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME3 ;
 ANTENNADIFFAREA                          1.293 LAYER ME4 ;
END DO36
PIN DI35
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 182.851 0.000 183.171 0.600 ;
  LAYER ME3 ;
  RECT 182.851 0.000 183.171 0.600 ;
  LAYER ME2 ;
  RECT 182.851 0.000 183.171 0.600 ;
  LAYER ME1 ;
  RECT 182.851 0.000 183.171 0.600 ;
 END
 ANTENNAPARTIALMETALAREA                  1.058 LAYER ME2 ;
 ANTENNAGATEAREA                          0.072 LAYER ME2 ;
 ANTENNAGATEAREA                          0.072 LAYER ME3 ;
 ANTENNAGATEAREA                          0.072 LAYER ME4 ;
 ANTENNADIFFAREA                          0.160 LAYER ME2 ;
 ANTENNADIFFAREA                          0.160 LAYER ME3 ;
 ANTENNADIFFAREA                          0.160 LAYER ME4 ;
 ANTENNAMAXAREACAR                       21.782 LAYER ME2 ;
 ANTENNAMAXAREACAR                       24.449 LAYER ME3 ;
 ANTENNAMAXAREACAR                       27.116 LAYER ME4 ;
END DI35
PIN DO35
  DIRECTION OUTPUT ;
 PORT
  LAYER ME4 ;
  RECT 182.289 0.000 182.609 0.600 ;
  LAYER ME3 ;
  RECT 182.289 0.000 182.609 0.600 ;
  LAYER ME2 ;
  RECT 182.289 0.000 182.609 0.600 ;
  LAYER ME1 ;
  RECT 182.289 0.000 182.609 0.600 ;
 END
 ANTENNAPARTIALMETALAREA                  5.273 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME3 ;
 ANTENNADIFFAREA                          1.293 LAYER ME4 ;
END DO35
PIN DI34
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 178.847 0.000 179.167 0.600 ;
  LAYER ME3 ;
  RECT 178.847 0.000 179.167 0.600 ;
  LAYER ME2 ;
  RECT 178.847 0.000 179.167 0.600 ;
  LAYER ME1 ;
  RECT 178.847 0.000 179.167 0.600 ;
 END
 ANTENNAPARTIALMETALAREA                  1.058 LAYER ME2 ;
 ANTENNAGATEAREA                          0.072 LAYER ME2 ;
 ANTENNAGATEAREA                          0.072 LAYER ME3 ;
 ANTENNAGATEAREA                          0.072 LAYER ME4 ;
 ANTENNADIFFAREA                          0.160 LAYER ME2 ;
 ANTENNADIFFAREA                          0.160 LAYER ME3 ;
 ANTENNADIFFAREA                          0.160 LAYER ME4 ;
 ANTENNAMAXAREACAR                       21.782 LAYER ME2 ;
 ANTENNAMAXAREACAR                       24.449 LAYER ME3 ;
 ANTENNAMAXAREACAR                       27.116 LAYER ME4 ;
END DI34
PIN DO34
  DIRECTION OUTPUT ;
 PORT
  LAYER ME4 ;
  RECT 178.285 0.000 178.605 0.600 ;
  LAYER ME3 ;
  RECT 178.285 0.000 178.605 0.600 ;
  LAYER ME2 ;
  RECT 178.285 0.000 178.605 0.600 ;
  LAYER ME1 ;
  RECT 178.285 0.000 178.605 0.600 ;
 END
 ANTENNAPARTIALMETALAREA                  5.273 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME3 ;
 ANTENNADIFFAREA                          1.293 LAYER ME4 ;
END DO34
PIN DI33
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 174.281 0.000 174.601 0.600 ;
  LAYER ME3 ;
  RECT 174.281 0.000 174.601 0.600 ;
  LAYER ME2 ;
  RECT 174.281 0.000 174.601 0.600 ;
  LAYER ME1 ;
  RECT 174.281 0.000 174.601 0.600 ;
 END
 ANTENNAPARTIALMETALAREA                  0.346 LAYER ME1 ;
 ANTENNAPARTIALMETALAREA                  1.466 LAYER ME2 ;
 ANTENNAPARTIALMETALAREA                  0.508 LAYER ME3 ;
 ANTENNAGATEAREA                          0.072 LAYER ME3 ;
 ANTENNAGATEAREA                          0.072 LAYER ME4 ;
 ANTENNADIFFAREA                          0.218 LAYER ME1 ;
 ANTENNADIFFAREA                          0.218 LAYER ME2 ;
 ANTENNADIFFAREA                          0.218 LAYER ME3 ;
 ANTENNADIFFAREA                          0.218 LAYER ME4 ;
 ANTENNAMAXAREACAR                       17.267 LAYER ME3 ;
 ANTENNAMAXAREACAR                       19.933 LAYER ME4 ;
END DI33
PIN DO33
  DIRECTION OUTPUT ;
 PORT
  LAYER ME4 ;
  RECT 174.843 0.000 175.163 0.600 ;
  LAYER ME3 ;
  RECT 174.843 0.000 175.163 0.600 ;
  LAYER ME2 ;
  RECT 174.843 0.000 175.163 0.600 ;
  LAYER ME1 ;
  RECT 174.843 0.000 175.163 0.600 ;
 END
 ANTENNAPARTIALMETALAREA                  5.602 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME3 ;
 ANTENNADIFFAREA                          1.293 LAYER ME4 ;
END DO33
PIN WEB3
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 172.841 0.000 173.161 0.600 ;
  LAYER ME3 ;
  RECT 172.841 0.000 173.161 0.600 ;
  LAYER ME2 ;
  RECT 172.841 0.000 173.161 0.600 ;
  LAYER ME1 ;
  RECT 172.841 0.000 173.161 0.600 ;
 END
 ANTENNAPARTIALMETALAREA                  1.036 LAYER ME2 ;
 ANTENNAGATEAREA                          0.288 LAYER ME2 ;
 ANTENNAGATEAREA                          0.288 LAYER ME3 ;
 ANTENNAGATEAREA                          0.288 LAYER ME4 ;
 ANTENNADIFFAREA                          0.206 LAYER ME2 ;
 ANTENNADIFFAREA                          0.206 LAYER ME3 ;
 ANTENNADIFFAREA                          0.206 LAYER ME4 ;
 ANTENNAMAXAREACAR                        5.844 LAYER ME2 ;
 ANTENNAMAXAREACAR                        6.511 LAYER ME3 ;
 ANTENNAMAXAREACAR                        7.178 LAYER ME4 ;
END WEB3
PIN DI32
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 170.839 0.000 171.159 0.600 ;
  LAYER ME3 ;
  RECT 170.839 0.000 171.159 0.600 ;
  LAYER ME2 ;
  RECT 170.839 0.000 171.159 0.600 ;
  LAYER ME1 ;
  RECT 170.839 0.000 171.159 0.600 ;
 END
 ANTENNAPARTIALMETALAREA                  1.058 LAYER ME2 ;
 ANTENNAGATEAREA                          0.072 LAYER ME2 ;
 ANTENNAGATEAREA                          0.072 LAYER ME3 ;
 ANTENNAGATEAREA                          0.072 LAYER ME4 ;
 ANTENNADIFFAREA                          0.160 LAYER ME2 ;
 ANTENNADIFFAREA                          0.160 LAYER ME3 ;
 ANTENNADIFFAREA                          0.160 LAYER ME4 ;
 ANTENNAMAXAREACAR                       21.782 LAYER ME2 ;
 ANTENNAMAXAREACAR                       24.449 LAYER ME3 ;
 ANTENNAMAXAREACAR                       27.116 LAYER ME4 ;
END DI32
PIN DO32
  DIRECTION OUTPUT ;
 PORT
  LAYER ME4 ;
  RECT 170.277 0.000 170.597 0.600 ;
  LAYER ME3 ;
  RECT 170.277 0.000 170.597 0.600 ;
  LAYER ME2 ;
  RECT 170.277 0.000 170.597 0.600 ;
  LAYER ME1 ;
  RECT 170.277 0.000 170.597 0.600 ;
 END
 ANTENNAPARTIALMETALAREA                  5.273 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME3 ;
 ANTENNADIFFAREA                          1.293 LAYER ME4 ;
END DO32
PIN DI31
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 166.835 0.000 167.155 0.600 ;
  LAYER ME3 ;
  RECT 166.835 0.000 167.155 0.600 ;
  LAYER ME2 ;
  RECT 166.835 0.000 167.155 0.600 ;
  LAYER ME1 ;
  RECT 166.835 0.000 167.155 0.600 ;
 END
 ANTENNAPARTIALMETALAREA                  1.058 LAYER ME2 ;
 ANTENNAGATEAREA                          0.072 LAYER ME2 ;
 ANTENNAGATEAREA                          0.072 LAYER ME3 ;
 ANTENNAGATEAREA                          0.072 LAYER ME4 ;
 ANTENNADIFFAREA                          0.160 LAYER ME2 ;
 ANTENNADIFFAREA                          0.160 LAYER ME3 ;
 ANTENNADIFFAREA                          0.160 LAYER ME4 ;
 ANTENNAMAXAREACAR                       21.782 LAYER ME2 ;
 ANTENNAMAXAREACAR                       24.449 LAYER ME3 ;
 ANTENNAMAXAREACAR                       27.116 LAYER ME4 ;
END DI31
PIN DO31
  DIRECTION OUTPUT ;
 PORT
  LAYER ME4 ;
  RECT 166.273 0.000 166.593 0.600 ;
  LAYER ME3 ;
  RECT 166.273 0.000 166.593 0.600 ;
  LAYER ME2 ;
  RECT 166.273 0.000 166.593 0.600 ;
  LAYER ME1 ;
  RECT 166.273 0.000 166.593 0.600 ;
 END
 ANTENNAPARTIALMETALAREA                  5.273 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME3 ;
 ANTENNADIFFAREA                          1.293 LAYER ME4 ;
END DO31
PIN DI30
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 162.831 0.000 163.151 0.600 ;
  LAYER ME3 ;
  RECT 162.831 0.000 163.151 0.600 ;
  LAYER ME2 ;
  RECT 162.831 0.000 163.151 0.600 ;
  LAYER ME1 ;
  RECT 162.831 0.000 163.151 0.600 ;
 END
 ANTENNAPARTIALMETALAREA                  1.058 LAYER ME2 ;
 ANTENNAGATEAREA                          0.072 LAYER ME2 ;
 ANTENNAGATEAREA                          0.072 LAYER ME3 ;
 ANTENNAGATEAREA                          0.072 LAYER ME4 ;
 ANTENNADIFFAREA                          0.160 LAYER ME2 ;
 ANTENNADIFFAREA                          0.160 LAYER ME3 ;
 ANTENNADIFFAREA                          0.160 LAYER ME4 ;
 ANTENNAMAXAREACAR                       21.782 LAYER ME2 ;
 ANTENNAMAXAREACAR                       24.449 LAYER ME3 ;
 ANTENNAMAXAREACAR                       27.116 LAYER ME4 ;
END DI30
PIN DO30
  DIRECTION OUTPUT ;
 PORT
  LAYER ME4 ;
  RECT 162.269 0.000 162.589 0.600 ;
  LAYER ME3 ;
  RECT 162.269 0.000 162.589 0.600 ;
  LAYER ME2 ;
  RECT 162.269 0.000 162.589 0.600 ;
  LAYER ME1 ;
  RECT 162.269 0.000 162.589 0.600 ;
 END
 ANTENNAPARTIALMETALAREA                  5.273 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME3 ;
 ANTENNADIFFAREA                          1.293 LAYER ME4 ;
END DO30
PIN DI29
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 158.827 0.000 159.147 0.600 ;
  LAYER ME3 ;
  RECT 158.827 0.000 159.147 0.600 ;
  LAYER ME2 ;
  RECT 158.827 0.000 159.147 0.600 ;
  LAYER ME1 ;
  RECT 158.827 0.000 159.147 0.600 ;
 END
 ANTENNAPARTIALMETALAREA                  1.058 LAYER ME2 ;
 ANTENNAGATEAREA                          0.072 LAYER ME2 ;
 ANTENNAGATEAREA                          0.072 LAYER ME3 ;
 ANTENNAGATEAREA                          0.072 LAYER ME4 ;
 ANTENNADIFFAREA                          0.160 LAYER ME2 ;
 ANTENNADIFFAREA                          0.160 LAYER ME3 ;
 ANTENNADIFFAREA                          0.160 LAYER ME4 ;
 ANTENNAMAXAREACAR                       21.782 LAYER ME2 ;
 ANTENNAMAXAREACAR                       24.449 LAYER ME3 ;
 ANTENNAMAXAREACAR                       27.116 LAYER ME4 ;
END DI29
PIN DO29
  DIRECTION OUTPUT ;
 PORT
  LAYER ME4 ;
  RECT 158.265 0.000 158.585 0.600 ;
  LAYER ME3 ;
  RECT 158.265 0.000 158.585 0.600 ;
  LAYER ME2 ;
  RECT 158.265 0.000 158.585 0.600 ;
  LAYER ME1 ;
  RECT 158.265 0.000 158.585 0.600 ;
 END
 ANTENNAPARTIALMETALAREA                  5.273 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME3 ;
 ANTENNADIFFAREA                          1.293 LAYER ME4 ;
END DO29
PIN DI28
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 154.823 0.000 155.143 0.600 ;
  LAYER ME3 ;
  RECT 154.823 0.000 155.143 0.600 ;
  LAYER ME2 ;
  RECT 154.823 0.000 155.143 0.600 ;
  LAYER ME1 ;
  RECT 154.823 0.000 155.143 0.600 ;
 END
 ANTENNAPARTIALMETALAREA                  1.058 LAYER ME2 ;
 ANTENNAGATEAREA                          0.072 LAYER ME2 ;
 ANTENNAGATEAREA                          0.072 LAYER ME3 ;
 ANTENNAGATEAREA                          0.072 LAYER ME4 ;
 ANTENNADIFFAREA                          0.160 LAYER ME2 ;
 ANTENNADIFFAREA                          0.160 LAYER ME3 ;
 ANTENNADIFFAREA                          0.160 LAYER ME4 ;
 ANTENNAMAXAREACAR                       21.782 LAYER ME2 ;
 ANTENNAMAXAREACAR                       24.449 LAYER ME3 ;
 ANTENNAMAXAREACAR                       27.116 LAYER ME4 ;
END DI28
PIN DO28
  DIRECTION OUTPUT ;
 PORT
  LAYER ME4 ;
  RECT 154.261 0.000 154.581 0.600 ;
  LAYER ME3 ;
  RECT 154.261 0.000 154.581 0.600 ;
  LAYER ME2 ;
  RECT 154.261 0.000 154.581 0.600 ;
  LAYER ME1 ;
  RECT 154.261 0.000 154.581 0.600 ;
 END
 ANTENNAPARTIALMETALAREA                  5.273 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME3 ;
 ANTENNADIFFAREA                          1.293 LAYER ME4 ;
END DO28
PIN DI27
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 150.819 0.000 151.139 0.600 ;
  LAYER ME3 ;
  RECT 150.819 0.000 151.139 0.600 ;
  LAYER ME2 ;
  RECT 150.819 0.000 151.139 0.600 ;
  LAYER ME1 ;
  RECT 150.819 0.000 151.139 0.600 ;
 END
 ANTENNAPARTIALMETALAREA                  1.058 LAYER ME2 ;
 ANTENNAGATEAREA                          0.072 LAYER ME2 ;
 ANTENNAGATEAREA                          0.072 LAYER ME3 ;
 ANTENNAGATEAREA                          0.072 LAYER ME4 ;
 ANTENNADIFFAREA                          0.160 LAYER ME2 ;
 ANTENNADIFFAREA                          0.160 LAYER ME3 ;
 ANTENNADIFFAREA                          0.160 LAYER ME4 ;
 ANTENNAMAXAREACAR                       21.782 LAYER ME2 ;
 ANTENNAMAXAREACAR                       24.449 LAYER ME3 ;
 ANTENNAMAXAREACAR                       27.116 LAYER ME4 ;
END DI27
PIN DO27
  DIRECTION OUTPUT ;
 PORT
  LAYER ME4 ;
  RECT 150.257 0.000 150.577 0.600 ;
  LAYER ME3 ;
  RECT 150.257 0.000 150.577 0.600 ;
  LAYER ME2 ;
  RECT 150.257 0.000 150.577 0.600 ;
  LAYER ME1 ;
  RECT 150.257 0.000 150.577 0.600 ;
 END
 ANTENNAPARTIALMETALAREA                  5.273 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME3 ;
 ANTENNADIFFAREA                          1.293 LAYER ME4 ;
END DO27
PIN DI26
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 146.815 0.000 147.135 0.600 ;
  LAYER ME3 ;
  RECT 146.815 0.000 147.135 0.600 ;
  LAYER ME2 ;
  RECT 146.815 0.000 147.135 0.600 ;
  LAYER ME1 ;
  RECT 146.815 0.000 147.135 0.600 ;
 END
 ANTENNAPARTIALMETALAREA                  1.058 LAYER ME2 ;
 ANTENNAGATEAREA                          0.072 LAYER ME2 ;
 ANTENNAGATEAREA                          0.072 LAYER ME3 ;
 ANTENNAGATEAREA                          0.072 LAYER ME4 ;
 ANTENNADIFFAREA                          0.160 LAYER ME2 ;
 ANTENNADIFFAREA                          0.160 LAYER ME3 ;
 ANTENNADIFFAREA                          0.160 LAYER ME4 ;
 ANTENNAMAXAREACAR                       21.782 LAYER ME2 ;
 ANTENNAMAXAREACAR                       24.449 LAYER ME3 ;
 ANTENNAMAXAREACAR                       27.116 LAYER ME4 ;
END DI26
PIN DO26
  DIRECTION OUTPUT ;
 PORT
  LAYER ME4 ;
  RECT 146.253 0.000 146.573 0.600 ;
  LAYER ME3 ;
  RECT 146.253 0.000 146.573 0.600 ;
  LAYER ME2 ;
  RECT 146.253 0.000 146.573 0.600 ;
  LAYER ME1 ;
  RECT 146.253 0.000 146.573 0.600 ;
 END
 ANTENNAPARTIALMETALAREA                  5.273 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME3 ;
 ANTENNADIFFAREA                          1.293 LAYER ME4 ;
END DO26
PIN DI25
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 142.811 0.000 143.131 0.600 ;
  LAYER ME3 ;
  RECT 142.811 0.000 143.131 0.600 ;
  LAYER ME2 ;
  RECT 142.811 0.000 143.131 0.600 ;
  LAYER ME1 ;
  RECT 142.811 0.000 143.131 0.600 ;
 END
 ANTENNAPARTIALMETALAREA                  1.058 LAYER ME2 ;
 ANTENNAGATEAREA                          0.072 LAYER ME2 ;
 ANTENNAGATEAREA                          0.072 LAYER ME3 ;
 ANTENNAGATEAREA                          0.072 LAYER ME4 ;
 ANTENNADIFFAREA                          0.160 LAYER ME2 ;
 ANTENNADIFFAREA                          0.160 LAYER ME3 ;
 ANTENNADIFFAREA                          0.160 LAYER ME4 ;
 ANTENNAMAXAREACAR                       21.782 LAYER ME2 ;
 ANTENNAMAXAREACAR                       24.449 LAYER ME3 ;
 ANTENNAMAXAREACAR                       27.116 LAYER ME4 ;
END DI25
PIN DO25
  DIRECTION OUTPUT ;
 PORT
  LAYER ME4 ;
  RECT 142.249 0.000 142.569 0.600 ;
  LAYER ME3 ;
  RECT 142.249 0.000 142.569 0.600 ;
  LAYER ME2 ;
  RECT 142.249 0.000 142.569 0.600 ;
  LAYER ME1 ;
  RECT 142.249 0.000 142.569 0.600 ;
 END
 ANTENNAPARTIALMETALAREA                  5.273 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME3 ;
 ANTENNADIFFAREA                          1.293 LAYER ME4 ;
END DO25
PIN DI24
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 138.807 0.000 139.127 0.600 ;
  LAYER ME3 ;
  RECT 138.807 0.000 139.127 0.600 ;
  LAYER ME2 ;
  RECT 138.807 0.000 139.127 0.600 ;
  LAYER ME1 ;
  RECT 138.807 0.000 139.127 0.600 ;
 END
 ANTENNAPARTIALMETALAREA                  1.058 LAYER ME2 ;
 ANTENNAGATEAREA                          0.072 LAYER ME2 ;
 ANTENNAGATEAREA                          0.072 LAYER ME3 ;
 ANTENNAGATEAREA                          0.072 LAYER ME4 ;
 ANTENNADIFFAREA                          0.160 LAYER ME2 ;
 ANTENNADIFFAREA                          0.160 LAYER ME3 ;
 ANTENNADIFFAREA                          0.160 LAYER ME4 ;
 ANTENNAMAXAREACAR                       21.782 LAYER ME2 ;
 ANTENNAMAXAREACAR                       24.449 LAYER ME3 ;
 ANTENNAMAXAREACAR                       27.116 LAYER ME4 ;
END DI24
PIN DO24
  DIRECTION OUTPUT ;
 PORT
  LAYER ME4 ;
  RECT 138.245 0.000 138.565 0.600 ;
  LAYER ME3 ;
  RECT 138.245 0.000 138.565 0.600 ;
  LAYER ME2 ;
  RECT 138.245 0.000 138.565 0.600 ;
  LAYER ME1 ;
  RECT 138.245 0.000 138.565 0.600 ;
 END
 ANTENNAPARTIALMETALAREA                  5.273 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME3 ;
 ANTENNADIFFAREA                          1.293 LAYER ME4 ;
END DO24
PIN DI23
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 134.803 0.000 135.123 0.600 ;
  LAYER ME3 ;
  RECT 134.803 0.000 135.123 0.600 ;
  LAYER ME2 ;
  RECT 134.803 0.000 135.123 0.600 ;
  LAYER ME1 ;
  RECT 134.803 0.000 135.123 0.600 ;
 END
 ANTENNAPARTIALMETALAREA                  1.058 LAYER ME2 ;
 ANTENNAGATEAREA                          0.072 LAYER ME2 ;
 ANTENNAGATEAREA                          0.072 LAYER ME3 ;
 ANTENNAGATEAREA                          0.072 LAYER ME4 ;
 ANTENNADIFFAREA                          0.160 LAYER ME2 ;
 ANTENNADIFFAREA                          0.160 LAYER ME3 ;
 ANTENNADIFFAREA                          0.160 LAYER ME4 ;
 ANTENNAMAXAREACAR                       21.782 LAYER ME2 ;
 ANTENNAMAXAREACAR                       24.449 LAYER ME3 ;
 ANTENNAMAXAREACAR                       27.116 LAYER ME4 ;
END DI23
PIN DO23
  DIRECTION OUTPUT ;
 PORT
  LAYER ME4 ;
  RECT 134.241 0.000 134.561 0.600 ;
  LAYER ME3 ;
  RECT 134.241 0.000 134.561 0.600 ;
  LAYER ME2 ;
  RECT 134.241 0.000 134.561 0.600 ;
  LAYER ME1 ;
  RECT 134.241 0.000 134.561 0.600 ;
 END
 ANTENNAPARTIALMETALAREA                  5.273 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME3 ;
 ANTENNADIFFAREA                          1.293 LAYER ME4 ;
END DO23
PIN DI22
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 130.237 0.000 130.557 0.600 ;
  LAYER ME3 ;
  RECT 130.237 0.000 130.557 0.600 ;
  LAYER ME2 ;
  RECT 130.237 0.000 130.557 0.600 ;
  LAYER ME1 ;
  RECT 130.237 0.000 130.557 0.600 ;
 END
 ANTENNAPARTIALMETALAREA                  0.346 LAYER ME1 ;
 ANTENNAPARTIALMETALAREA                  1.466 LAYER ME2 ;
 ANTENNAPARTIALMETALAREA                  0.508 LAYER ME3 ;
 ANTENNAGATEAREA                          0.072 LAYER ME3 ;
 ANTENNAGATEAREA                          0.072 LAYER ME4 ;
 ANTENNADIFFAREA                          0.218 LAYER ME1 ;
 ANTENNADIFFAREA                          0.218 LAYER ME2 ;
 ANTENNADIFFAREA                          0.218 LAYER ME3 ;
 ANTENNADIFFAREA                          0.218 LAYER ME4 ;
 ANTENNAMAXAREACAR                       17.267 LAYER ME3 ;
 ANTENNAMAXAREACAR                       19.933 LAYER ME4 ;
END DI22
PIN DO22
  DIRECTION OUTPUT ;
 PORT
  LAYER ME4 ;
  RECT 130.799 0.000 131.119 0.600 ;
  LAYER ME3 ;
  RECT 130.799 0.000 131.119 0.600 ;
  LAYER ME2 ;
  RECT 130.799 0.000 131.119 0.600 ;
  LAYER ME1 ;
  RECT 130.799 0.000 131.119 0.600 ;
 END
 ANTENNAPARTIALMETALAREA                  5.602 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME3 ;
 ANTENNADIFFAREA                          1.293 LAYER ME4 ;
END DO22
PIN WEB2
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 128.797 0.000 129.117 0.600 ;
  LAYER ME3 ;
  RECT 128.797 0.000 129.117 0.600 ;
  LAYER ME2 ;
  RECT 128.797 0.000 129.117 0.600 ;
  LAYER ME1 ;
  RECT 128.797 0.000 129.117 0.600 ;
 END
 ANTENNAPARTIALMETALAREA                  1.036 LAYER ME2 ;
 ANTENNAGATEAREA                          0.288 LAYER ME2 ;
 ANTENNAGATEAREA                          0.288 LAYER ME3 ;
 ANTENNAGATEAREA                          0.288 LAYER ME4 ;
 ANTENNADIFFAREA                          0.206 LAYER ME2 ;
 ANTENNADIFFAREA                          0.206 LAYER ME3 ;
 ANTENNADIFFAREA                          0.206 LAYER ME4 ;
 ANTENNAMAXAREACAR                        5.844 LAYER ME2 ;
 ANTENNAMAXAREACAR                        6.511 LAYER ME3 ;
 ANTENNAMAXAREACAR                        7.178 LAYER ME4 ;
END WEB2
OBS
  LAYER ME3 ;
  RECT 0.000 0.000 219.675 111.491 ;
  LAYER ME2 ;
  RECT 0.000 0.000 219.675 111.491 ;
  LAYER ME1 ;
  RECT 0.000 0.000 219.675 111.491 ;
  LAYER ME4 ;
  RECT 0.000 0.000 103.830 111.491 ;
  LAYER ME4 ;
  RECT 105.484 0.000 106.604 111.491 ;
  LAYER ME4 ;
  RECT 108.199 0.000 108.919 111.491 ;
  LAYER ME4 ;
  RECT 109.649 0.000 110.369 111.491 ;
  LAYER ME4 ;
  RECT 112.429 0.000 113.029 111.491 ;
  LAYER ME4 ;
  RECT 115.643 0.000 117.329 111.491 ;
  LAYER ME4 ;
  RECT 118.719 0.000 119.839 111.491 ;
  LAYER ME4 ;
  RECT 121.114 0.000 121.834 111.491 ;
  LAYER ME4 ;
  RECT 122.829 0.000 123.549 111.491 ;
  LAYER ME4 ;
  RECT 124.749 0.000 219.675 111.491 ;
END
END SYKB110_128X11X4CM2
END LIBRARY





