# ________________________________________________________________________________________________
# 
# 
#             Synchronous High-Density Single-Port SRAM Compiler
# 
#                 UMC 0.11um LL AE Logic Process
# 
# ________________________________________________________________________________________________
# 
#               
#         Copyright (C) 2024 Faraday Technology Corporation. All Rights Reserved.       
#                
#         This source code is an unpublished work belongs to Faraday Technology Corporation       
#         It is considered a trade secret and is not to be divulged or       
#         used by parties who have not received written authorization from       
#         Faraday Technology Corporation       
#                
#         Faraday's home page can be found at: http://www.faraday-tech.com/       
#                
# ________________________________________________________________________________________________
# 
#        IP Name            :  FSR0K_D_SH                
#        IP Version         :  1.3.0                     
#        IP Release Status  :  Active                    
#        Word               :  1024                      
#        Bit                :  16                        
#        Byte               :  8                         
#        Mux                :  1                         
#        Output Loading     :  0.01                      
#        Clock Input Slew   :  0.016                     
#        Data Input Slew    :  0.016                     
#        Ring Type          :  Ring Shape Model          
#        Ring Width         :  2                         
#        Bus Format         :  0                         
#        Memaker Path       :  /home/mem/Desktop/memlib  
#        GUI Version        :  m20230904                 
#        Date               :  2024/10/31 12:57:12       
# ________________________________________________________________________________________________
# 

VERSION 5.5 ;
NAMESCASESENSITIVE ON ;
MACRO SHKD110_1024X16X8BM1
CLASS BLOCK ;
FOREIGN SHKD110_1024X16X8BM1 0.000 0.000 ;
ORIGIN 0.000 0.000 ;
SIZE 2684.940 BY 197.930 ;
SYMMETRY x y r90 ;
SITE core ;
PIN DO127
  DIRECTION OUTPUT ;
 PORT
  LAYER ME4 ;
  RECT 2672.800 0.000 2673.600 1.000 ;
  LAYER ME3 ;
  RECT 2672.800 0.000 2673.600 1.000 ;
  LAYER ME2 ;
  RECT 2672.800 0.000 2673.600 1.000 ;
  LAYER ME1 ;
  RECT 2672.800 0.000 2673.600 1.000 ;
 END
 ANTENNAPARTIALMETALAREA                  4.176 LAYER ME2 ;
 ANTENNADIFFAREA                          5.472 LAYER ME2 ;
 ANTENNADIFFAREA                          5.472 LAYER ME3 ;
 ANTENNADIFFAREA                          5.472 LAYER ME4 ;
END DO127
PIN DI127
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 2658.400 0.000 2659.200 1.000 ;
  LAYER ME3 ;
  RECT 2658.400 0.000 2659.200 1.000 ;
  LAYER ME2 ;
  RECT 2658.400 0.000 2659.200 1.000 ;
  LAYER ME1 ;
  RECT 2658.400 0.000 2659.200 1.000 ;
 END
 ANTENNAPARTIALMETALAREA                  3.126 LAYER ME2 ;
 ANTENNAGATEAREA                          0.086 LAYER ME2 ;
 ANTENNAGATEAREA                          0.086 LAYER ME3 ;
 ANTENNAGATEAREA                          0.086 LAYER ME4 ;
 ANTENNADIFFAREA                          0.160 LAYER ME2 ;
 ANTENNADIFFAREA                          0.160 LAYER ME3 ;
 ANTENNADIFFAREA                          0.160 LAYER ME4 ;
 ANTENNAMAXAREACAR                       48.523 LAYER ME2 ;
 ANTENNAMAXAREACAR                       57.782 LAYER ME3 ;
 ANTENNAMAXAREACAR                       67.042 LAYER ME4 ;
END DI127
PIN DO126
  DIRECTION OUTPUT ;
 PORT
  LAYER ME4 ;
  RECT 2653.200 0.000 2654.000 1.000 ;
  LAYER ME3 ;
  RECT 2653.200 0.000 2654.000 1.000 ;
  LAYER ME2 ;
  RECT 2653.200 0.000 2654.000 1.000 ;
  LAYER ME1 ;
  RECT 2653.200 0.000 2654.000 1.000 ;
 END
 ANTENNAPARTIALMETALAREA                  4.152 LAYER ME2 ;
 ANTENNADIFFAREA                          5.472 LAYER ME2 ;
 ANTENNADIFFAREA                          5.472 LAYER ME3 ;
 ANTENNADIFFAREA                          5.472 LAYER ME4 ;
END DO126
PIN DI126
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 2638.400 0.000 2639.200 1.000 ;
  LAYER ME3 ;
  RECT 2638.400 0.000 2639.200 1.000 ;
  LAYER ME2 ;
  RECT 2638.400 0.000 2639.200 1.000 ;
  LAYER ME1 ;
  RECT 2638.400 0.000 2639.200 1.000 ;
 END
 ANTENNAPARTIALMETALAREA                  3.138 LAYER ME2 ;
 ANTENNAGATEAREA                          0.086 LAYER ME2 ;
 ANTENNAGATEAREA                          0.086 LAYER ME3 ;
 ANTENNAGATEAREA                          0.086 LAYER ME4 ;
 ANTENNADIFFAREA                          0.160 LAYER ME2 ;
 ANTENNADIFFAREA                          0.160 LAYER ME3 ;
 ANTENNADIFFAREA                          0.160 LAYER ME4 ;
 ANTENNAMAXAREACAR                       48.662 LAYER ME2 ;
 ANTENNAMAXAREACAR                       57.921 LAYER ME3 ;
 ANTENNAMAXAREACAR                       67.181 LAYER ME4 ;
END DI126
PIN DO125
  DIRECTION OUTPUT ;
 PORT
  LAYER ME4 ;
  RECT 2632.000 0.000 2632.800 1.000 ;
  LAYER ME3 ;
  RECT 2632.000 0.000 2632.800 1.000 ;
  LAYER ME2 ;
  RECT 2632.000 0.000 2632.800 1.000 ;
  LAYER ME1 ;
  RECT 2632.000 0.000 2632.800 1.000 ;
 END
 ANTENNAPARTIALMETALAREA                  4.152 LAYER ME2 ;
 ANTENNADIFFAREA                          5.472 LAYER ME2 ;
 ANTENNADIFFAREA                          5.472 LAYER ME3 ;
 ANTENNADIFFAREA                          5.472 LAYER ME4 ;
END DO125
PIN DI125
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 2617.600 0.000 2618.400 1.000 ;
  LAYER ME3 ;
  RECT 2617.600 0.000 2618.400 1.000 ;
  LAYER ME2 ;
  RECT 2617.600 0.000 2618.400 1.000 ;
  LAYER ME1 ;
  RECT 2617.600 0.000 2618.400 1.000 ;
 END
 ANTENNAPARTIALMETALAREA                  3.150 LAYER ME2 ;
 ANTENNAGATEAREA                          0.086 LAYER ME2 ;
 ANTENNAGATEAREA                          0.086 LAYER ME3 ;
 ANTENNAGATEAREA                          0.086 LAYER ME4 ;
 ANTENNADIFFAREA                          0.160 LAYER ME2 ;
 ANTENNADIFFAREA                          0.160 LAYER ME3 ;
 ANTENNADIFFAREA                          0.160 LAYER ME4 ;
 ANTENNAMAXAREACAR                       48.801 LAYER ME2 ;
 ANTENNAMAXAREACAR                       58.060 LAYER ME3 ;
 ANTENNAMAXAREACAR                       67.319 LAYER ME4 ;
END DI125
PIN DO124
  DIRECTION OUTPUT ;
 PORT
  LAYER ME4 ;
  RECT 2612.400 0.000 2613.200 1.000 ;
  LAYER ME3 ;
  RECT 2612.400 0.000 2613.200 1.000 ;
  LAYER ME2 ;
  RECT 2612.400 0.000 2613.200 1.000 ;
  LAYER ME1 ;
  RECT 2612.400 0.000 2613.200 1.000 ;
 END
 ANTENNAPARTIALMETALAREA                  4.176 LAYER ME2 ;
 ANTENNADIFFAREA                          5.472 LAYER ME2 ;
 ANTENNADIFFAREA                          5.472 LAYER ME3 ;
 ANTENNADIFFAREA                          5.472 LAYER ME4 ;
END DO124
PIN DI124
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 2597.600 0.000 2598.400 1.000 ;
  LAYER ME3 ;
  RECT 2597.600 0.000 2598.400 1.000 ;
  LAYER ME2 ;
  RECT 2597.600 0.000 2598.400 1.000 ;
  LAYER ME1 ;
  RECT 2597.600 0.000 2598.400 1.000 ;
 END
 ANTENNAPARTIALMETALAREA                  3.118 LAYER ME2 ;
 ANTENNAGATEAREA                          0.086 LAYER ME2 ;
 ANTENNAGATEAREA                          0.086 LAYER ME3 ;
 ANTENNAGATEAREA                          0.086 LAYER ME4 ;
 ANTENNADIFFAREA                          0.160 LAYER ME2 ;
 ANTENNADIFFAREA                          0.160 LAYER ME3 ;
 ANTENNADIFFAREA                          0.160 LAYER ME4 ;
 ANTENNAMAXAREACAR                       48.431 LAYER ME2 ;
 ANTENNAMAXAREACAR                       57.690 LAYER ME3 ;
 ANTENNAMAXAREACAR                       66.949 LAYER ME4 ;
END DI124
PIN DO123
  DIRECTION OUTPUT ;
 PORT
  LAYER ME4 ;
  RECT 2591.200 0.000 2592.000 1.000 ;
  LAYER ME3 ;
  RECT 2591.200 0.000 2592.000 1.000 ;
  LAYER ME2 ;
  RECT 2591.200 0.000 2592.000 1.000 ;
  LAYER ME1 ;
  RECT 2591.200 0.000 2592.000 1.000 ;
 END
 ANTENNAPARTIALMETALAREA                  4.152 LAYER ME2 ;
 ANTENNADIFFAREA                          5.472 LAYER ME2 ;
 ANTENNADIFFAREA                          5.472 LAYER ME3 ;
 ANTENNADIFFAREA                          5.472 LAYER ME4 ;
END DO123
PIN DI123
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 2576.400 0.000 2577.200 1.000 ;
  LAYER ME3 ;
  RECT 2576.400 0.000 2577.200 1.000 ;
  LAYER ME2 ;
  RECT 2576.400 0.000 2577.200 1.000 ;
  LAYER ME1 ;
  RECT 2576.400 0.000 2577.200 1.000 ;
 END
 ANTENNAPARTIALMETALAREA                  3.138 LAYER ME2 ;
 ANTENNAGATEAREA                          0.086 LAYER ME2 ;
 ANTENNAGATEAREA                          0.086 LAYER ME3 ;
 ANTENNAGATEAREA                          0.086 LAYER ME4 ;
 ANTENNADIFFAREA                          0.160 LAYER ME2 ;
 ANTENNADIFFAREA                          0.160 LAYER ME3 ;
 ANTENNADIFFAREA                          0.160 LAYER ME4 ;
 ANTENNAMAXAREACAR                       48.662 LAYER ME2 ;
 ANTENNAMAXAREACAR                       57.921 LAYER ME3 ;
 ANTENNAMAXAREACAR                       67.181 LAYER ME4 ;
END DI123
PIN DO122
  DIRECTION OUTPUT ;
 PORT
  LAYER ME4 ;
  RECT 2571.200 0.000 2572.000 1.000 ;
  LAYER ME3 ;
  RECT 2571.200 0.000 2572.000 1.000 ;
  LAYER ME2 ;
  RECT 2571.200 0.000 2572.000 1.000 ;
  LAYER ME1 ;
  RECT 2571.200 0.000 2572.000 1.000 ;
 END
 ANTENNAPARTIALMETALAREA                  4.160 LAYER ME2 ;
 ANTENNADIFFAREA                          5.472 LAYER ME2 ;
 ANTENNADIFFAREA                          5.472 LAYER ME3 ;
 ANTENNADIFFAREA                          5.472 LAYER ME4 ;
END DO122
PIN DI122
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 2556.800 0.000 2557.600 1.000 ;
  LAYER ME3 ;
  RECT 2556.800 0.000 2557.600 1.000 ;
  LAYER ME2 ;
  RECT 2556.800 0.000 2557.600 1.000 ;
  LAYER ME1 ;
  RECT 2556.800 0.000 2557.600 1.000 ;
 END
 ANTENNAPARTIALMETALAREA                  3.142 LAYER ME2 ;
 ANTENNAGATEAREA                          0.086 LAYER ME2 ;
 ANTENNAGATEAREA                          0.086 LAYER ME3 ;
 ANTENNAGATEAREA                          0.086 LAYER ME4 ;
 ANTENNADIFFAREA                          0.160 LAYER ME2 ;
 ANTENNADIFFAREA                          0.160 LAYER ME3 ;
 ANTENNADIFFAREA                          0.160 LAYER ME4 ;
 ANTENNAMAXAREACAR                       48.708 LAYER ME2 ;
 ANTENNAMAXAREACAR                       57.968 LAYER ME3 ;
 ANTENNAMAXAREACAR                       67.227 LAYER ME4 ;
END DI122
PIN DO121
  DIRECTION OUTPUT ;
 PORT
  LAYER ME4 ;
  RECT 2550.400 0.000 2551.200 1.000 ;
  LAYER ME3 ;
  RECT 2550.400 0.000 2551.200 1.000 ;
  LAYER ME2 ;
  RECT 2550.400 0.000 2551.200 1.000 ;
  LAYER ME1 ;
  RECT 2550.400 0.000 2551.200 1.000 ;
 END
 ANTENNAPARTIALMETALAREA                  4.176 LAYER ME2 ;
 ANTENNADIFFAREA                          5.472 LAYER ME2 ;
 ANTENNADIFFAREA                          5.472 LAYER ME3 ;
 ANTENNADIFFAREA                          5.472 LAYER ME4 ;
END DO121
PIN DI121
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 2535.600 0.000 2536.400 1.000 ;
  LAYER ME3 ;
  RECT 2535.600 0.000 2536.400 1.000 ;
  LAYER ME2 ;
  RECT 2535.600 0.000 2536.400 1.000 ;
  LAYER ME1 ;
  RECT 2535.600 0.000 2536.400 1.000 ;
 END
 ANTENNAPARTIALMETALAREA                  3.118 LAYER ME2 ;
 ANTENNAGATEAREA                          0.086 LAYER ME2 ;
 ANTENNAGATEAREA                          0.086 LAYER ME3 ;
 ANTENNAGATEAREA                          0.086 LAYER ME4 ;
 ANTENNADIFFAREA                          0.160 LAYER ME2 ;
 ANTENNADIFFAREA                          0.160 LAYER ME3 ;
 ANTENNADIFFAREA                          0.160 LAYER ME4 ;
 ANTENNAMAXAREACAR                       48.431 LAYER ME2 ;
 ANTENNAMAXAREACAR                       57.690 LAYER ME3 ;
 ANTENNAMAXAREACAR                       66.949 LAYER ME4 ;
END DI121
PIN DO120
  DIRECTION OUTPUT ;
 PORT
  LAYER ME4 ;
  RECT 2530.400 0.000 2531.200 1.000 ;
  LAYER ME3 ;
  RECT 2530.400 0.000 2531.200 1.000 ;
  LAYER ME2 ;
  RECT 2530.400 0.000 2531.200 1.000 ;
  LAYER ME1 ;
  RECT 2530.400 0.000 2531.200 1.000 ;
 END
 ANTENNAPARTIALMETALAREA                  4.144 LAYER ME2 ;
 ANTENNADIFFAREA                          5.472 LAYER ME2 ;
 ANTENNADIFFAREA                          5.472 LAYER ME3 ;
 ANTENNADIFFAREA                          5.472 LAYER ME4 ;
END DO120
PIN DI120
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 2515.600 0.000 2516.400 1.000 ;
  LAYER ME3 ;
  RECT 2515.600 0.000 2516.400 1.000 ;
  LAYER ME2 ;
  RECT 2515.600 0.000 2516.400 1.000 ;
  LAYER ME1 ;
  RECT 2515.600 0.000 2516.400 1.000 ;
 END
 ANTENNAPARTIALMETALAREA                  3.146 LAYER ME2 ;
 ANTENNAGATEAREA                          0.086 LAYER ME2 ;
 ANTENNAGATEAREA                          0.086 LAYER ME3 ;
 ANTENNAGATEAREA                          0.086 LAYER ME4 ;
 ANTENNADIFFAREA                          0.160 LAYER ME2 ;
 ANTENNADIFFAREA                          0.160 LAYER ME3 ;
 ANTENNADIFFAREA                          0.160 LAYER ME4 ;
 ANTENNAMAXAREACAR                       48.755 LAYER ME2 ;
 ANTENNAMAXAREACAR                       58.014 LAYER ME3 ;
 ANTENNAMAXAREACAR                       67.273 LAYER ME4 ;
END DI120
PIN DO119
  DIRECTION OUTPUT ;
 PORT
  LAYER ME4 ;
  RECT 2509.200 0.000 2510.000 1.000 ;
  LAYER ME3 ;
  RECT 2509.200 0.000 2510.000 1.000 ;
  LAYER ME2 ;
  RECT 2509.200 0.000 2510.000 1.000 ;
  LAYER ME1 ;
  RECT 2509.200 0.000 2510.000 1.000 ;
 END
 ANTENNAPARTIALMETALAREA                  4.160 LAYER ME2 ;
 ANTENNADIFFAREA                          5.472 LAYER ME2 ;
 ANTENNADIFFAREA                          5.472 LAYER ME3 ;
 ANTENNADIFFAREA                          5.472 LAYER ME4 ;
END DO119
PIN DI119
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 2494.800 0.000 2495.600 1.000 ;
  LAYER ME3 ;
  RECT 2494.800 0.000 2495.600 1.000 ;
  LAYER ME2 ;
  RECT 2494.800 0.000 2495.600 1.000 ;
  LAYER ME1 ;
  RECT 2494.800 0.000 2495.600 1.000 ;
 END
 ANTENNAPARTIALMETALAREA                  3.142 LAYER ME2 ;
 ANTENNAGATEAREA                          0.086 LAYER ME2 ;
 ANTENNAGATEAREA                          0.086 LAYER ME3 ;
 ANTENNAGATEAREA                          0.086 LAYER ME4 ;
 ANTENNADIFFAREA                          0.160 LAYER ME2 ;
 ANTENNADIFFAREA                          0.160 LAYER ME3 ;
 ANTENNADIFFAREA                          0.160 LAYER ME4 ;
 ANTENNAMAXAREACAR                       48.708 LAYER ME2 ;
 ANTENNAMAXAREACAR                       57.968 LAYER ME3 ;
 ANTENNAMAXAREACAR                       67.227 LAYER ME4 ;
END DI119
PIN DO118
  DIRECTION OUTPUT ;
 PORT
  LAYER ME4 ;
  RECT 2489.600 0.000 2490.400 1.000 ;
  LAYER ME3 ;
  RECT 2489.600 0.000 2490.400 1.000 ;
  LAYER ME2 ;
  RECT 2489.600 0.000 2490.400 1.000 ;
  LAYER ME1 ;
  RECT 2489.600 0.000 2490.400 1.000 ;
 END
 ANTENNAPARTIALMETALAREA                  4.168 LAYER ME2 ;
 ANTENNADIFFAREA                          5.472 LAYER ME2 ;
 ANTENNADIFFAREA                          5.472 LAYER ME3 ;
 ANTENNADIFFAREA                          5.472 LAYER ME4 ;
END DO118
PIN DI118
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 2474.800 0.000 2475.600 1.000 ;
  LAYER ME3 ;
  RECT 2474.800 0.000 2475.600 1.000 ;
  LAYER ME2 ;
  RECT 2474.800 0.000 2475.600 1.000 ;
  LAYER ME1 ;
  RECT 2474.800 0.000 2475.600 1.000 ;
 END
 ANTENNAPARTIALMETALAREA                  3.122 LAYER ME2 ;
 ANTENNAGATEAREA                          0.086 LAYER ME2 ;
 ANTENNAGATEAREA                          0.086 LAYER ME3 ;
 ANTENNAGATEAREA                          0.086 LAYER ME4 ;
 ANTENNADIFFAREA                          0.160 LAYER ME2 ;
 ANTENNADIFFAREA                          0.160 LAYER ME3 ;
 ANTENNADIFFAREA                          0.160 LAYER ME4 ;
 ANTENNAMAXAREACAR                       48.477 LAYER ME2 ;
 ANTENNAMAXAREACAR                       57.736 LAYER ME3 ;
 ANTENNAMAXAREACAR                       66.995 LAYER ME4 ;
END DI118
PIN DO117
  DIRECTION OUTPUT ;
 PORT
  LAYER ME4 ;
  RECT 2468.400 0.000 2469.200 1.000 ;
  LAYER ME3 ;
  RECT 2468.400 0.000 2469.200 1.000 ;
  LAYER ME2 ;
  RECT 2468.400 0.000 2469.200 1.000 ;
  LAYER ME1 ;
  RECT 2468.400 0.000 2469.200 1.000 ;
 END
 ANTENNAPARTIALMETALAREA                  4.144 LAYER ME2 ;
 ANTENNADIFFAREA                          5.472 LAYER ME2 ;
 ANTENNADIFFAREA                          5.472 LAYER ME3 ;
 ANTENNADIFFAREA                          5.472 LAYER ME4 ;
END DO117
PIN DI117
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 2453.600 0.000 2454.400 1.000 ;
  LAYER ME3 ;
  RECT 2453.600 0.000 2454.400 1.000 ;
  LAYER ME2 ;
  RECT 2453.600 0.000 2454.400 1.000 ;
  LAYER ME1 ;
  RECT 2453.600 0.000 2454.400 1.000 ;
 END
 ANTENNAPARTIALMETALAREA                  3.146 LAYER ME2 ;
 ANTENNAGATEAREA                          0.086 LAYER ME2 ;
 ANTENNAGATEAREA                          0.086 LAYER ME3 ;
 ANTENNAGATEAREA                          0.086 LAYER ME4 ;
 ANTENNADIFFAREA                          0.160 LAYER ME2 ;
 ANTENNADIFFAREA                          0.160 LAYER ME3 ;
 ANTENNADIFFAREA                          0.160 LAYER ME4 ;
 ANTENNAMAXAREACAR                       48.755 LAYER ME2 ;
 ANTENNAMAXAREACAR                       58.014 LAYER ME3 ;
 ANTENNAMAXAREACAR                       67.273 LAYER ME4 ;
END DI117
PIN DO116
  DIRECTION OUTPUT ;
 PORT
  LAYER ME4 ;
  RECT 2448.400 0.000 2449.200 1.000 ;
  LAYER ME3 ;
  RECT 2448.400 0.000 2449.200 1.000 ;
  LAYER ME2 ;
  RECT 2448.400 0.000 2449.200 1.000 ;
  LAYER ME1 ;
  RECT 2448.400 0.000 2449.200 1.000 ;
 END
 ANTENNAPARTIALMETALAREA                  4.168 LAYER ME2 ;
 ANTENNADIFFAREA                          5.472 LAYER ME2 ;
 ANTENNADIFFAREA                          5.472 LAYER ME3 ;
 ANTENNADIFFAREA                          5.472 LAYER ME4 ;
END DO116
PIN DI116
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 2434.000 0.000 2434.800 1.000 ;
  LAYER ME3 ;
  RECT 2434.000 0.000 2434.800 1.000 ;
  LAYER ME2 ;
  RECT 2434.000 0.000 2434.800 1.000 ;
  LAYER ME1 ;
  RECT 2434.000 0.000 2434.800 1.000 ;
 END
 ANTENNAPARTIALMETALAREA                  3.134 LAYER ME2 ;
 ANTENNAGATEAREA                          0.086 LAYER ME2 ;
 ANTENNAGATEAREA                          0.086 LAYER ME3 ;
 ANTENNAGATEAREA                          0.086 LAYER ME4 ;
 ANTENNADIFFAREA                          0.160 LAYER ME2 ;
 ANTENNADIFFAREA                          0.160 LAYER ME3 ;
 ANTENNADIFFAREA                          0.160 LAYER ME4 ;
 ANTENNAMAXAREACAR                       48.616 LAYER ME2 ;
 ANTENNAMAXAREACAR                       57.875 LAYER ME3 ;
 ANTENNAMAXAREACAR                       67.134 LAYER ME4 ;
END DI116
PIN DO115
  DIRECTION OUTPUT ;
 PORT
  LAYER ME4 ;
  RECT 2427.600 0.000 2428.400 1.000 ;
  LAYER ME3 ;
  RECT 2427.600 0.000 2428.400 1.000 ;
  LAYER ME2 ;
  RECT 2427.600 0.000 2428.400 1.000 ;
  LAYER ME1 ;
  RECT 2427.600 0.000 2428.400 1.000 ;
 END
 ANTENNAPARTIALMETALAREA                  4.168 LAYER ME2 ;
 ANTENNADIFFAREA                          5.472 LAYER ME2 ;
 ANTENNADIFFAREA                          5.472 LAYER ME3 ;
 ANTENNADIFFAREA                          5.472 LAYER ME4 ;
END DO115
PIN DI115
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 2412.800 0.000 2413.600 1.000 ;
  LAYER ME3 ;
  RECT 2412.800 0.000 2413.600 1.000 ;
  LAYER ME2 ;
  RECT 2412.800 0.000 2413.600 1.000 ;
  LAYER ME1 ;
  RECT 2412.800 0.000 2413.600 1.000 ;
 END
 ANTENNAPARTIALMETALAREA                  3.122 LAYER ME2 ;
 ANTENNAGATEAREA                          0.086 LAYER ME2 ;
 ANTENNAGATEAREA                          0.086 LAYER ME3 ;
 ANTENNAGATEAREA                          0.086 LAYER ME4 ;
 ANTENNADIFFAREA                          0.160 LAYER ME2 ;
 ANTENNADIFFAREA                          0.160 LAYER ME3 ;
 ANTENNADIFFAREA                          0.160 LAYER ME4 ;
 ANTENNAMAXAREACAR                       48.477 LAYER ME2 ;
 ANTENNAMAXAREACAR                       57.736 LAYER ME3 ;
 ANTENNAMAXAREACAR                       66.995 LAYER ME4 ;
END DI115
PIN DO114
  DIRECTION OUTPUT ;
 PORT
  LAYER ME4 ;
  RECT 2407.600 0.000 2408.400 1.000 ;
  LAYER ME3 ;
  RECT 2407.600 0.000 2408.400 1.000 ;
  LAYER ME2 ;
  RECT 2407.600 0.000 2408.400 1.000 ;
  LAYER ME1 ;
  RECT 2407.600 0.000 2408.400 1.000 ;
 END
 ANTENNAPARTIALMETALAREA                  4.144 LAYER ME2 ;
 ANTENNADIFFAREA                          5.472 LAYER ME2 ;
 ANTENNADIFFAREA                          5.472 LAYER ME3 ;
 ANTENNADIFFAREA                          5.472 LAYER ME4 ;
END DO114
PIN DI114
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 2392.800 0.000 2393.600 1.000 ;
  LAYER ME3 ;
  RECT 2392.800 0.000 2393.600 1.000 ;
  LAYER ME2 ;
  RECT 2392.800 0.000 2393.600 1.000 ;
  LAYER ME1 ;
  RECT 2392.800 0.000 2393.600 1.000 ;
 END
 ANTENNAPARTIALMETALAREA                  3.154 LAYER ME2 ;
 ANTENNAGATEAREA                          0.086 LAYER ME2 ;
 ANTENNAGATEAREA                          0.086 LAYER ME3 ;
 ANTENNAGATEAREA                          0.086 LAYER ME4 ;
 ANTENNADIFFAREA                          0.160 LAYER ME2 ;
 ANTENNADIFFAREA                          0.160 LAYER ME3 ;
 ANTENNADIFFAREA                          0.160 LAYER ME4 ;
 ANTENNAMAXAREACAR                       48.847 LAYER ME2 ;
 ANTENNAMAXAREACAR                       58.106 LAYER ME3 ;
 ANTENNAMAXAREACAR                       67.366 LAYER ME4 ;
END DI114
PIN DO113
  DIRECTION OUTPUT ;
 PORT
  LAYER ME4 ;
  RECT 2386.400 0.000 2387.200 1.000 ;
  LAYER ME3 ;
  RECT 2386.400 0.000 2387.200 1.000 ;
  LAYER ME2 ;
  RECT 2386.400 0.000 2387.200 1.000 ;
  LAYER ME1 ;
  RECT 2386.400 0.000 2387.200 1.000 ;
 END
 ANTENNAPARTIALMETALAREA                  4.168 LAYER ME2 ;
 ANTENNADIFFAREA                          5.472 LAYER ME2 ;
 ANTENNADIFFAREA                          5.472 LAYER ME3 ;
 ANTENNADIFFAREA                          5.472 LAYER ME4 ;
END DO113
PIN DI113
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 2372.000 0.000 2372.800 1.000 ;
  LAYER ME3 ;
  RECT 2372.000 0.000 2372.800 1.000 ;
  LAYER ME2 ;
  RECT 2372.000 0.000 2372.800 1.000 ;
  LAYER ME1 ;
  RECT 2372.000 0.000 2372.800 1.000 ;
 END
 ANTENNAPARTIALMETALAREA                  3.134 LAYER ME2 ;
 ANTENNAGATEAREA                          0.086 LAYER ME2 ;
 ANTENNAGATEAREA                          0.086 LAYER ME3 ;
 ANTENNAGATEAREA                          0.086 LAYER ME4 ;
 ANTENNADIFFAREA                          0.160 LAYER ME2 ;
 ANTENNADIFFAREA                          0.160 LAYER ME3 ;
 ANTENNADIFFAREA                          0.160 LAYER ME4 ;
 ANTENNAMAXAREACAR                       48.616 LAYER ME2 ;
 ANTENNAMAXAREACAR                       57.875 LAYER ME3 ;
 ANTENNAMAXAREACAR                       67.134 LAYER ME4 ;
END DI113
PIN DO112
  DIRECTION OUTPUT ;
 PORT
  LAYER ME4 ;
  RECT 2366.800 0.000 2367.600 1.000 ;
  LAYER ME3 ;
  RECT 2366.800 0.000 2367.600 1.000 ;
  LAYER ME2 ;
  RECT 2366.800 0.000 2367.600 1.000 ;
  LAYER ME1 ;
  RECT 2366.800 0.000 2367.600 1.000 ;
 END
 ANTENNAPARTIALMETALAREA                  4.160 LAYER ME2 ;
 ANTENNADIFFAREA                          5.472 LAYER ME2 ;
 ANTENNADIFFAREA                          5.472 LAYER ME3 ;
 ANTENNADIFFAREA                          5.472 LAYER ME4 ;
END DO112
PIN WEB7
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 2353.600 0.000 2354.400 1.000 ;
  LAYER ME3 ;
  RECT 2353.600 0.000 2354.400 1.000 ;
  LAYER ME2 ;
  RECT 2353.600 0.000 2354.400 1.000 ;
  LAYER ME1 ;
  RECT 2353.600 0.000 2354.400 1.000 ;
 END
 ANTENNAPARTIALMETALAREA                  2.868 LAYER ME2 ;
 ANTENNAGATEAREA                          0.072 LAYER ME2 ;
 ANTENNAGATEAREA                          0.072 LAYER ME3 ;
 ANTENNAGATEAREA                          0.072 LAYER ME4 ;
 ANTENNADIFFAREA                          0.160 LAYER ME2 ;
 ANTENNADIFFAREA                          0.160 LAYER ME3 ;
 ANTENNADIFFAREA                          0.160 LAYER ME4 ;
 ANTENNAMAXAREACAR                       54.844 LAYER ME2 ;
 ANTENNAMAXAREACAR                       65.956 LAYER ME3 ;
 ANTENNAMAXAREACAR                       77.067 LAYER ME4 ;
END WEB7
PIN DI112
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 2352.000 0.000 2352.800 1.000 ;
  LAYER ME3 ;
  RECT 2352.000 0.000 2352.800 1.000 ;
  LAYER ME2 ;
  RECT 2352.000 0.000 2352.800 1.000 ;
  LAYER ME1 ;
  RECT 2352.000 0.000 2352.800 1.000 ;
 END
 ANTENNAPARTIALMETALAREA                  3.130 LAYER ME2 ;
 ANTENNAGATEAREA                          0.086 LAYER ME2 ;
 ANTENNAGATEAREA                          0.086 LAYER ME3 ;
 ANTENNAGATEAREA                          0.086 LAYER ME4 ;
 ANTENNADIFFAREA                          0.160 LAYER ME2 ;
 ANTENNADIFFAREA                          0.160 LAYER ME3 ;
 ANTENNADIFFAREA                          0.160 LAYER ME4 ;
 ANTENNAMAXAREACAR                       48.569 LAYER ME2 ;
 ANTENNAMAXAREACAR                       57.829 LAYER ME3 ;
 ANTENNAMAXAREACAR                       67.088 LAYER ME4 ;
END DI112
PIN DO111
  DIRECTION OUTPUT ;
 PORT
  LAYER ME4 ;
  RECT 2345.600 0.000 2346.400 1.000 ;
  LAYER ME3 ;
  RECT 2345.600 0.000 2346.400 1.000 ;
  LAYER ME2 ;
  RECT 2345.600 0.000 2346.400 1.000 ;
  LAYER ME1 ;
  RECT 2345.600 0.000 2346.400 1.000 ;
 END
 ANTENNAPARTIALMETALAREA                  4.144 LAYER ME2 ;
 ANTENNADIFFAREA                          5.472 LAYER ME2 ;
 ANTENNADIFFAREA                          5.472 LAYER ME3 ;
 ANTENNADIFFAREA                          5.472 LAYER ME4 ;
END DO111
PIN DI111
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 2330.800 0.000 2331.600 1.000 ;
  LAYER ME3 ;
  RECT 2330.800 0.000 2331.600 1.000 ;
  LAYER ME2 ;
  RECT 2330.800 0.000 2331.600 1.000 ;
  LAYER ME1 ;
  RECT 2330.800 0.000 2331.600 1.000 ;
 END
 ANTENNAPARTIALMETALAREA                  3.154 LAYER ME2 ;
 ANTENNAGATEAREA                          0.086 LAYER ME2 ;
 ANTENNAGATEAREA                          0.086 LAYER ME3 ;
 ANTENNAGATEAREA                          0.086 LAYER ME4 ;
 ANTENNADIFFAREA                          0.160 LAYER ME2 ;
 ANTENNADIFFAREA                          0.160 LAYER ME3 ;
 ANTENNADIFFAREA                          0.160 LAYER ME4 ;
 ANTENNAMAXAREACAR                       48.847 LAYER ME2 ;
 ANTENNAMAXAREACAR                       58.106 LAYER ME3 ;
 ANTENNAMAXAREACAR                       67.366 LAYER ME4 ;
END DI111
PIN DO110
  DIRECTION OUTPUT ;
 PORT
  LAYER ME4 ;
  RECT 2325.600 0.000 2326.400 1.000 ;
  LAYER ME3 ;
  RECT 2325.600 0.000 2326.400 1.000 ;
  LAYER ME2 ;
  RECT 2325.600 0.000 2326.400 1.000 ;
  LAYER ME1 ;
  RECT 2325.600 0.000 2326.400 1.000 ;
 END
 ANTENNAPARTIALMETALAREA                  4.176 LAYER ME2 ;
 ANTENNADIFFAREA                          5.472 LAYER ME2 ;
 ANTENNADIFFAREA                          5.472 LAYER ME3 ;
 ANTENNADIFFAREA                          5.472 LAYER ME4 ;
END DO110
PIN DI110
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 2311.200 0.000 2312.000 1.000 ;
  LAYER ME3 ;
  RECT 2311.200 0.000 2312.000 1.000 ;
  LAYER ME2 ;
  RECT 2311.200 0.000 2312.000 1.000 ;
  LAYER ME1 ;
  RECT 2311.200 0.000 2312.000 1.000 ;
 END
 ANTENNAPARTIALMETALAREA                  3.126 LAYER ME2 ;
 ANTENNAGATEAREA                          0.086 LAYER ME2 ;
 ANTENNAGATEAREA                          0.086 LAYER ME3 ;
 ANTENNAGATEAREA                          0.086 LAYER ME4 ;
 ANTENNADIFFAREA                          0.160 LAYER ME2 ;
 ANTENNADIFFAREA                          0.160 LAYER ME3 ;
 ANTENNADIFFAREA                          0.160 LAYER ME4 ;
 ANTENNAMAXAREACAR                       48.523 LAYER ME2 ;
 ANTENNAMAXAREACAR                       57.782 LAYER ME3 ;
 ANTENNAMAXAREACAR                       67.042 LAYER ME4 ;
END DI110
PIN DO109
  DIRECTION OUTPUT ;
 PORT
  LAYER ME4 ;
  RECT 2304.800 0.000 2305.600 1.000 ;
  LAYER ME3 ;
  RECT 2304.800 0.000 2305.600 1.000 ;
  LAYER ME2 ;
  RECT 2304.800 0.000 2305.600 1.000 ;
  LAYER ME1 ;
  RECT 2304.800 0.000 2305.600 1.000 ;
 END
 ANTENNAPARTIALMETALAREA                  4.160 LAYER ME2 ;
 ANTENNADIFFAREA                          5.472 LAYER ME2 ;
 ANTENNADIFFAREA                          5.472 LAYER ME3 ;
 ANTENNADIFFAREA                          5.472 LAYER ME4 ;
END DO109
PIN DI109
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 2290.000 0.000 2290.800 1.000 ;
  LAYER ME3 ;
  RECT 2290.000 0.000 2290.800 1.000 ;
  LAYER ME2 ;
  RECT 2290.000 0.000 2290.800 1.000 ;
  LAYER ME1 ;
  RECT 2290.000 0.000 2290.800 1.000 ;
 END
 ANTENNAPARTIALMETALAREA                  3.130 LAYER ME2 ;
 ANTENNAGATEAREA                          0.086 LAYER ME2 ;
 ANTENNAGATEAREA                          0.086 LAYER ME3 ;
 ANTENNAGATEAREA                          0.086 LAYER ME4 ;
 ANTENNADIFFAREA                          0.160 LAYER ME2 ;
 ANTENNADIFFAREA                          0.160 LAYER ME3 ;
 ANTENNADIFFAREA                          0.160 LAYER ME4 ;
 ANTENNAMAXAREACAR                       48.569 LAYER ME2 ;
 ANTENNAMAXAREACAR                       57.829 LAYER ME3 ;
 ANTENNAMAXAREACAR                       67.088 LAYER ME4 ;
END DI109
PIN DO108
  DIRECTION OUTPUT ;
 PORT
  LAYER ME4 ;
  RECT 2284.800 0.000 2285.600 1.000 ;
  LAYER ME3 ;
  RECT 2284.800 0.000 2285.600 1.000 ;
  LAYER ME2 ;
  RECT 2284.800 0.000 2285.600 1.000 ;
  LAYER ME1 ;
  RECT 2284.800 0.000 2285.600 1.000 ;
 END
 ANTENNAPARTIALMETALAREA                  4.152 LAYER ME2 ;
 ANTENNADIFFAREA                          5.472 LAYER ME2 ;
 ANTENNADIFFAREA                          5.472 LAYER ME3 ;
 ANTENNADIFFAREA                          5.472 LAYER ME4 ;
END DO108
PIN DI108
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 2270.400 0.000 2271.200 1.000 ;
  LAYER ME3 ;
  RECT 2270.400 0.000 2271.200 1.000 ;
  LAYER ME2 ;
  RECT 2270.400 0.000 2271.200 1.000 ;
  LAYER ME1 ;
  RECT 2270.400 0.000 2271.200 1.000 ;
 END
 ANTENNAPARTIALMETALAREA                  3.150 LAYER ME2 ;
 ANTENNAGATEAREA                          0.086 LAYER ME2 ;
 ANTENNAGATEAREA                          0.086 LAYER ME3 ;
 ANTENNAGATEAREA                          0.086 LAYER ME4 ;
 ANTENNADIFFAREA                          0.160 LAYER ME2 ;
 ANTENNADIFFAREA                          0.160 LAYER ME3 ;
 ANTENNADIFFAREA                          0.160 LAYER ME4 ;
 ANTENNAMAXAREACAR                       48.801 LAYER ME2 ;
 ANTENNAMAXAREACAR                       58.060 LAYER ME3 ;
 ANTENNAMAXAREACAR                       67.319 LAYER ME4 ;
END DI108
PIN DO107
  DIRECTION OUTPUT ;
 PORT
  LAYER ME4 ;
  RECT 2263.600 0.000 2264.400 1.000 ;
  LAYER ME3 ;
  RECT 2263.600 0.000 2264.400 1.000 ;
  LAYER ME2 ;
  RECT 2263.600 0.000 2264.400 1.000 ;
  LAYER ME1 ;
  RECT 2263.600 0.000 2264.400 1.000 ;
 END
 ANTENNAPARTIALMETALAREA                  4.176 LAYER ME2 ;
 ANTENNADIFFAREA                          5.472 LAYER ME2 ;
 ANTENNADIFFAREA                          5.472 LAYER ME3 ;
 ANTENNADIFFAREA                          5.472 LAYER ME4 ;
END DO107
PIN DI107
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 2249.200 0.000 2250.000 1.000 ;
  LAYER ME3 ;
  RECT 2249.200 0.000 2250.000 1.000 ;
  LAYER ME2 ;
  RECT 2249.200 0.000 2250.000 1.000 ;
  LAYER ME1 ;
  RECT 2249.200 0.000 2250.000 1.000 ;
 END
 ANTENNAPARTIALMETALAREA                  3.126 LAYER ME2 ;
 ANTENNAGATEAREA                          0.086 LAYER ME2 ;
 ANTENNAGATEAREA                          0.086 LAYER ME3 ;
 ANTENNAGATEAREA                          0.086 LAYER ME4 ;
 ANTENNADIFFAREA                          0.160 LAYER ME2 ;
 ANTENNADIFFAREA                          0.160 LAYER ME3 ;
 ANTENNADIFFAREA                          0.160 LAYER ME4 ;
 ANTENNAMAXAREACAR                       48.523 LAYER ME2 ;
 ANTENNAMAXAREACAR                       57.782 LAYER ME3 ;
 ANTENNAMAXAREACAR                       67.042 LAYER ME4 ;
END DI107
PIN DO106
  DIRECTION OUTPUT ;
 PORT
  LAYER ME4 ;
  RECT 2244.000 0.000 2244.800 1.000 ;
  LAYER ME3 ;
  RECT 2244.000 0.000 2244.800 1.000 ;
  LAYER ME2 ;
  RECT 2244.000 0.000 2244.800 1.000 ;
  LAYER ME1 ;
  RECT 2244.000 0.000 2244.800 1.000 ;
 END
 ANTENNAPARTIALMETALAREA                  4.152 LAYER ME2 ;
 ANTENNADIFFAREA                          5.472 LAYER ME2 ;
 ANTENNADIFFAREA                          5.472 LAYER ME3 ;
 ANTENNADIFFAREA                          5.472 LAYER ME4 ;
END DO106
PIN DI106
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 2229.200 0.000 2230.000 1.000 ;
  LAYER ME3 ;
  RECT 2229.200 0.000 2230.000 1.000 ;
  LAYER ME2 ;
  RECT 2229.200 0.000 2230.000 1.000 ;
  LAYER ME1 ;
  RECT 2229.200 0.000 2230.000 1.000 ;
 END
 ANTENNAPARTIALMETALAREA                  3.138 LAYER ME2 ;
 ANTENNAGATEAREA                          0.086 LAYER ME2 ;
 ANTENNAGATEAREA                          0.086 LAYER ME3 ;
 ANTENNAGATEAREA                          0.086 LAYER ME4 ;
 ANTENNADIFFAREA                          0.160 LAYER ME2 ;
 ANTENNADIFFAREA                          0.160 LAYER ME3 ;
 ANTENNADIFFAREA                          0.160 LAYER ME4 ;
 ANTENNAMAXAREACAR                       48.662 LAYER ME2 ;
 ANTENNAMAXAREACAR                       57.921 LAYER ME3 ;
 ANTENNAMAXAREACAR                       67.181 LAYER ME4 ;
END DI106
PIN DO105
  DIRECTION OUTPUT ;
 PORT
  LAYER ME4 ;
  RECT 2222.800 0.000 2223.600 1.000 ;
  LAYER ME3 ;
  RECT 2222.800 0.000 2223.600 1.000 ;
  LAYER ME2 ;
  RECT 2222.800 0.000 2223.600 1.000 ;
  LAYER ME1 ;
  RECT 2222.800 0.000 2223.600 1.000 ;
 END
 ANTENNAPARTIALMETALAREA                  4.152 LAYER ME2 ;
 ANTENNADIFFAREA                          5.472 LAYER ME2 ;
 ANTENNADIFFAREA                          5.472 LAYER ME3 ;
 ANTENNADIFFAREA                          5.472 LAYER ME4 ;
END DO105
PIN DI105
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 2208.400 0.000 2209.200 1.000 ;
  LAYER ME3 ;
  RECT 2208.400 0.000 2209.200 1.000 ;
  LAYER ME2 ;
  RECT 2208.400 0.000 2209.200 1.000 ;
  LAYER ME1 ;
  RECT 2208.400 0.000 2209.200 1.000 ;
 END
 ANTENNAPARTIALMETALAREA                  3.150 LAYER ME2 ;
 ANTENNAGATEAREA                          0.086 LAYER ME2 ;
 ANTENNAGATEAREA                          0.086 LAYER ME3 ;
 ANTENNAGATEAREA                          0.086 LAYER ME4 ;
 ANTENNADIFFAREA                          0.160 LAYER ME2 ;
 ANTENNADIFFAREA                          0.160 LAYER ME3 ;
 ANTENNADIFFAREA                          0.160 LAYER ME4 ;
 ANTENNAMAXAREACAR                       48.801 LAYER ME2 ;
 ANTENNAMAXAREACAR                       58.060 LAYER ME3 ;
 ANTENNAMAXAREACAR                       67.319 LAYER ME4 ;
END DI105
PIN DO104
  DIRECTION OUTPUT ;
 PORT
  LAYER ME4 ;
  RECT 2203.200 0.000 2204.000 1.000 ;
  LAYER ME3 ;
  RECT 2203.200 0.000 2204.000 1.000 ;
  LAYER ME2 ;
  RECT 2203.200 0.000 2204.000 1.000 ;
  LAYER ME1 ;
  RECT 2203.200 0.000 2204.000 1.000 ;
 END
 ANTENNAPARTIALMETALAREA                  4.176 LAYER ME2 ;
 ANTENNADIFFAREA                          5.472 LAYER ME2 ;
 ANTENNADIFFAREA                          5.472 LAYER ME3 ;
 ANTENNADIFFAREA                          5.472 LAYER ME4 ;
END DO104
PIN DI104
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 2188.400 0.000 2189.200 1.000 ;
  LAYER ME3 ;
  RECT 2188.400 0.000 2189.200 1.000 ;
  LAYER ME2 ;
  RECT 2188.400 0.000 2189.200 1.000 ;
  LAYER ME1 ;
  RECT 2188.400 0.000 2189.200 1.000 ;
 END
 ANTENNAPARTIALMETALAREA                  3.118 LAYER ME2 ;
 ANTENNAGATEAREA                          0.086 LAYER ME2 ;
 ANTENNAGATEAREA                          0.086 LAYER ME3 ;
 ANTENNAGATEAREA                          0.086 LAYER ME4 ;
 ANTENNADIFFAREA                          0.160 LAYER ME2 ;
 ANTENNADIFFAREA                          0.160 LAYER ME3 ;
 ANTENNADIFFAREA                          0.160 LAYER ME4 ;
 ANTENNAMAXAREACAR                       48.431 LAYER ME2 ;
 ANTENNAMAXAREACAR                       57.690 LAYER ME3 ;
 ANTENNAMAXAREACAR                       66.949 LAYER ME4 ;
END DI104
PIN DO103
  DIRECTION OUTPUT ;
 PORT
  LAYER ME4 ;
  RECT 2182.000 0.000 2182.800 1.000 ;
  LAYER ME3 ;
  RECT 2182.000 0.000 2182.800 1.000 ;
  LAYER ME2 ;
  RECT 2182.000 0.000 2182.800 1.000 ;
  LAYER ME1 ;
  RECT 2182.000 0.000 2182.800 1.000 ;
 END
 ANTENNAPARTIALMETALAREA                  4.152 LAYER ME2 ;
 ANTENNADIFFAREA                          5.472 LAYER ME2 ;
 ANTENNADIFFAREA                          5.472 LAYER ME3 ;
 ANTENNADIFFAREA                          5.472 LAYER ME4 ;
END DO103
PIN DI103
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 2167.200 0.000 2168.000 1.000 ;
  LAYER ME3 ;
  RECT 2167.200 0.000 2168.000 1.000 ;
  LAYER ME2 ;
  RECT 2167.200 0.000 2168.000 1.000 ;
  LAYER ME1 ;
  RECT 2167.200 0.000 2168.000 1.000 ;
 END
 ANTENNAPARTIALMETALAREA                  3.138 LAYER ME2 ;
 ANTENNAGATEAREA                          0.086 LAYER ME2 ;
 ANTENNAGATEAREA                          0.086 LAYER ME3 ;
 ANTENNAGATEAREA                          0.086 LAYER ME4 ;
 ANTENNADIFFAREA                          0.160 LAYER ME2 ;
 ANTENNADIFFAREA                          0.160 LAYER ME3 ;
 ANTENNADIFFAREA                          0.160 LAYER ME4 ;
 ANTENNAMAXAREACAR                       48.662 LAYER ME2 ;
 ANTENNAMAXAREACAR                       57.921 LAYER ME3 ;
 ANTENNAMAXAREACAR                       67.181 LAYER ME4 ;
END DI103
PIN DO102
  DIRECTION OUTPUT ;
 PORT
  LAYER ME4 ;
  RECT 2162.000 0.000 2162.800 1.000 ;
  LAYER ME3 ;
  RECT 2162.000 0.000 2162.800 1.000 ;
  LAYER ME2 ;
  RECT 2162.000 0.000 2162.800 1.000 ;
  LAYER ME1 ;
  RECT 2162.000 0.000 2162.800 1.000 ;
 END
 ANTENNAPARTIALMETALAREA                  4.160 LAYER ME2 ;
 ANTENNADIFFAREA                          5.472 LAYER ME2 ;
 ANTENNADIFFAREA                          5.472 LAYER ME3 ;
 ANTENNADIFFAREA                          5.472 LAYER ME4 ;
END DO102
PIN DI102
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 2147.600 0.000 2148.400 1.000 ;
  LAYER ME3 ;
  RECT 2147.600 0.000 2148.400 1.000 ;
  LAYER ME2 ;
  RECT 2147.600 0.000 2148.400 1.000 ;
  LAYER ME1 ;
  RECT 2147.600 0.000 2148.400 1.000 ;
 END
 ANTENNAPARTIALMETALAREA                  3.142 LAYER ME2 ;
 ANTENNAGATEAREA                          0.086 LAYER ME2 ;
 ANTENNAGATEAREA                          0.086 LAYER ME3 ;
 ANTENNAGATEAREA                          0.086 LAYER ME4 ;
 ANTENNADIFFAREA                          0.160 LAYER ME2 ;
 ANTENNADIFFAREA                          0.160 LAYER ME3 ;
 ANTENNADIFFAREA                          0.160 LAYER ME4 ;
 ANTENNAMAXAREACAR                       48.708 LAYER ME2 ;
 ANTENNAMAXAREACAR                       57.968 LAYER ME3 ;
 ANTENNAMAXAREACAR                       67.227 LAYER ME4 ;
END DI102
PIN DO101
  DIRECTION OUTPUT ;
 PORT
  LAYER ME4 ;
  RECT 2141.200 0.000 2142.000 1.000 ;
  LAYER ME3 ;
  RECT 2141.200 0.000 2142.000 1.000 ;
  LAYER ME2 ;
  RECT 2141.200 0.000 2142.000 1.000 ;
  LAYER ME1 ;
  RECT 2141.200 0.000 2142.000 1.000 ;
 END
 ANTENNAPARTIALMETALAREA                  4.176 LAYER ME2 ;
 ANTENNADIFFAREA                          5.472 LAYER ME2 ;
 ANTENNADIFFAREA                          5.472 LAYER ME3 ;
 ANTENNADIFFAREA                          5.472 LAYER ME4 ;
END DO101
PIN DI101
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 2126.400 0.000 2127.200 1.000 ;
  LAYER ME3 ;
  RECT 2126.400 0.000 2127.200 1.000 ;
  LAYER ME2 ;
  RECT 2126.400 0.000 2127.200 1.000 ;
  LAYER ME1 ;
  RECT 2126.400 0.000 2127.200 1.000 ;
 END
 ANTENNAPARTIALMETALAREA                  3.118 LAYER ME2 ;
 ANTENNAGATEAREA                          0.086 LAYER ME2 ;
 ANTENNAGATEAREA                          0.086 LAYER ME3 ;
 ANTENNAGATEAREA                          0.086 LAYER ME4 ;
 ANTENNADIFFAREA                          0.160 LAYER ME2 ;
 ANTENNADIFFAREA                          0.160 LAYER ME3 ;
 ANTENNADIFFAREA                          0.160 LAYER ME4 ;
 ANTENNAMAXAREACAR                       48.431 LAYER ME2 ;
 ANTENNAMAXAREACAR                       57.690 LAYER ME3 ;
 ANTENNAMAXAREACAR                       66.949 LAYER ME4 ;
END DI101
PIN DO100
  DIRECTION OUTPUT ;
 PORT
  LAYER ME4 ;
  RECT 2121.200 0.000 2122.000 1.000 ;
  LAYER ME3 ;
  RECT 2121.200 0.000 2122.000 1.000 ;
  LAYER ME2 ;
  RECT 2121.200 0.000 2122.000 1.000 ;
  LAYER ME1 ;
  RECT 2121.200 0.000 2122.000 1.000 ;
 END
 ANTENNAPARTIALMETALAREA                  4.144 LAYER ME2 ;
 ANTENNADIFFAREA                          5.472 LAYER ME2 ;
 ANTENNADIFFAREA                          5.472 LAYER ME3 ;
 ANTENNADIFFAREA                          5.472 LAYER ME4 ;
END DO100
PIN DI100
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 2106.400 0.000 2107.200 1.000 ;
  LAYER ME3 ;
  RECT 2106.400 0.000 2107.200 1.000 ;
  LAYER ME2 ;
  RECT 2106.400 0.000 2107.200 1.000 ;
  LAYER ME1 ;
  RECT 2106.400 0.000 2107.200 1.000 ;
 END
 ANTENNAPARTIALMETALAREA                  3.146 LAYER ME2 ;
 ANTENNAGATEAREA                          0.086 LAYER ME2 ;
 ANTENNAGATEAREA                          0.086 LAYER ME3 ;
 ANTENNAGATEAREA                          0.086 LAYER ME4 ;
 ANTENNADIFFAREA                          0.160 LAYER ME2 ;
 ANTENNADIFFAREA                          0.160 LAYER ME3 ;
 ANTENNADIFFAREA                          0.160 LAYER ME4 ;
 ANTENNAMAXAREACAR                       48.755 LAYER ME2 ;
 ANTENNAMAXAREACAR                       58.014 LAYER ME3 ;
 ANTENNAMAXAREACAR                       67.273 LAYER ME4 ;
END DI100
PIN DO99
  DIRECTION OUTPUT ;
 PORT
  LAYER ME4 ;
  RECT 2100.000 0.000 2100.800 1.000 ;
  LAYER ME3 ;
  RECT 2100.000 0.000 2100.800 1.000 ;
  LAYER ME2 ;
  RECT 2100.000 0.000 2100.800 1.000 ;
  LAYER ME1 ;
  RECT 2100.000 0.000 2100.800 1.000 ;
 END
 ANTENNAPARTIALMETALAREA                  4.160 LAYER ME2 ;
 ANTENNADIFFAREA                          5.472 LAYER ME2 ;
 ANTENNADIFFAREA                          5.472 LAYER ME3 ;
 ANTENNADIFFAREA                          5.472 LAYER ME4 ;
END DO99
PIN DI99
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 2085.600 0.000 2086.400 1.000 ;
  LAYER ME3 ;
  RECT 2085.600 0.000 2086.400 1.000 ;
  LAYER ME2 ;
  RECT 2085.600 0.000 2086.400 1.000 ;
  LAYER ME1 ;
  RECT 2085.600 0.000 2086.400 1.000 ;
 END
 ANTENNAPARTIALMETALAREA                  3.142 LAYER ME2 ;
 ANTENNAGATEAREA                          0.086 LAYER ME2 ;
 ANTENNAGATEAREA                          0.086 LAYER ME3 ;
 ANTENNAGATEAREA                          0.086 LAYER ME4 ;
 ANTENNADIFFAREA                          0.160 LAYER ME2 ;
 ANTENNADIFFAREA                          0.160 LAYER ME3 ;
 ANTENNADIFFAREA                          0.160 LAYER ME4 ;
 ANTENNAMAXAREACAR                       48.708 LAYER ME2 ;
 ANTENNAMAXAREACAR                       57.968 LAYER ME3 ;
 ANTENNAMAXAREACAR                       67.227 LAYER ME4 ;
END DI99
PIN DO98
  DIRECTION OUTPUT ;
 PORT
  LAYER ME4 ;
  RECT 2080.400 0.000 2081.200 1.000 ;
  LAYER ME3 ;
  RECT 2080.400 0.000 2081.200 1.000 ;
  LAYER ME2 ;
  RECT 2080.400 0.000 2081.200 1.000 ;
  LAYER ME1 ;
  RECT 2080.400 0.000 2081.200 1.000 ;
 END
 ANTENNAPARTIALMETALAREA                  4.168 LAYER ME2 ;
 ANTENNADIFFAREA                          5.472 LAYER ME2 ;
 ANTENNADIFFAREA                          5.472 LAYER ME3 ;
 ANTENNADIFFAREA                          5.472 LAYER ME4 ;
END DO98
PIN DI98
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 2065.600 0.000 2066.400 1.000 ;
  LAYER ME3 ;
  RECT 2065.600 0.000 2066.400 1.000 ;
  LAYER ME2 ;
  RECT 2065.600 0.000 2066.400 1.000 ;
  LAYER ME1 ;
  RECT 2065.600 0.000 2066.400 1.000 ;
 END
 ANTENNAPARTIALMETALAREA                  3.122 LAYER ME2 ;
 ANTENNAGATEAREA                          0.086 LAYER ME2 ;
 ANTENNAGATEAREA                          0.086 LAYER ME3 ;
 ANTENNAGATEAREA                          0.086 LAYER ME4 ;
 ANTENNADIFFAREA                          0.160 LAYER ME2 ;
 ANTENNADIFFAREA                          0.160 LAYER ME3 ;
 ANTENNADIFFAREA                          0.160 LAYER ME4 ;
 ANTENNAMAXAREACAR                       48.477 LAYER ME2 ;
 ANTENNAMAXAREACAR                       57.736 LAYER ME3 ;
 ANTENNAMAXAREACAR                       66.995 LAYER ME4 ;
END DI98
PIN DO97
  DIRECTION OUTPUT ;
 PORT
  LAYER ME4 ;
  RECT 2059.200 0.000 2060.000 1.000 ;
  LAYER ME3 ;
  RECT 2059.200 0.000 2060.000 1.000 ;
  LAYER ME2 ;
  RECT 2059.200 0.000 2060.000 1.000 ;
  LAYER ME1 ;
  RECT 2059.200 0.000 2060.000 1.000 ;
 END
 ANTENNAPARTIALMETALAREA                  4.144 LAYER ME2 ;
 ANTENNADIFFAREA                          5.472 LAYER ME2 ;
 ANTENNADIFFAREA                          5.472 LAYER ME3 ;
 ANTENNADIFFAREA                          5.472 LAYER ME4 ;
END DO97
PIN DI97
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 2044.400 0.000 2045.200 1.000 ;
  LAYER ME3 ;
  RECT 2044.400 0.000 2045.200 1.000 ;
  LAYER ME2 ;
  RECT 2044.400 0.000 2045.200 1.000 ;
  LAYER ME1 ;
  RECT 2044.400 0.000 2045.200 1.000 ;
 END
 ANTENNAPARTIALMETALAREA                  3.146 LAYER ME2 ;
 ANTENNAGATEAREA                          0.086 LAYER ME2 ;
 ANTENNAGATEAREA                          0.086 LAYER ME3 ;
 ANTENNAGATEAREA                          0.086 LAYER ME4 ;
 ANTENNADIFFAREA                          0.160 LAYER ME2 ;
 ANTENNADIFFAREA                          0.160 LAYER ME3 ;
 ANTENNADIFFAREA                          0.160 LAYER ME4 ;
 ANTENNAMAXAREACAR                       48.755 LAYER ME2 ;
 ANTENNAMAXAREACAR                       58.014 LAYER ME3 ;
 ANTENNAMAXAREACAR                       67.273 LAYER ME4 ;
END DI97
PIN DO96
  DIRECTION OUTPUT ;
 PORT
  LAYER ME4 ;
  RECT 2039.200 0.000 2040.000 1.000 ;
  LAYER ME3 ;
  RECT 2039.200 0.000 2040.000 1.000 ;
  LAYER ME2 ;
  RECT 2039.200 0.000 2040.000 1.000 ;
  LAYER ME1 ;
  RECT 2039.200 0.000 2040.000 1.000 ;
 END
 ANTENNAPARTIALMETALAREA                  4.168 LAYER ME2 ;
 ANTENNADIFFAREA                          5.472 LAYER ME2 ;
 ANTENNADIFFAREA                          5.472 LAYER ME3 ;
 ANTENNADIFFAREA                          5.472 LAYER ME4 ;
END DO96
PIN WEB6
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 2026.400 0.000 2027.200 1.000 ;
  LAYER ME3 ;
  RECT 2026.400 0.000 2027.200 1.000 ;
  LAYER ME2 ;
  RECT 2026.400 0.000 2027.200 1.000 ;
  LAYER ME1 ;
  RECT 2026.400 0.000 2027.200 1.000 ;
 END
 ANTENNAPARTIALMETALAREA                  2.836 LAYER ME2 ;
 ANTENNAGATEAREA                          0.072 LAYER ME2 ;
 ANTENNAGATEAREA                          0.072 LAYER ME3 ;
 ANTENNAGATEAREA                          0.072 LAYER ME4 ;
 ANTENNADIFFAREA                          0.160 LAYER ME2 ;
 ANTENNADIFFAREA                          0.160 LAYER ME3 ;
 ANTENNADIFFAREA                          0.160 LAYER ME4 ;
 ANTENNAMAXAREACAR                       54.400 LAYER ME2 ;
 ANTENNAMAXAREACAR                       65.511 LAYER ME3 ;
 ANTENNAMAXAREACAR                       76.622 LAYER ME4 ;
END WEB6
PIN DI96
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 2024.800 0.000 2025.600 1.000 ;
  LAYER ME3 ;
  RECT 2024.800 0.000 2025.600 1.000 ;
  LAYER ME2 ;
  RECT 2024.800 0.000 2025.600 1.000 ;
  LAYER ME1 ;
  RECT 2024.800 0.000 2025.600 1.000 ;
 END
 ANTENNAPARTIALMETALAREA                  3.134 LAYER ME2 ;
 ANTENNAGATEAREA                          0.086 LAYER ME2 ;
 ANTENNAGATEAREA                          0.086 LAYER ME3 ;
 ANTENNAGATEAREA                          0.086 LAYER ME4 ;
 ANTENNADIFFAREA                          0.160 LAYER ME2 ;
 ANTENNADIFFAREA                          0.160 LAYER ME3 ;
 ANTENNADIFFAREA                          0.160 LAYER ME4 ;
 ANTENNAMAXAREACAR                       48.616 LAYER ME2 ;
 ANTENNAMAXAREACAR                       57.875 LAYER ME3 ;
 ANTENNAMAXAREACAR                       67.134 LAYER ME4 ;
END DI96
PIN DO95
  DIRECTION OUTPUT ;
 PORT
  LAYER ME4 ;
  RECT 2018.400 0.000 2019.200 1.000 ;
  LAYER ME3 ;
  RECT 2018.400 0.000 2019.200 1.000 ;
  LAYER ME2 ;
  RECT 2018.400 0.000 2019.200 1.000 ;
  LAYER ME1 ;
  RECT 2018.400 0.000 2019.200 1.000 ;
 END
 ANTENNAPARTIALMETALAREA                  4.168 LAYER ME2 ;
 ANTENNADIFFAREA                          5.472 LAYER ME2 ;
 ANTENNADIFFAREA                          5.472 LAYER ME3 ;
 ANTENNADIFFAREA                          5.472 LAYER ME4 ;
END DO95
PIN DI95
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 2003.600 0.000 2004.400 1.000 ;
  LAYER ME3 ;
  RECT 2003.600 0.000 2004.400 1.000 ;
  LAYER ME2 ;
  RECT 2003.600 0.000 2004.400 1.000 ;
  LAYER ME1 ;
  RECT 2003.600 0.000 2004.400 1.000 ;
 END
 ANTENNAPARTIALMETALAREA                  3.122 LAYER ME2 ;
 ANTENNAGATEAREA                          0.086 LAYER ME2 ;
 ANTENNAGATEAREA                          0.086 LAYER ME3 ;
 ANTENNAGATEAREA                          0.086 LAYER ME4 ;
 ANTENNADIFFAREA                          0.160 LAYER ME2 ;
 ANTENNADIFFAREA                          0.160 LAYER ME3 ;
 ANTENNADIFFAREA                          0.160 LAYER ME4 ;
 ANTENNAMAXAREACAR                       48.477 LAYER ME2 ;
 ANTENNAMAXAREACAR                       57.736 LAYER ME3 ;
 ANTENNAMAXAREACAR                       66.995 LAYER ME4 ;
END DI95
PIN DO94
  DIRECTION OUTPUT ;
 PORT
  LAYER ME4 ;
  RECT 1998.400 0.000 1999.200 1.000 ;
  LAYER ME3 ;
  RECT 1998.400 0.000 1999.200 1.000 ;
  LAYER ME2 ;
  RECT 1998.400 0.000 1999.200 1.000 ;
  LAYER ME1 ;
  RECT 1998.400 0.000 1999.200 1.000 ;
 END
 ANTENNAPARTIALMETALAREA                  4.144 LAYER ME2 ;
 ANTENNADIFFAREA                          5.472 LAYER ME2 ;
 ANTENNADIFFAREA                          5.472 LAYER ME3 ;
 ANTENNADIFFAREA                          5.472 LAYER ME4 ;
END DO94
PIN DI94
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 1983.600 0.000 1984.400 1.000 ;
  LAYER ME3 ;
  RECT 1983.600 0.000 1984.400 1.000 ;
  LAYER ME2 ;
  RECT 1983.600 0.000 1984.400 1.000 ;
  LAYER ME1 ;
  RECT 1983.600 0.000 1984.400 1.000 ;
 END
 ANTENNAPARTIALMETALAREA                  3.154 LAYER ME2 ;
 ANTENNAGATEAREA                          0.086 LAYER ME2 ;
 ANTENNAGATEAREA                          0.086 LAYER ME3 ;
 ANTENNAGATEAREA                          0.086 LAYER ME4 ;
 ANTENNADIFFAREA                          0.160 LAYER ME2 ;
 ANTENNADIFFAREA                          0.160 LAYER ME3 ;
 ANTENNADIFFAREA                          0.160 LAYER ME4 ;
 ANTENNAMAXAREACAR                       48.847 LAYER ME2 ;
 ANTENNAMAXAREACAR                       58.106 LAYER ME3 ;
 ANTENNAMAXAREACAR                       67.366 LAYER ME4 ;
END DI94
PIN DO93
  DIRECTION OUTPUT ;
 PORT
  LAYER ME4 ;
  RECT 1977.200 0.000 1978.000 1.000 ;
  LAYER ME3 ;
  RECT 1977.200 0.000 1978.000 1.000 ;
  LAYER ME2 ;
  RECT 1977.200 0.000 1978.000 1.000 ;
  LAYER ME1 ;
  RECT 1977.200 0.000 1978.000 1.000 ;
 END
 ANTENNAPARTIALMETALAREA                  4.168 LAYER ME2 ;
 ANTENNADIFFAREA                          5.472 LAYER ME2 ;
 ANTENNADIFFAREA                          5.472 LAYER ME3 ;
 ANTENNADIFFAREA                          5.472 LAYER ME4 ;
END DO93
PIN DI93
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 1962.800 0.000 1963.600 1.000 ;
  LAYER ME3 ;
  RECT 1962.800 0.000 1963.600 1.000 ;
  LAYER ME2 ;
  RECT 1962.800 0.000 1963.600 1.000 ;
  LAYER ME1 ;
  RECT 1962.800 0.000 1963.600 1.000 ;
 END
 ANTENNAPARTIALMETALAREA                  3.134 LAYER ME2 ;
 ANTENNAGATEAREA                          0.086 LAYER ME2 ;
 ANTENNAGATEAREA                          0.086 LAYER ME3 ;
 ANTENNAGATEAREA                          0.086 LAYER ME4 ;
 ANTENNADIFFAREA                          0.160 LAYER ME2 ;
 ANTENNADIFFAREA                          0.160 LAYER ME3 ;
 ANTENNADIFFAREA                          0.160 LAYER ME4 ;
 ANTENNAMAXAREACAR                       48.616 LAYER ME2 ;
 ANTENNAMAXAREACAR                       57.875 LAYER ME3 ;
 ANTENNAMAXAREACAR                       67.134 LAYER ME4 ;
END DI93
PIN DO92
  DIRECTION OUTPUT ;
 PORT
  LAYER ME4 ;
  RECT 1957.600 0.000 1958.400 1.000 ;
  LAYER ME3 ;
  RECT 1957.600 0.000 1958.400 1.000 ;
  LAYER ME2 ;
  RECT 1957.600 0.000 1958.400 1.000 ;
  LAYER ME1 ;
  RECT 1957.600 0.000 1958.400 1.000 ;
 END
 ANTENNAPARTIALMETALAREA                  4.160 LAYER ME2 ;
 ANTENNADIFFAREA                          5.472 LAYER ME2 ;
 ANTENNADIFFAREA                          5.472 LAYER ME3 ;
 ANTENNADIFFAREA                          5.472 LAYER ME4 ;
END DO92
PIN DI92
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 1942.800 0.000 1943.600 1.000 ;
  LAYER ME3 ;
  RECT 1942.800 0.000 1943.600 1.000 ;
  LAYER ME2 ;
  RECT 1942.800 0.000 1943.600 1.000 ;
  LAYER ME1 ;
  RECT 1942.800 0.000 1943.600 1.000 ;
 END
 ANTENNAPARTIALMETALAREA                  3.130 LAYER ME2 ;
 ANTENNAGATEAREA                          0.086 LAYER ME2 ;
 ANTENNAGATEAREA                          0.086 LAYER ME3 ;
 ANTENNAGATEAREA                          0.086 LAYER ME4 ;
 ANTENNADIFFAREA                          0.160 LAYER ME2 ;
 ANTENNADIFFAREA                          0.160 LAYER ME3 ;
 ANTENNADIFFAREA                          0.160 LAYER ME4 ;
 ANTENNAMAXAREACAR                       48.569 LAYER ME2 ;
 ANTENNAMAXAREACAR                       57.829 LAYER ME3 ;
 ANTENNAMAXAREACAR                       67.088 LAYER ME4 ;
END DI92
PIN DO91
  DIRECTION OUTPUT ;
 PORT
  LAYER ME4 ;
  RECT 1936.400 0.000 1937.200 1.000 ;
  LAYER ME3 ;
  RECT 1936.400 0.000 1937.200 1.000 ;
  LAYER ME2 ;
  RECT 1936.400 0.000 1937.200 1.000 ;
  LAYER ME1 ;
  RECT 1936.400 0.000 1937.200 1.000 ;
 END
 ANTENNAPARTIALMETALAREA                  4.144 LAYER ME2 ;
 ANTENNADIFFAREA                          5.472 LAYER ME2 ;
 ANTENNADIFFAREA                          5.472 LAYER ME3 ;
 ANTENNADIFFAREA                          5.472 LAYER ME4 ;
END DO91
PIN DI91
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 1921.600 0.000 1922.400 1.000 ;
  LAYER ME3 ;
  RECT 1921.600 0.000 1922.400 1.000 ;
  LAYER ME2 ;
  RECT 1921.600 0.000 1922.400 1.000 ;
  LAYER ME1 ;
  RECT 1921.600 0.000 1922.400 1.000 ;
 END
 ANTENNAPARTIALMETALAREA                  3.154 LAYER ME2 ;
 ANTENNAGATEAREA                          0.086 LAYER ME2 ;
 ANTENNAGATEAREA                          0.086 LAYER ME3 ;
 ANTENNAGATEAREA                          0.086 LAYER ME4 ;
 ANTENNADIFFAREA                          0.160 LAYER ME2 ;
 ANTENNADIFFAREA                          0.160 LAYER ME3 ;
 ANTENNADIFFAREA                          0.160 LAYER ME4 ;
 ANTENNAMAXAREACAR                       48.847 LAYER ME2 ;
 ANTENNAMAXAREACAR                       58.106 LAYER ME3 ;
 ANTENNAMAXAREACAR                       67.366 LAYER ME4 ;
END DI91
PIN DO90
  DIRECTION OUTPUT ;
 PORT
  LAYER ME4 ;
  RECT 1916.400 0.000 1917.200 1.000 ;
  LAYER ME3 ;
  RECT 1916.400 0.000 1917.200 1.000 ;
  LAYER ME2 ;
  RECT 1916.400 0.000 1917.200 1.000 ;
  LAYER ME1 ;
  RECT 1916.400 0.000 1917.200 1.000 ;
 END
 ANTENNAPARTIALMETALAREA                  4.176 LAYER ME2 ;
 ANTENNADIFFAREA                          5.472 LAYER ME2 ;
 ANTENNADIFFAREA                          5.472 LAYER ME3 ;
 ANTENNADIFFAREA                          5.472 LAYER ME4 ;
END DO90
PIN DI90
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 1902.000 0.000 1902.800 1.000 ;
  LAYER ME3 ;
  RECT 1902.000 0.000 1902.800 1.000 ;
  LAYER ME2 ;
  RECT 1902.000 0.000 1902.800 1.000 ;
  LAYER ME1 ;
  RECT 1902.000 0.000 1902.800 1.000 ;
 END
 ANTENNAPARTIALMETALAREA                  3.126 LAYER ME2 ;
 ANTENNAGATEAREA                          0.086 LAYER ME2 ;
 ANTENNAGATEAREA                          0.086 LAYER ME3 ;
 ANTENNAGATEAREA                          0.086 LAYER ME4 ;
 ANTENNADIFFAREA                          0.160 LAYER ME2 ;
 ANTENNADIFFAREA                          0.160 LAYER ME3 ;
 ANTENNADIFFAREA                          0.160 LAYER ME4 ;
 ANTENNAMAXAREACAR                       48.523 LAYER ME2 ;
 ANTENNAMAXAREACAR                       57.782 LAYER ME3 ;
 ANTENNAMAXAREACAR                       67.042 LAYER ME4 ;
END DI90
PIN DO89
  DIRECTION OUTPUT ;
 PORT
  LAYER ME4 ;
  RECT 1895.600 0.000 1896.400 1.000 ;
  LAYER ME3 ;
  RECT 1895.600 0.000 1896.400 1.000 ;
  LAYER ME2 ;
  RECT 1895.600 0.000 1896.400 1.000 ;
  LAYER ME1 ;
  RECT 1895.600 0.000 1896.400 1.000 ;
 END
 ANTENNAPARTIALMETALAREA                  4.160 LAYER ME2 ;
 ANTENNADIFFAREA                          5.472 LAYER ME2 ;
 ANTENNADIFFAREA                          5.472 LAYER ME3 ;
 ANTENNADIFFAREA                          5.472 LAYER ME4 ;
END DO89
PIN DI89
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 1880.800 0.000 1881.600 1.000 ;
  LAYER ME3 ;
  RECT 1880.800 0.000 1881.600 1.000 ;
  LAYER ME2 ;
  RECT 1880.800 0.000 1881.600 1.000 ;
  LAYER ME1 ;
  RECT 1880.800 0.000 1881.600 1.000 ;
 END
 ANTENNAPARTIALMETALAREA                  3.130 LAYER ME2 ;
 ANTENNAGATEAREA                          0.086 LAYER ME2 ;
 ANTENNAGATEAREA                          0.086 LAYER ME3 ;
 ANTENNAGATEAREA                          0.086 LAYER ME4 ;
 ANTENNADIFFAREA                          0.160 LAYER ME2 ;
 ANTENNADIFFAREA                          0.160 LAYER ME3 ;
 ANTENNADIFFAREA                          0.160 LAYER ME4 ;
 ANTENNAMAXAREACAR                       48.569 LAYER ME2 ;
 ANTENNAMAXAREACAR                       57.829 LAYER ME3 ;
 ANTENNAMAXAREACAR                       67.088 LAYER ME4 ;
END DI89
PIN DO88
  DIRECTION OUTPUT ;
 PORT
  LAYER ME4 ;
  RECT 1875.600 0.000 1876.400 1.000 ;
  LAYER ME3 ;
  RECT 1875.600 0.000 1876.400 1.000 ;
  LAYER ME2 ;
  RECT 1875.600 0.000 1876.400 1.000 ;
  LAYER ME1 ;
  RECT 1875.600 0.000 1876.400 1.000 ;
 END
 ANTENNAPARTIALMETALAREA                  4.152 LAYER ME2 ;
 ANTENNADIFFAREA                          5.472 LAYER ME2 ;
 ANTENNADIFFAREA                          5.472 LAYER ME3 ;
 ANTENNADIFFAREA                          5.472 LAYER ME4 ;
END DO88
PIN DI88
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 1861.200 0.000 1862.000 1.000 ;
  LAYER ME3 ;
  RECT 1861.200 0.000 1862.000 1.000 ;
  LAYER ME2 ;
  RECT 1861.200 0.000 1862.000 1.000 ;
  LAYER ME1 ;
  RECT 1861.200 0.000 1862.000 1.000 ;
 END
 ANTENNAPARTIALMETALAREA                  3.150 LAYER ME2 ;
 ANTENNAGATEAREA                          0.086 LAYER ME2 ;
 ANTENNAGATEAREA                          0.086 LAYER ME3 ;
 ANTENNAGATEAREA                          0.086 LAYER ME4 ;
 ANTENNADIFFAREA                          0.160 LAYER ME2 ;
 ANTENNADIFFAREA                          0.160 LAYER ME3 ;
 ANTENNADIFFAREA                          0.160 LAYER ME4 ;
 ANTENNAMAXAREACAR                       48.801 LAYER ME2 ;
 ANTENNAMAXAREACAR                       58.060 LAYER ME3 ;
 ANTENNAMAXAREACAR                       67.319 LAYER ME4 ;
END DI88
PIN DO87
  DIRECTION OUTPUT ;
 PORT
  LAYER ME4 ;
  RECT 1854.400 0.000 1855.200 1.000 ;
  LAYER ME3 ;
  RECT 1854.400 0.000 1855.200 1.000 ;
  LAYER ME2 ;
  RECT 1854.400 0.000 1855.200 1.000 ;
  LAYER ME1 ;
  RECT 1854.400 0.000 1855.200 1.000 ;
 END
 ANTENNAPARTIALMETALAREA                  4.176 LAYER ME2 ;
 ANTENNADIFFAREA                          5.472 LAYER ME2 ;
 ANTENNADIFFAREA                          5.472 LAYER ME3 ;
 ANTENNADIFFAREA                          5.472 LAYER ME4 ;
END DO87
PIN DI87
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 1840.000 0.000 1840.800 1.000 ;
  LAYER ME3 ;
  RECT 1840.000 0.000 1840.800 1.000 ;
  LAYER ME2 ;
  RECT 1840.000 0.000 1840.800 1.000 ;
  LAYER ME1 ;
  RECT 1840.000 0.000 1840.800 1.000 ;
 END
 ANTENNAPARTIALMETALAREA                  3.126 LAYER ME2 ;
 ANTENNAGATEAREA                          0.086 LAYER ME2 ;
 ANTENNAGATEAREA                          0.086 LAYER ME3 ;
 ANTENNAGATEAREA                          0.086 LAYER ME4 ;
 ANTENNADIFFAREA                          0.160 LAYER ME2 ;
 ANTENNADIFFAREA                          0.160 LAYER ME3 ;
 ANTENNADIFFAREA                          0.160 LAYER ME4 ;
 ANTENNAMAXAREACAR                       48.523 LAYER ME2 ;
 ANTENNAMAXAREACAR                       57.782 LAYER ME3 ;
 ANTENNAMAXAREACAR                       67.042 LAYER ME4 ;
END DI87
PIN DO86
  DIRECTION OUTPUT ;
 PORT
  LAYER ME4 ;
  RECT 1834.800 0.000 1835.600 1.000 ;
  LAYER ME3 ;
  RECT 1834.800 0.000 1835.600 1.000 ;
  LAYER ME2 ;
  RECT 1834.800 0.000 1835.600 1.000 ;
  LAYER ME1 ;
  RECT 1834.800 0.000 1835.600 1.000 ;
 END
 ANTENNAPARTIALMETALAREA                  4.152 LAYER ME2 ;
 ANTENNADIFFAREA                          5.472 LAYER ME2 ;
 ANTENNADIFFAREA                          5.472 LAYER ME3 ;
 ANTENNADIFFAREA                          5.472 LAYER ME4 ;
END DO86
PIN DI86
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 1820.000 0.000 1820.800 1.000 ;
  LAYER ME3 ;
  RECT 1820.000 0.000 1820.800 1.000 ;
  LAYER ME2 ;
  RECT 1820.000 0.000 1820.800 1.000 ;
  LAYER ME1 ;
  RECT 1820.000 0.000 1820.800 1.000 ;
 END
 ANTENNAPARTIALMETALAREA                  3.138 LAYER ME2 ;
 ANTENNAGATEAREA                          0.086 LAYER ME2 ;
 ANTENNAGATEAREA                          0.086 LAYER ME3 ;
 ANTENNAGATEAREA                          0.086 LAYER ME4 ;
 ANTENNADIFFAREA                          0.160 LAYER ME2 ;
 ANTENNADIFFAREA                          0.160 LAYER ME3 ;
 ANTENNADIFFAREA                          0.160 LAYER ME4 ;
 ANTENNAMAXAREACAR                       48.662 LAYER ME2 ;
 ANTENNAMAXAREACAR                       57.921 LAYER ME3 ;
 ANTENNAMAXAREACAR                       67.181 LAYER ME4 ;
END DI86
PIN DO85
  DIRECTION OUTPUT ;
 PORT
  LAYER ME4 ;
  RECT 1813.600 0.000 1814.400 1.000 ;
  LAYER ME3 ;
  RECT 1813.600 0.000 1814.400 1.000 ;
  LAYER ME2 ;
  RECT 1813.600 0.000 1814.400 1.000 ;
  LAYER ME1 ;
  RECT 1813.600 0.000 1814.400 1.000 ;
 END
 ANTENNAPARTIALMETALAREA                  4.152 LAYER ME2 ;
 ANTENNADIFFAREA                          5.472 LAYER ME2 ;
 ANTENNADIFFAREA                          5.472 LAYER ME3 ;
 ANTENNADIFFAREA                          5.472 LAYER ME4 ;
END DO85
PIN DI85
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 1799.200 0.000 1800.000 1.000 ;
  LAYER ME3 ;
  RECT 1799.200 0.000 1800.000 1.000 ;
  LAYER ME2 ;
  RECT 1799.200 0.000 1800.000 1.000 ;
  LAYER ME1 ;
  RECT 1799.200 0.000 1800.000 1.000 ;
 END
 ANTENNAPARTIALMETALAREA                  3.150 LAYER ME2 ;
 ANTENNAGATEAREA                          0.086 LAYER ME2 ;
 ANTENNAGATEAREA                          0.086 LAYER ME3 ;
 ANTENNAGATEAREA                          0.086 LAYER ME4 ;
 ANTENNADIFFAREA                          0.160 LAYER ME2 ;
 ANTENNADIFFAREA                          0.160 LAYER ME3 ;
 ANTENNADIFFAREA                          0.160 LAYER ME4 ;
 ANTENNAMAXAREACAR                       48.801 LAYER ME2 ;
 ANTENNAMAXAREACAR                       58.060 LAYER ME3 ;
 ANTENNAMAXAREACAR                       67.319 LAYER ME4 ;
END DI85
PIN DO84
  DIRECTION OUTPUT ;
 PORT
  LAYER ME4 ;
  RECT 1794.000 0.000 1794.800 1.000 ;
  LAYER ME3 ;
  RECT 1794.000 0.000 1794.800 1.000 ;
  LAYER ME2 ;
  RECT 1794.000 0.000 1794.800 1.000 ;
  LAYER ME1 ;
  RECT 1794.000 0.000 1794.800 1.000 ;
 END
 ANTENNAPARTIALMETALAREA                  4.176 LAYER ME2 ;
 ANTENNADIFFAREA                          5.472 LAYER ME2 ;
 ANTENNADIFFAREA                          5.472 LAYER ME3 ;
 ANTENNADIFFAREA                          5.472 LAYER ME4 ;
END DO84
PIN DI84
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 1779.200 0.000 1780.000 1.000 ;
  LAYER ME3 ;
  RECT 1779.200 0.000 1780.000 1.000 ;
  LAYER ME2 ;
  RECT 1779.200 0.000 1780.000 1.000 ;
  LAYER ME1 ;
  RECT 1779.200 0.000 1780.000 1.000 ;
 END
 ANTENNAPARTIALMETALAREA                  3.118 LAYER ME2 ;
 ANTENNAGATEAREA                          0.086 LAYER ME2 ;
 ANTENNAGATEAREA                          0.086 LAYER ME3 ;
 ANTENNAGATEAREA                          0.086 LAYER ME4 ;
 ANTENNADIFFAREA                          0.160 LAYER ME2 ;
 ANTENNADIFFAREA                          0.160 LAYER ME3 ;
 ANTENNADIFFAREA                          0.160 LAYER ME4 ;
 ANTENNAMAXAREACAR                       48.431 LAYER ME2 ;
 ANTENNAMAXAREACAR                       57.690 LAYER ME3 ;
 ANTENNAMAXAREACAR                       66.949 LAYER ME4 ;
END DI84
PIN DO83
  DIRECTION OUTPUT ;
 PORT
  LAYER ME4 ;
  RECT 1772.800 0.000 1773.600 1.000 ;
  LAYER ME3 ;
  RECT 1772.800 0.000 1773.600 1.000 ;
  LAYER ME2 ;
  RECT 1772.800 0.000 1773.600 1.000 ;
  LAYER ME1 ;
  RECT 1772.800 0.000 1773.600 1.000 ;
 END
 ANTENNAPARTIALMETALAREA                  4.152 LAYER ME2 ;
 ANTENNADIFFAREA                          5.472 LAYER ME2 ;
 ANTENNADIFFAREA                          5.472 LAYER ME3 ;
 ANTENNADIFFAREA                          5.472 LAYER ME4 ;
END DO83
PIN DI83
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 1758.000 0.000 1758.800 1.000 ;
  LAYER ME3 ;
  RECT 1758.000 0.000 1758.800 1.000 ;
  LAYER ME2 ;
  RECT 1758.000 0.000 1758.800 1.000 ;
  LAYER ME1 ;
  RECT 1758.000 0.000 1758.800 1.000 ;
 END
 ANTENNAPARTIALMETALAREA                  3.138 LAYER ME2 ;
 ANTENNAGATEAREA                          0.086 LAYER ME2 ;
 ANTENNAGATEAREA                          0.086 LAYER ME3 ;
 ANTENNAGATEAREA                          0.086 LAYER ME4 ;
 ANTENNADIFFAREA                          0.160 LAYER ME2 ;
 ANTENNADIFFAREA                          0.160 LAYER ME3 ;
 ANTENNADIFFAREA                          0.160 LAYER ME4 ;
 ANTENNAMAXAREACAR                       48.662 LAYER ME2 ;
 ANTENNAMAXAREACAR                       57.921 LAYER ME3 ;
 ANTENNAMAXAREACAR                       67.181 LAYER ME4 ;
END DI83
PIN DO82
  DIRECTION OUTPUT ;
 PORT
  LAYER ME4 ;
  RECT 1752.800 0.000 1753.600 1.000 ;
  LAYER ME3 ;
  RECT 1752.800 0.000 1753.600 1.000 ;
  LAYER ME2 ;
  RECT 1752.800 0.000 1753.600 1.000 ;
  LAYER ME1 ;
  RECT 1752.800 0.000 1753.600 1.000 ;
 END
 ANTENNAPARTIALMETALAREA                  4.160 LAYER ME2 ;
 ANTENNADIFFAREA                          5.472 LAYER ME2 ;
 ANTENNADIFFAREA                          5.472 LAYER ME3 ;
 ANTENNADIFFAREA                          5.472 LAYER ME4 ;
END DO82
PIN DI82
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 1738.400 0.000 1739.200 1.000 ;
  LAYER ME3 ;
  RECT 1738.400 0.000 1739.200 1.000 ;
  LAYER ME2 ;
  RECT 1738.400 0.000 1739.200 1.000 ;
  LAYER ME1 ;
  RECT 1738.400 0.000 1739.200 1.000 ;
 END
 ANTENNAPARTIALMETALAREA                  3.142 LAYER ME2 ;
 ANTENNAGATEAREA                          0.086 LAYER ME2 ;
 ANTENNAGATEAREA                          0.086 LAYER ME3 ;
 ANTENNAGATEAREA                          0.086 LAYER ME4 ;
 ANTENNADIFFAREA                          0.160 LAYER ME2 ;
 ANTENNADIFFAREA                          0.160 LAYER ME3 ;
 ANTENNADIFFAREA                          0.160 LAYER ME4 ;
 ANTENNAMAXAREACAR                       48.708 LAYER ME2 ;
 ANTENNAMAXAREACAR                       57.968 LAYER ME3 ;
 ANTENNAMAXAREACAR                       67.227 LAYER ME4 ;
END DI82
PIN DO81
  DIRECTION OUTPUT ;
 PORT
  LAYER ME4 ;
  RECT 1732.000 0.000 1732.800 1.000 ;
  LAYER ME3 ;
  RECT 1732.000 0.000 1732.800 1.000 ;
  LAYER ME2 ;
  RECT 1732.000 0.000 1732.800 1.000 ;
  LAYER ME1 ;
  RECT 1732.000 0.000 1732.800 1.000 ;
 END
 ANTENNAPARTIALMETALAREA                  4.176 LAYER ME2 ;
 ANTENNADIFFAREA                          5.472 LAYER ME2 ;
 ANTENNADIFFAREA                          5.472 LAYER ME3 ;
 ANTENNADIFFAREA                          5.472 LAYER ME4 ;
END DO81
PIN DI81
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 1717.200 0.000 1718.000 1.000 ;
  LAYER ME3 ;
  RECT 1717.200 0.000 1718.000 1.000 ;
  LAYER ME2 ;
  RECT 1717.200 0.000 1718.000 1.000 ;
  LAYER ME1 ;
  RECT 1717.200 0.000 1718.000 1.000 ;
 END
 ANTENNAPARTIALMETALAREA                  3.118 LAYER ME2 ;
 ANTENNAGATEAREA                          0.086 LAYER ME2 ;
 ANTENNAGATEAREA                          0.086 LAYER ME3 ;
 ANTENNAGATEAREA                          0.086 LAYER ME4 ;
 ANTENNADIFFAREA                          0.160 LAYER ME2 ;
 ANTENNADIFFAREA                          0.160 LAYER ME3 ;
 ANTENNADIFFAREA                          0.160 LAYER ME4 ;
 ANTENNAMAXAREACAR                       48.431 LAYER ME2 ;
 ANTENNAMAXAREACAR                       57.690 LAYER ME3 ;
 ANTENNAMAXAREACAR                       66.949 LAYER ME4 ;
END DI81
PIN DO80
  DIRECTION OUTPUT ;
 PORT
  LAYER ME4 ;
  RECT 1712.000 0.000 1712.800 1.000 ;
  LAYER ME3 ;
  RECT 1712.000 0.000 1712.800 1.000 ;
  LAYER ME2 ;
  RECT 1712.000 0.000 1712.800 1.000 ;
  LAYER ME1 ;
  RECT 1712.000 0.000 1712.800 1.000 ;
 END
 ANTENNAPARTIALMETALAREA                  4.144 LAYER ME2 ;
 ANTENNADIFFAREA                          5.472 LAYER ME2 ;
 ANTENNADIFFAREA                          5.472 LAYER ME3 ;
 ANTENNADIFFAREA                          5.472 LAYER ME4 ;
END DO80
PIN WEB5
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 1699.200 0.000 1700.000 1.000 ;
  LAYER ME3 ;
  RECT 1699.200 0.000 1700.000 1.000 ;
  LAYER ME2 ;
  RECT 1699.200 0.000 1700.000 1.000 ;
  LAYER ME1 ;
  RECT 1699.200 0.000 1700.000 1.000 ;
 END
 ANTENNAPARTIALMETALAREA                  2.856 LAYER ME2 ;
 ANTENNAGATEAREA                          0.072 LAYER ME2 ;
 ANTENNAGATEAREA                          0.072 LAYER ME3 ;
 ANTENNAGATEAREA                          0.072 LAYER ME4 ;
 ANTENNADIFFAREA                          0.160 LAYER ME2 ;
 ANTENNADIFFAREA                          0.160 LAYER ME3 ;
 ANTENNADIFFAREA                          0.160 LAYER ME4 ;
 ANTENNAMAXAREACAR                       54.678 LAYER ME2 ;
 ANTENNAMAXAREACAR                       65.789 LAYER ME3 ;
 ANTENNAMAXAREACAR                       76.900 LAYER ME4 ;
END WEB5
PIN DI80
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 1697.200 0.000 1698.000 1.000 ;
  LAYER ME3 ;
  RECT 1697.200 0.000 1698.000 1.000 ;
  LAYER ME2 ;
  RECT 1697.200 0.000 1698.000 1.000 ;
  LAYER ME1 ;
  RECT 1697.200 0.000 1698.000 1.000 ;
 END
 ANTENNAPARTIALMETALAREA                  3.146 LAYER ME2 ;
 ANTENNAGATEAREA                          0.086 LAYER ME2 ;
 ANTENNAGATEAREA                          0.086 LAYER ME3 ;
 ANTENNAGATEAREA                          0.086 LAYER ME4 ;
 ANTENNADIFFAREA                          0.160 LAYER ME2 ;
 ANTENNADIFFAREA                          0.160 LAYER ME3 ;
 ANTENNADIFFAREA                          0.160 LAYER ME4 ;
 ANTENNAMAXAREACAR                       48.755 LAYER ME2 ;
 ANTENNAMAXAREACAR                       58.014 LAYER ME3 ;
 ANTENNAMAXAREACAR                       67.273 LAYER ME4 ;
END DI80
PIN DO79
  DIRECTION OUTPUT ;
 PORT
  LAYER ME4 ;
  RECT 1690.800 0.000 1691.600 1.000 ;
  LAYER ME3 ;
  RECT 1690.800 0.000 1691.600 1.000 ;
  LAYER ME2 ;
  RECT 1690.800 0.000 1691.600 1.000 ;
  LAYER ME1 ;
  RECT 1690.800 0.000 1691.600 1.000 ;
 END
 ANTENNAPARTIALMETALAREA                  4.160 LAYER ME2 ;
 ANTENNADIFFAREA                          5.472 LAYER ME2 ;
 ANTENNADIFFAREA                          5.472 LAYER ME3 ;
 ANTENNADIFFAREA                          5.472 LAYER ME4 ;
END DO79
PIN DI79
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 1676.400 0.000 1677.200 1.000 ;
  LAYER ME3 ;
  RECT 1676.400 0.000 1677.200 1.000 ;
  LAYER ME2 ;
  RECT 1676.400 0.000 1677.200 1.000 ;
  LAYER ME1 ;
  RECT 1676.400 0.000 1677.200 1.000 ;
 END
 ANTENNAPARTIALMETALAREA                  3.142 LAYER ME2 ;
 ANTENNAGATEAREA                          0.086 LAYER ME2 ;
 ANTENNAGATEAREA                          0.086 LAYER ME3 ;
 ANTENNAGATEAREA                          0.086 LAYER ME4 ;
 ANTENNADIFFAREA                          0.160 LAYER ME2 ;
 ANTENNADIFFAREA                          0.160 LAYER ME3 ;
 ANTENNADIFFAREA                          0.160 LAYER ME4 ;
 ANTENNAMAXAREACAR                       48.708 LAYER ME2 ;
 ANTENNAMAXAREACAR                       57.968 LAYER ME3 ;
 ANTENNAMAXAREACAR                       67.227 LAYER ME4 ;
END DI79
PIN DO78
  DIRECTION OUTPUT ;
 PORT
  LAYER ME4 ;
  RECT 1671.200 0.000 1672.000 1.000 ;
  LAYER ME3 ;
  RECT 1671.200 0.000 1672.000 1.000 ;
  LAYER ME2 ;
  RECT 1671.200 0.000 1672.000 1.000 ;
  LAYER ME1 ;
  RECT 1671.200 0.000 1672.000 1.000 ;
 END
 ANTENNAPARTIALMETALAREA                  4.168 LAYER ME2 ;
 ANTENNADIFFAREA                          5.472 LAYER ME2 ;
 ANTENNADIFFAREA                          5.472 LAYER ME3 ;
 ANTENNADIFFAREA                          5.472 LAYER ME4 ;
END DO78
PIN DI78
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 1656.400 0.000 1657.200 1.000 ;
  LAYER ME3 ;
  RECT 1656.400 0.000 1657.200 1.000 ;
  LAYER ME2 ;
  RECT 1656.400 0.000 1657.200 1.000 ;
  LAYER ME1 ;
  RECT 1656.400 0.000 1657.200 1.000 ;
 END
 ANTENNAPARTIALMETALAREA                  3.122 LAYER ME2 ;
 ANTENNAGATEAREA                          0.086 LAYER ME2 ;
 ANTENNAGATEAREA                          0.086 LAYER ME3 ;
 ANTENNAGATEAREA                          0.086 LAYER ME4 ;
 ANTENNADIFFAREA                          0.160 LAYER ME2 ;
 ANTENNADIFFAREA                          0.160 LAYER ME3 ;
 ANTENNADIFFAREA                          0.160 LAYER ME4 ;
 ANTENNAMAXAREACAR                       48.477 LAYER ME2 ;
 ANTENNAMAXAREACAR                       57.736 LAYER ME3 ;
 ANTENNAMAXAREACAR                       66.995 LAYER ME4 ;
END DI78
PIN DO77
  DIRECTION OUTPUT ;
 PORT
  LAYER ME4 ;
  RECT 1650.000 0.000 1650.800 1.000 ;
  LAYER ME3 ;
  RECT 1650.000 0.000 1650.800 1.000 ;
  LAYER ME2 ;
  RECT 1650.000 0.000 1650.800 1.000 ;
  LAYER ME1 ;
  RECT 1650.000 0.000 1650.800 1.000 ;
 END
 ANTENNAPARTIALMETALAREA                  4.144 LAYER ME2 ;
 ANTENNADIFFAREA                          5.472 LAYER ME2 ;
 ANTENNADIFFAREA                          5.472 LAYER ME3 ;
 ANTENNADIFFAREA                          5.472 LAYER ME4 ;
END DO77
PIN DI77
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 1635.200 0.000 1636.000 1.000 ;
  LAYER ME3 ;
  RECT 1635.200 0.000 1636.000 1.000 ;
  LAYER ME2 ;
  RECT 1635.200 0.000 1636.000 1.000 ;
  LAYER ME1 ;
  RECT 1635.200 0.000 1636.000 1.000 ;
 END
 ANTENNAPARTIALMETALAREA                  3.146 LAYER ME2 ;
 ANTENNAGATEAREA                          0.086 LAYER ME2 ;
 ANTENNAGATEAREA                          0.086 LAYER ME3 ;
 ANTENNAGATEAREA                          0.086 LAYER ME4 ;
 ANTENNADIFFAREA                          0.160 LAYER ME2 ;
 ANTENNADIFFAREA                          0.160 LAYER ME3 ;
 ANTENNADIFFAREA                          0.160 LAYER ME4 ;
 ANTENNAMAXAREACAR                       48.755 LAYER ME2 ;
 ANTENNAMAXAREACAR                       58.014 LAYER ME3 ;
 ANTENNAMAXAREACAR                       67.273 LAYER ME4 ;
END DI77
PIN DO76
  DIRECTION OUTPUT ;
 PORT
  LAYER ME4 ;
  RECT 1630.000 0.000 1630.800 1.000 ;
  LAYER ME3 ;
  RECT 1630.000 0.000 1630.800 1.000 ;
  LAYER ME2 ;
  RECT 1630.000 0.000 1630.800 1.000 ;
  LAYER ME1 ;
  RECT 1630.000 0.000 1630.800 1.000 ;
 END
 ANTENNAPARTIALMETALAREA                  4.168 LAYER ME2 ;
 ANTENNADIFFAREA                          5.472 LAYER ME2 ;
 ANTENNADIFFAREA                          5.472 LAYER ME3 ;
 ANTENNADIFFAREA                          5.472 LAYER ME4 ;
END DO76
PIN DI76
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 1615.600 0.000 1616.400 1.000 ;
  LAYER ME3 ;
  RECT 1615.600 0.000 1616.400 1.000 ;
  LAYER ME2 ;
  RECT 1615.600 0.000 1616.400 1.000 ;
  LAYER ME1 ;
  RECT 1615.600 0.000 1616.400 1.000 ;
 END
 ANTENNAPARTIALMETALAREA                  3.134 LAYER ME2 ;
 ANTENNAGATEAREA                          0.086 LAYER ME2 ;
 ANTENNAGATEAREA                          0.086 LAYER ME3 ;
 ANTENNAGATEAREA                          0.086 LAYER ME4 ;
 ANTENNADIFFAREA                          0.160 LAYER ME2 ;
 ANTENNADIFFAREA                          0.160 LAYER ME3 ;
 ANTENNADIFFAREA                          0.160 LAYER ME4 ;
 ANTENNAMAXAREACAR                       48.616 LAYER ME2 ;
 ANTENNAMAXAREACAR                       57.875 LAYER ME3 ;
 ANTENNAMAXAREACAR                       67.134 LAYER ME4 ;
END DI76
PIN DO75
  DIRECTION OUTPUT ;
 PORT
  LAYER ME4 ;
  RECT 1609.200 0.000 1610.000 1.000 ;
  LAYER ME3 ;
  RECT 1609.200 0.000 1610.000 1.000 ;
  LAYER ME2 ;
  RECT 1609.200 0.000 1610.000 1.000 ;
  LAYER ME1 ;
  RECT 1609.200 0.000 1610.000 1.000 ;
 END
 ANTENNAPARTIALMETALAREA                  4.168 LAYER ME2 ;
 ANTENNADIFFAREA                          5.472 LAYER ME2 ;
 ANTENNADIFFAREA                          5.472 LAYER ME3 ;
 ANTENNADIFFAREA                          5.472 LAYER ME4 ;
END DO75
PIN DI75
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 1594.400 0.000 1595.200 1.000 ;
  LAYER ME3 ;
  RECT 1594.400 0.000 1595.200 1.000 ;
  LAYER ME2 ;
  RECT 1594.400 0.000 1595.200 1.000 ;
  LAYER ME1 ;
  RECT 1594.400 0.000 1595.200 1.000 ;
 END
 ANTENNAPARTIALMETALAREA                  3.122 LAYER ME2 ;
 ANTENNAGATEAREA                          0.086 LAYER ME2 ;
 ANTENNAGATEAREA                          0.086 LAYER ME3 ;
 ANTENNAGATEAREA                          0.086 LAYER ME4 ;
 ANTENNADIFFAREA                          0.160 LAYER ME2 ;
 ANTENNADIFFAREA                          0.160 LAYER ME3 ;
 ANTENNADIFFAREA                          0.160 LAYER ME4 ;
 ANTENNAMAXAREACAR                       48.477 LAYER ME2 ;
 ANTENNAMAXAREACAR                       57.736 LAYER ME3 ;
 ANTENNAMAXAREACAR                       66.995 LAYER ME4 ;
END DI75
PIN DO74
  DIRECTION OUTPUT ;
 PORT
  LAYER ME4 ;
  RECT 1589.200 0.000 1590.000 1.000 ;
  LAYER ME3 ;
  RECT 1589.200 0.000 1590.000 1.000 ;
  LAYER ME2 ;
  RECT 1589.200 0.000 1590.000 1.000 ;
  LAYER ME1 ;
  RECT 1589.200 0.000 1590.000 1.000 ;
 END
 ANTENNAPARTIALMETALAREA                  4.144 LAYER ME2 ;
 ANTENNADIFFAREA                          5.472 LAYER ME2 ;
 ANTENNADIFFAREA                          5.472 LAYER ME3 ;
 ANTENNADIFFAREA                          5.472 LAYER ME4 ;
END DO74
PIN DI74
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 1574.400 0.000 1575.200 1.000 ;
  LAYER ME3 ;
  RECT 1574.400 0.000 1575.200 1.000 ;
  LAYER ME2 ;
  RECT 1574.400 0.000 1575.200 1.000 ;
  LAYER ME1 ;
  RECT 1574.400 0.000 1575.200 1.000 ;
 END
 ANTENNAPARTIALMETALAREA                  3.154 LAYER ME2 ;
 ANTENNAGATEAREA                          0.086 LAYER ME2 ;
 ANTENNAGATEAREA                          0.086 LAYER ME3 ;
 ANTENNAGATEAREA                          0.086 LAYER ME4 ;
 ANTENNADIFFAREA                          0.160 LAYER ME2 ;
 ANTENNADIFFAREA                          0.160 LAYER ME3 ;
 ANTENNADIFFAREA                          0.160 LAYER ME4 ;
 ANTENNAMAXAREACAR                       48.847 LAYER ME2 ;
 ANTENNAMAXAREACAR                       58.106 LAYER ME3 ;
 ANTENNAMAXAREACAR                       67.366 LAYER ME4 ;
END DI74
PIN DO73
  DIRECTION OUTPUT ;
 PORT
  LAYER ME4 ;
  RECT 1568.000 0.000 1568.800 1.000 ;
  LAYER ME3 ;
  RECT 1568.000 0.000 1568.800 1.000 ;
  LAYER ME2 ;
  RECT 1568.000 0.000 1568.800 1.000 ;
  LAYER ME1 ;
  RECT 1568.000 0.000 1568.800 1.000 ;
 END
 ANTENNAPARTIALMETALAREA                  4.168 LAYER ME2 ;
 ANTENNADIFFAREA                          5.472 LAYER ME2 ;
 ANTENNADIFFAREA                          5.472 LAYER ME3 ;
 ANTENNADIFFAREA                          5.472 LAYER ME4 ;
END DO73
PIN DI73
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 1553.600 0.000 1554.400 1.000 ;
  LAYER ME3 ;
  RECT 1553.600 0.000 1554.400 1.000 ;
  LAYER ME2 ;
  RECT 1553.600 0.000 1554.400 1.000 ;
  LAYER ME1 ;
  RECT 1553.600 0.000 1554.400 1.000 ;
 END
 ANTENNAPARTIALMETALAREA                  3.134 LAYER ME2 ;
 ANTENNAGATEAREA                          0.086 LAYER ME2 ;
 ANTENNAGATEAREA                          0.086 LAYER ME3 ;
 ANTENNAGATEAREA                          0.086 LAYER ME4 ;
 ANTENNADIFFAREA                          0.160 LAYER ME2 ;
 ANTENNADIFFAREA                          0.160 LAYER ME3 ;
 ANTENNADIFFAREA                          0.160 LAYER ME4 ;
 ANTENNAMAXAREACAR                       48.616 LAYER ME2 ;
 ANTENNAMAXAREACAR                       57.875 LAYER ME3 ;
 ANTENNAMAXAREACAR                       67.134 LAYER ME4 ;
END DI73
PIN DO72
  DIRECTION OUTPUT ;
 PORT
  LAYER ME4 ;
  RECT 1548.400 0.000 1549.200 1.000 ;
  LAYER ME3 ;
  RECT 1548.400 0.000 1549.200 1.000 ;
  LAYER ME2 ;
  RECT 1548.400 0.000 1549.200 1.000 ;
  LAYER ME1 ;
  RECT 1548.400 0.000 1549.200 1.000 ;
 END
 ANTENNAPARTIALMETALAREA                  4.160 LAYER ME2 ;
 ANTENNADIFFAREA                          5.472 LAYER ME2 ;
 ANTENNADIFFAREA                          5.472 LAYER ME3 ;
 ANTENNADIFFAREA                          5.472 LAYER ME4 ;
END DO72
PIN DI72
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 1533.600 0.000 1534.400 1.000 ;
  LAYER ME3 ;
  RECT 1533.600 0.000 1534.400 1.000 ;
  LAYER ME2 ;
  RECT 1533.600 0.000 1534.400 1.000 ;
  LAYER ME1 ;
  RECT 1533.600 0.000 1534.400 1.000 ;
 END
 ANTENNAPARTIALMETALAREA                  3.130 LAYER ME2 ;
 ANTENNAGATEAREA                          0.086 LAYER ME2 ;
 ANTENNAGATEAREA                          0.086 LAYER ME3 ;
 ANTENNAGATEAREA                          0.086 LAYER ME4 ;
 ANTENNADIFFAREA                          0.160 LAYER ME2 ;
 ANTENNADIFFAREA                          0.160 LAYER ME3 ;
 ANTENNADIFFAREA                          0.160 LAYER ME4 ;
 ANTENNAMAXAREACAR                       48.569 LAYER ME2 ;
 ANTENNAMAXAREACAR                       57.829 LAYER ME3 ;
 ANTENNAMAXAREACAR                       67.088 LAYER ME4 ;
END DI72
PIN DO71
  DIRECTION OUTPUT ;
 PORT
  LAYER ME4 ;
  RECT 1527.200 0.000 1528.000 1.000 ;
  LAYER ME3 ;
  RECT 1527.200 0.000 1528.000 1.000 ;
  LAYER ME2 ;
  RECT 1527.200 0.000 1528.000 1.000 ;
  LAYER ME1 ;
  RECT 1527.200 0.000 1528.000 1.000 ;
 END
 ANTENNAPARTIALMETALAREA                  4.144 LAYER ME2 ;
 ANTENNADIFFAREA                          5.472 LAYER ME2 ;
 ANTENNADIFFAREA                          5.472 LAYER ME3 ;
 ANTENNADIFFAREA                          5.472 LAYER ME4 ;
END DO71
PIN DI71
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 1512.400 0.000 1513.200 1.000 ;
  LAYER ME3 ;
  RECT 1512.400 0.000 1513.200 1.000 ;
  LAYER ME2 ;
  RECT 1512.400 0.000 1513.200 1.000 ;
  LAYER ME1 ;
  RECT 1512.400 0.000 1513.200 1.000 ;
 END
 ANTENNAPARTIALMETALAREA                  3.154 LAYER ME2 ;
 ANTENNAGATEAREA                          0.086 LAYER ME2 ;
 ANTENNAGATEAREA                          0.086 LAYER ME3 ;
 ANTENNAGATEAREA                          0.086 LAYER ME4 ;
 ANTENNADIFFAREA                          0.160 LAYER ME2 ;
 ANTENNADIFFAREA                          0.160 LAYER ME3 ;
 ANTENNADIFFAREA                          0.160 LAYER ME4 ;
 ANTENNAMAXAREACAR                       48.847 LAYER ME2 ;
 ANTENNAMAXAREACAR                       58.106 LAYER ME3 ;
 ANTENNAMAXAREACAR                       67.366 LAYER ME4 ;
END DI71
PIN DO70
  DIRECTION OUTPUT ;
 PORT
  LAYER ME4 ;
  RECT 1507.200 0.000 1508.000 1.000 ;
  LAYER ME3 ;
  RECT 1507.200 0.000 1508.000 1.000 ;
  LAYER ME2 ;
  RECT 1507.200 0.000 1508.000 1.000 ;
  LAYER ME1 ;
  RECT 1507.200 0.000 1508.000 1.000 ;
 END
 ANTENNAPARTIALMETALAREA                  4.176 LAYER ME2 ;
 ANTENNADIFFAREA                          5.472 LAYER ME2 ;
 ANTENNADIFFAREA                          5.472 LAYER ME3 ;
 ANTENNADIFFAREA                          5.472 LAYER ME4 ;
END DO70
PIN DI70
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 1492.800 0.000 1493.600 1.000 ;
  LAYER ME3 ;
  RECT 1492.800 0.000 1493.600 1.000 ;
  LAYER ME2 ;
  RECT 1492.800 0.000 1493.600 1.000 ;
  LAYER ME1 ;
  RECT 1492.800 0.000 1493.600 1.000 ;
 END
 ANTENNAPARTIALMETALAREA                  3.126 LAYER ME2 ;
 ANTENNAGATEAREA                          0.086 LAYER ME2 ;
 ANTENNAGATEAREA                          0.086 LAYER ME3 ;
 ANTENNAGATEAREA                          0.086 LAYER ME4 ;
 ANTENNADIFFAREA                          0.160 LAYER ME2 ;
 ANTENNADIFFAREA                          0.160 LAYER ME3 ;
 ANTENNADIFFAREA                          0.160 LAYER ME4 ;
 ANTENNAMAXAREACAR                       48.523 LAYER ME2 ;
 ANTENNAMAXAREACAR                       57.782 LAYER ME3 ;
 ANTENNAMAXAREACAR                       67.042 LAYER ME4 ;
END DI70
PIN DO69
  DIRECTION OUTPUT ;
 PORT
  LAYER ME4 ;
  RECT 1486.400 0.000 1487.200 1.000 ;
  LAYER ME3 ;
  RECT 1486.400 0.000 1487.200 1.000 ;
  LAYER ME2 ;
  RECT 1486.400 0.000 1487.200 1.000 ;
  LAYER ME1 ;
  RECT 1486.400 0.000 1487.200 1.000 ;
 END
 ANTENNAPARTIALMETALAREA                  4.160 LAYER ME2 ;
 ANTENNADIFFAREA                          5.472 LAYER ME2 ;
 ANTENNADIFFAREA                          5.472 LAYER ME3 ;
 ANTENNADIFFAREA                          5.472 LAYER ME4 ;
END DO69
PIN DI69
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 1471.600 0.000 1472.400 1.000 ;
  LAYER ME3 ;
  RECT 1471.600 0.000 1472.400 1.000 ;
  LAYER ME2 ;
  RECT 1471.600 0.000 1472.400 1.000 ;
  LAYER ME1 ;
  RECT 1471.600 0.000 1472.400 1.000 ;
 END
 ANTENNAPARTIALMETALAREA                  3.130 LAYER ME2 ;
 ANTENNAGATEAREA                          0.086 LAYER ME2 ;
 ANTENNAGATEAREA                          0.086 LAYER ME3 ;
 ANTENNAGATEAREA                          0.086 LAYER ME4 ;
 ANTENNADIFFAREA                          0.160 LAYER ME2 ;
 ANTENNADIFFAREA                          0.160 LAYER ME3 ;
 ANTENNADIFFAREA                          0.160 LAYER ME4 ;
 ANTENNAMAXAREACAR                       48.569 LAYER ME2 ;
 ANTENNAMAXAREACAR                       57.829 LAYER ME3 ;
 ANTENNAMAXAREACAR                       67.088 LAYER ME4 ;
END DI69
PIN DO68
  DIRECTION OUTPUT ;
 PORT
  LAYER ME4 ;
  RECT 1466.400 0.000 1467.200 1.000 ;
  LAYER ME3 ;
  RECT 1466.400 0.000 1467.200 1.000 ;
  LAYER ME2 ;
  RECT 1466.400 0.000 1467.200 1.000 ;
  LAYER ME1 ;
  RECT 1466.400 0.000 1467.200 1.000 ;
 END
 ANTENNAPARTIALMETALAREA                  4.152 LAYER ME2 ;
 ANTENNADIFFAREA                          5.472 LAYER ME2 ;
 ANTENNADIFFAREA                          5.472 LAYER ME3 ;
 ANTENNADIFFAREA                          5.472 LAYER ME4 ;
END DO68
PIN DI68
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 1452.000 0.000 1452.800 1.000 ;
  LAYER ME3 ;
  RECT 1452.000 0.000 1452.800 1.000 ;
  LAYER ME2 ;
  RECT 1452.000 0.000 1452.800 1.000 ;
  LAYER ME1 ;
  RECT 1452.000 0.000 1452.800 1.000 ;
 END
 ANTENNAPARTIALMETALAREA                  3.150 LAYER ME2 ;
 ANTENNAGATEAREA                          0.086 LAYER ME2 ;
 ANTENNAGATEAREA                          0.086 LAYER ME3 ;
 ANTENNAGATEAREA                          0.086 LAYER ME4 ;
 ANTENNADIFFAREA                          0.160 LAYER ME2 ;
 ANTENNADIFFAREA                          0.160 LAYER ME3 ;
 ANTENNADIFFAREA                          0.160 LAYER ME4 ;
 ANTENNAMAXAREACAR                       48.801 LAYER ME2 ;
 ANTENNAMAXAREACAR                       58.060 LAYER ME3 ;
 ANTENNAMAXAREACAR                       67.319 LAYER ME4 ;
END DI68
PIN DO67
  DIRECTION OUTPUT ;
 PORT
  LAYER ME4 ;
  RECT 1445.200 0.000 1446.000 1.000 ;
  LAYER ME3 ;
  RECT 1445.200 0.000 1446.000 1.000 ;
  LAYER ME2 ;
  RECT 1445.200 0.000 1446.000 1.000 ;
  LAYER ME1 ;
  RECT 1445.200 0.000 1446.000 1.000 ;
 END
 ANTENNAPARTIALMETALAREA                  4.176 LAYER ME2 ;
 ANTENNADIFFAREA                          5.472 LAYER ME2 ;
 ANTENNADIFFAREA                          5.472 LAYER ME3 ;
 ANTENNADIFFAREA                          5.472 LAYER ME4 ;
END DO67
PIN DI67
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 1430.800 0.000 1431.600 1.000 ;
  LAYER ME3 ;
  RECT 1430.800 0.000 1431.600 1.000 ;
  LAYER ME2 ;
  RECT 1430.800 0.000 1431.600 1.000 ;
  LAYER ME1 ;
  RECT 1430.800 0.000 1431.600 1.000 ;
 END
 ANTENNAPARTIALMETALAREA                  3.126 LAYER ME2 ;
 ANTENNAGATEAREA                          0.086 LAYER ME2 ;
 ANTENNAGATEAREA                          0.086 LAYER ME3 ;
 ANTENNAGATEAREA                          0.086 LAYER ME4 ;
 ANTENNADIFFAREA                          0.160 LAYER ME2 ;
 ANTENNADIFFAREA                          0.160 LAYER ME3 ;
 ANTENNADIFFAREA                          0.160 LAYER ME4 ;
 ANTENNAMAXAREACAR                       48.523 LAYER ME2 ;
 ANTENNAMAXAREACAR                       57.782 LAYER ME3 ;
 ANTENNAMAXAREACAR                       67.042 LAYER ME4 ;
END DI67
PIN DO66
  DIRECTION OUTPUT ;
 PORT
  LAYER ME4 ;
  RECT 1425.600 0.000 1426.400 1.000 ;
  LAYER ME3 ;
  RECT 1425.600 0.000 1426.400 1.000 ;
  LAYER ME2 ;
  RECT 1425.600 0.000 1426.400 1.000 ;
  LAYER ME1 ;
  RECT 1425.600 0.000 1426.400 1.000 ;
 END
 ANTENNAPARTIALMETALAREA                  4.152 LAYER ME2 ;
 ANTENNADIFFAREA                          5.472 LAYER ME2 ;
 ANTENNADIFFAREA                          5.472 LAYER ME3 ;
 ANTENNADIFFAREA                          5.472 LAYER ME4 ;
END DO66
PIN DI66
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 1410.800 0.000 1411.600 1.000 ;
  LAYER ME3 ;
  RECT 1410.800 0.000 1411.600 1.000 ;
  LAYER ME2 ;
  RECT 1410.800 0.000 1411.600 1.000 ;
  LAYER ME1 ;
  RECT 1410.800 0.000 1411.600 1.000 ;
 END
 ANTENNAPARTIALMETALAREA                  3.138 LAYER ME2 ;
 ANTENNAGATEAREA                          0.086 LAYER ME2 ;
 ANTENNAGATEAREA                          0.086 LAYER ME3 ;
 ANTENNAGATEAREA                          0.086 LAYER ME4 ;
 ANTENNADIFFAREA                          0.160 LAYER ME2 ;
 ANTENNADIFFAREA                          0.160 LAYER ME3 ;
 ANTENNADIFFAREA                          0.160 LAYER ME4 ;
 ANTENNAMAXAREACAR                       48.662 LAYER ME2 ;
 ANTENNAMAXAREACAR                       57.921 LAYER ME3 ;
 ANTENNAMAXAREACAR                       67.181 LAYER ME4 ;
END DI66
PIN DO65
  DIRECTION OUTPUT ;
 PORT
  LAYER ME4 ;
  RECT 1404.400 0.000 1405.200 1.000 ;
  LAYER ME3 ;
  RECT 1404.400 0.000 1405.200 1.000 ;
  LAYER ME2 ;
  RECT 1404.400 0.000 1405.200 1.000 ;
  LAYER ME1 ;
  RECT 1404.400 0.000 1405.200 1.000 ;
 END
 ANTENNAPARTIALMETALAREA                  4.152 LAYER ME2 ;
 ANTENNADIFFAREA                          5.472 LAYER ME2 ;
 ANTENNADIFFAREA                          5.472 LAYER ME3 ;
 ANTENNADIFFAREA                          5.472 LAYER ME4 ;
END DO65
PIN DI65
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 1390.000 0.000 1390.800 1.000 ;
  LAYER ME3 ;
  RECT 1390.000 0.000 1390.800 1.000 ;
  LAYER ME2 ;
  RECT 1390.000 0.000 1390.800 1.000 ;
  LAYER ME1 ;
  RECT 1390.000 0.000 1390.800 1.000 ;
 END
 ANTENNAPARTIALMETALAREA                  3.150 LAYER ME2 ;
 ANTENNAGATEAREA                          0.086 LAYER ME2 ;
 ANTENNAGATEAREA                          0.086 LAYER ME3 ;
 ANTENNAGATEAREA                          0.086 LAYER ME4 ;
 ANTENNADIFFAREA                          0.160 LAYER ME2 ;
 ANTENNADIFFAREA                          0.160 LAYER ME3 ;
 ANTENNADIFFAREA                          0.160 LAYER ME4 ;
 ANTENNAMAXAREACAR                       48.801 LAYER ME2 ;
 ANTENNAMAXAREACAR                       58.060 LAYER ME3 ;
 ANTENNAMAXAREACAR                       67.319 LAYER ME4 ;
END DI65
PIN DO64
  DIRECTION OUTPUT ;
 PORT
  LAYER ME4 ;
  RECT 1384.800 0.000 1385.600 1.000 ;
  LAYER ME3 ;
  RECT 1384.800 0.000 1385.600 1.000 ;
  LAYER ME2 ;
  RECT 1384.800 0.000 1385.600 1.000 ;
  LAYER ME1 ;
  RECT 1384.800 0.000 1385.600 1.000 ;
 END
 ANTENNAPARTIALMETALAREA                  4.176 LAYER ME2 ;
 ANTENNADIFFAREA                          5.472 LAYER ME2 ;
 ANTENNADIFFAREA                          5.472 LAYER ME3 ;
 ANTENNADIFFAREA                          5.472 LAYER ME4 ;
END DO64
PIN WEB4
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 1371.600 0.000 1372.400 1.000 ;
  LAYER ME3 ;
  RECT 1371.600 0.000 1372.400 1.000 ;
  LAYER ME2 ;
  RECT 1371.600 0.000 1372.400 1.000 ;
  LAYER ME1 ;
  RECT 1371.600 0.000 1372.400 1.000 ;
 END
 ANTENNAPARTIALMETALAREA                  2.852 LAYER ME2 ;
 ANTENNAGATEAREA                          0.072 LAYER ME2 ;
 ANTENNAGATEAREA                          0.072 LAYER ME3 ;
 ANTENNAGATEAREA                          0.072 LAYER ME4 ;
 ANTENNADIFFAREA                          0.160 LAYER ME2 ;
 ANTENNADIFFAREA                          0.160 LAYER ME3 ;
 ANTENNADIFFAREA                          0.160 LAYER ME4 ;
 ANTENNAMAXAREACAR                       54.622 LAYER ME2 ;
 ANTENNAMAXAREACAR                       65.733 LAYER ME3 ;
 ANTENNAMAXAREACAR                       76.844 LAYER ME4 ;
END WEB4
PIN DI64
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 1370.000 0.000 1370.800 1.000 ;
  LAYER ME3 ;
  RECT 1370.000 0.000 1370.800 1.000 ;
  LAYER ME2 ;
  RECT 1370.000 0.000 1370.800 1.000 ;
  LAYER ME1 ;
  RECT 1370.000 0.000 1370.800 1.000 ;
 END
 ANTENNAPARTIALMETALAREA                  3.118 LAYER ME2 ;
 ANTENNAGATEAREA                          0.086 LAYER ME2 ;
 ANTENNAGATEAREA                          0.086 LAYER ME3 ;
 ANTENNAGATEAREA                          0.086 LAYER ME4 ;
 ANTENNADIFFAREA                          0.160 LAYER ME2 ;
 ANTENNADIFFAREA                          0.160 LAYER ME3 ;
 ANTENNADIFFAREA                          0.160 LAYER ME4 ;
 ANTENNAMAXAREACAR                       48.431 LAYER ME2 ;
 ANTENNAMAXAREACAR                       57.690 LAYER ME3 ;
 ANTENNAMAXAREACAR                       66.949 LAYER ME4 ;
END DI64
PIN A3
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 1349.200 0.000 1350.000 1.000 ;
  LAYER ME3 ;
  RECT 1349.200 0.000 1350.000 1.000 ;
  LAYER ME2 ;
  RECT 1349.200 0.000 1350.000 1.000 ;
  LAYER ME1 ;
  RECT 1349.200 0.000 1350.000 1.000 ;
 END
 ANTENNAPARTIALMETALAREA                  2.028 LAYER ME2 ;
 ANTENNAGATEAREA                          0.180 LAYER ME2 ;
 ANTENNAGATEAREA                          0.180 LAYER ME3 ;
 ANTENNAGATEAREA                          0.180 LAYER ME4 ;
 ANTENNADIFFAREA                          0.160 LAYER ME2 ;
 ANTENNADIFFAREA                          0.160 LAYER ME3 ;
 ANTENNADIFFAREA                          0.160 LAYER ME4 ;
 ANTENNAMAXAREACAR                       17.116 LAYER ME2 ;
 ANTENNAMAXAREACAR                       21.560 LAYER ME3 ;
 ANTENNAMAXAREACAR                       26.004 LAYER ME4 ;
END A3
PIN A1
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 1348.000 0.000 1348.800 1.000 ;
  LAYER ME3 ;
  RECT 1348.000 0.000 1348.800 1.000 ;
  LAYER ME2 ;
  RECT 1348.000 0.000 1348.800 1.000 ;
  LAYER ME1 ;
  RECT 1348.000 0.000 1348.800 1.000 ;
 END
 ANTENNAPARTIALMETALAREA                  7.298 LAYER ME2 ;
 ANTENNAGATEAREA                          0.192 LAYER ME2 ;
 ANTENNAGATEAREA                          0.192 LAYER ME3 ;
 ANTENNAGATEAREA                          0.192 LAYER ME4 ;
 ANTENNADIFFAREA                          0.160 LAYER ME2 ;
 ANTENNADIFFAREA                          0.160 LAYER ME3 ;
 ANTENNADIFFAREA                          0.160 LAYER ME4 ;
 ANTENNAMAXAREACAR                       43.452 LAYER ME2 ;
 ANTENNAMAXAREACAR                       47.619 LAYER ME3 ;
 ANTENNAMAXAREACAR                       51.785 LAYER ME4 ;
END A1
PIN OE
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 1346.800 0.000 1347.600 1.000 ;
  LAYER ME3 ;
  RECT 1346.800 0.000 1347.600 1.000 ;
  LAYER ME2 ;
  RECT 1346.800 0.000 1347.600 1.000 ;
  LAYER ME1 ;
  RECT 1346.800 0.000 1347.600 1.000 ;
 END
 ANTENNAPARTIALMETALAREA                  3.370 LAYER ME2 ;
 ANTENNAGATEAREA                          0.840 LAYER ME2 ;
 ANTENNAGATEAREA                          0.840 LAYER ME3 ;
 ANTENNAGATEAREA                          0.840 LAYER ME4 ;
 ANTENNADIFFAREA                          0.160 LAYER ME2 ;
 ANTENNADIFFAREA                          0.160 LAYER ME3 ;
 ANTENNADIFFAREA                          0.160 LAYER ME4 ;
 ANTENNAMAXAREACAR                        5.336 LAYER ME2 ;
 ANTENNAMAXAREACAR                        6.288 LAYER ME3 ;
 ANTENNAMAXAREACAR                        7.240 LAYER ME4 ;
END OE
PIN CS
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 1345.600 0.000 1346.400 1.000 ;
  LAYER ME3 ;
  RECT 1345.600 0.000 1346.400 1.000 ;
  LAYER ME2 ;
  RECT 1345.600 0.000 1346.400 1.000 ;
  LAYER ME1 ;
  RECT 1345.600 0.000 1346.400 1.000 ;
 END
 ANTENNAPARTIALMETALAREA                  5.076 LAYER ME2 ;
 ANTENNAGATEAREA                          1.680 LAYER ME2 ;
 ANTENNAGATEAREA                          1.680 LAYER ME3 ;
 ANTENNAGATEAREA                          1.680 LAYER ME4 ;
 ANTENNADIFFAREA                          0.160 LAYER ME2 ;
 ANTENNADIFFAREA                          0.160 LAYER ME3 ;
 ANTENNADIFFAREA                          0.160 LAYER ME4 ;
 ANTENNAMAXAREACAR                        3.648 LAYER ME2 ;
 ANTENNAMAXAREACAR                        4.124 LAYER ME3 ;
 ANTENNAMAXAREACAR                        4.600 LAYER ME4 ;
END CS
PIN A2
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 1344.400 0.000 1345.200 1.000 ;
  LAYER ME3 ;
  RECT 1344.400 0.000 1345.200 1.000 ;
  LAYER ME2 ;
  RECT 1344.400 0.000 1345.200 1.000 ;
  LAYER ME1 ;
  RECT 1344.400 0.000 1345.200 1.000 ;
 END
 ANTENNAPARTIALMETALAREA                  7.366 LAYER ME2 ;
 ANTENNAGATEAREA                          0.192 LAYER ME2 ;
 ANTENNAGATEAREA                          0.192 LAYER ME3 ;
 ANTENNAGATEAREA                          0.192 LAYER ME4 ;
 ANTENNADIFFAREA                          0.160 LAYER ME2 ;
 ANTENNADIFFAREA                          0.160 LAYER ME3 ;
 ANTENNADIFFAREA                          0.160 LAYER ME4 ;
 ANTENNAMAXAREACAR                       43.806 LAYER ME2 ;
 ANTENNAMAXAREACAR                       47.973 LAYER ME3 ;
 ANTENNAMAXAREACAR                       52.140 LAYER ME4 ;
END A2
PIN A0
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 1343.200 0.000 1344.000 1.000 ;
  LAYER ME3 ;
  RECT 1343.200 0.000 1344.000 1.000 ;
  LAYER ME2 ;
  RECT 1343.200 0.000 1344.000 1.000 ;
  LAYER ME1 ;
  RECT 1343.200 0.000 1344.000 1.000 ;
 END
 ANTENNAPARTIALMETALAREA                  7.418 LAYER ME2 ;
 ANTENNAGATEAREA                          0.192 LAYER ME2 ;
 ANTENNAGATEAREA                          0.192 LAYER ME3 ;
 ANTENNAGATEAREA                          0.192 LAYER ME4 ;
 ANTENNADIFFAREA                          0.160 LAYER ME2 ;
 ANTENNADIFFAREA                          0.160 LAYER ME3 ;
 ANTENNADIFFAREA                          0.160 LAYER ME4 ;
 ANTENNAMAXAREACAR                       44.077 LAYER ME2 ;
 ANTENNAMAXAREACAR                       48.244 LAYER ME3 ;
 ANTENNAMAXAREACAR                       52.410 LAYER ME4 ;
END A0
PIN CK
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 1337.200 0.000 1338.000 1.000 ;
  LAYER ME3 ;
  RECT 1337.200 0.000 1338.000 1.000 ;
  LAYER ME2 ;
  RECT 1337.200 0.000 1338.000 1.000 ;
  LAYER ME1 ;
  RECT 1337.200 0.000 1338.000 1.000 ;
 END
 ANTENNAPARTIALMETALAREA                  5.506 LAYER ME2 ;
 ANTENNAGATEAREA                          1.908 LAYER ME2 ;
 ANTENNAGATEAREA                          1.908 LAYER ME3 ;
 ANTENNAGATEAREA                          1.908 LAYER ME4 ;
 ANTENNADIFFAREA                          0.160 LAYER ME2 ;
 ANTENNADIFFAREA                          0.160 LAYER ME3 ;
 ANTENNADIFFAREA                          0.160 LAYER ME4 ;
 ANTENNAMAXAREACAR                       59.337 LAYER ME2 ;
 ANTENNAMAXAREACAR                       66.744 LAYER ME3 ;
 ANTENNAMAXAREACAR                       74.152 LAYER ME4 ;
END CK
PIN A4
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 1330.000 0.000 1330.800 1.000 ;
  LAYER ME3 ;
  RECT 1330.000 0.000 1330.800 1.000 ;
  LAYER ME2 ;
  RECT 1330.000 0.000 1330.800 1.000 ;
  LAYER ME1 ;
  RECT 1330.000 0.000 1330.800 1.000 ;
 END
 ANTENNAPARTIALMETALAREA                  2.212 LAYER ME2 ;
 ANTENNAGATEAREA                          0.180 LAYER ME2 ;
 ANTENNAGATEAREA                          0.180 LAYER ME3 ;
 ANTENNAGATEAREA                          0.180 LAYER ME4 ;
 ANTENNADIFFAREA                          0.160 LAYER ME2 ;
 ANTENNADIFFAREA                          0.160 LAYER ME3 ;
 ANTENNADIFFAREA                          0.160 LAYER ME4 ;
 ANTENNAMAXAREACAR                       18.181 LAYER ME2 ;
 ANTENNAMAXAREACAR                       22.626 LAYER ME3 ;
 ANTENNAMAXAREACAR                       27.070 LAYER ME4 ;
END A4
PIN A5
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 1327.200 0.000 1328.000 1.000 ;
  LAYER ME3 ;
  RECT 1327.200 0.000 1328.000 1.000 ;
  LAYER ME2 ;
  RECT 1327.200 0.000 1328.000 1.000 ;
  LAYER ME1 ;
  RECT 1327.200 0.000 1328.000 1.000 ;
 END
 ANTENNAPARTIALMETALAREA                  2.406 LAYER ME2 ;
 ANTENNAGATEAREA                          0.180 LAYER ME2 ;
 ANTENNAGATEAREA                          0.180 LAYER ME3 ;
 ANTENNAGATEAREA                          0.180 LAYER ME4 ;
 ANTENNADIFFAREA                          0.160 LAYER ME2 ;
 ANTENNADIFFAREA                          0.160 LAYER ME3 ;
 ANTENNADIFFAREA                          0.160 LAYER ME4 ;
 ANTENNAMAXAREACAR                       19.319 LAYER ME2 ;
 ANTENNAMAXAREACAR                       23.763 LAYER ME3 ;
 ANTENNAMAXAREACAR                       28.208 LAYER ME4 ;
END A5
PIN A6
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 1324.400 0.000 1325.200 1.000 ;
  LAYER ME3 ;
  RECT 1324.400 0.000 1325.200 1.000 ;
  LAYER ME2 ;
  RECT 1324.400 0.000 1325.200 1.000 ;
  LAYER ME1 ;
  RECT 1324.400 0.000 1325.200 1.000 ;
 END
 ANTENNAPARTIALMETALAREA                  2.394 LAYER ME2 ;
 ANTENNAGATEAREA                          0.180 LAYER ME2 ;
 ANTENNAGATEAREA                          0.180 LAYER ME3 ;
 ANTENNAGATEAREA                          0.180 LAYER ME4 ;
 ANTENNADIFFAREA                          0.160 LAYER ME2 ;
 ANTENNADIFFAREA                          0.160 LAYER ME3 ;
 ANTENNADIFFAREA                          0.160 LAYER ME4 ;
 ANTENNAMAXAREACAR                       19.156 LAYER ME2 ;
 ANTENNAMAXAREACAR                       23.600 LAYER ME3 ;
 ANTENNAMAXAREACAR                       28.044 LAYER ME4 ;
END A6
PIN A7
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 1322.000 0.000 1322.800 1.000 ;
  LAYER ME3 ;
  RECT 1322.000 0.000 1322.800 1.000 ;
  LAYER ME2 ;
  RECT 1322.000 0.000 1322.800 1.000 ;
  LAYER ME1 ;
  RECT 1322.000 0.000 1322.800 1.000 ;
 END
 ANTENNAPARTIALMETALAREA                  2.378 LAYER ME2 ;
 ANTENNAGATEAREA                          0.180 LAYER ME2 ;
 ANTENNAGATEAREA                          0.180 LAYER ME3 ;
 ANTENNAGATEAREA                          0.180 LAYER ME4 ;
 ANTENNADIFFAREA                          0.160 LAYER ME2 ;
 ANTENNADIFFAREA                          0.160 LAYER ME3 ;
 ANTENNADIFFAREA                          0.160 LAYER ME4 ;
 ANTENNAMAXAREACAR                       19.067 LAYER ME2 ;
 ANTENNAMAXAREACAR                       23.511 LAYER ME3 ;
 ANTENNAMAXAREACAR                       27.956 LAYER ME4 ;
END A7
PIN A8
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 1320.400 0.000 1321.200 1.000 ;
  LAYER ME3 ;
  RECT 1320.400 0.000 1321.200 1.000 ;
  LAYER ME2 ;
  RECT 1320.400 0.000 1321.200 1.000 ;
  LAYER ME1 ;
  RECT 1320.400 0.000 1321.200 1.000 ;
 END
 ANTENNAPARTIALMETALAREA                  2.394 LAYER ME2 ;
 ANTENNAGATEAREA                          0.180 LAYER ME2 ;
 ANTENNAGATEAREA                          0.180 LAYER ME3 ;
 ANTENNAGATEAREA                          0.180 LAYER ME4 ;
 ANTENNADIFFAREA                          0.160 LAYER ME2 ;
 ANTENNADIFFAREA                          0.160 LAYER ME3 ;
 ANTENNADIFFAREA                          0.160 LAYER ME4 ;
 ANTENNAMAXAREACAR                       19.156 LAYER ME2 ;
 ANTENNAMAXAREACAR                       23.600 LAYER ME3 ;
 ANTENNAMAXAREACAR                       28.044 LAYER ME4 ;
END A8
PIN A9
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 1318.000 0.000 1318.800 1.000 ;
  LAYER ME3 ;
  RECT 1318.000 0.000 1318.800 1.000 ;
  LAYER ME2 ;
  RECT 1318.000 0.000 1318.800 1.000 ;
  LAYER ME1 ;
  RECT 1318.000 0.000 1318.800 1.000 ;
 END
 ANTENNAPARTIALMETALAREA                  2.378 LAYER ME2 ;
 ANTENNAGATEAREA                          0.180 LAYER ME2 ;
 ANTENNAGATEAREA                          0.180 LAYER ME3 ;
 ANTENNAGATEAREA                          0.180 LAYER ME4 ;
 ANTENNADIFFAREA                          0.160 LAYER ME2 ;
 ANTENNADIFFAREA                          0.160 LAYER ME3 ;
 ANTENNADIFFAREA                          0.160 LAYER ME4 ;
 ANTENNAMAXAREACAR                       19.067 LAYER ME2 ;
 ANTENNAMAXAREACAR                       23.511 LAYER ME3 ;
 ANTENNAMAXAREACAR                       27.956 LAYER ME4 ;
END A9
PIN DO63
  DIRECTION OUTPUT ;
 PORT
  LAYER ME4 ;
  RECT 1311.200 0.000 1312.000 1.000 ;
  LAYER ME3 ;
  RECT 1311.200 0.000 1312.000 1.000 ;
  LAYER ME2 ;
  RECT 1311.200 0.000 1312.000 1.000 ;
  LAYER ME1 ;
  RECT 1311.200 0.000 1312.000 1.000 ;
 END
 ANTENNAPARTIALMETALAREA                  4.148 LAYER ME2 ;
 ANTENNADIFFAREA                          5.472 LAYER ME2 ;
 ANTENNADIFFAREA                          5.472 LAYER ME3 ;
 ANTENNADIFFAREA                          5.472 LAYER ME4 ;
END DO63
PIN DI63
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 1296.400 0.000 1297.200 1.000 ;
  LAYER ME3 ;
  RECT 1296.400 0.000 1297.200 1.000 ;
  LAYER ME2 ;
  RECT 1296.400 0.000 1297.200 1.000 ;
  LAYER ME1 ;
  RECT 1296.400 0.000 1297.200 1.000 ;
 END
 ANTENNAPARTIALMETALAREA                  3.142 LAYER ME2 ;
 ANTENNAGATEAREA                          0.086 LAYER ME2 ;
 ANTENNAGATEAREA                          0.086 LAYER ME3 ;
 ANTENNAGATEAREA                          0.086 LAYER ME4 ;
 ANTENNADIFFAREA                          0.160 LAYER ME2 ;
 ANTENNADIFFAREA                          0.160 LAYER ME3 ;
 ANTENNADIFFAREA                          0.160 LAYER ME4 ;
 ANTENNAMAXAREACAR                       48.708 LAYER ME2 ;
 ANTENNAMAXAREACAR                       57.968 LAYER ME3 ;
 ANTENNAMAXAREACAR                       67.227 LAYER ME4 ;
END DI63
PIN DO62
  DIRECTION OUTPUT ;
 PORT
  LAYER ME4 ;
  RECT 1291.200 0.000 1292.000 1.000 ;
  LAYER ME3 ;
  RECT 1291.200 0.000 1292.000 1.000 ;
  LAYER ME2 ;
  RECT 1291.200 0.000 1292.000 1.000 ;
  LAYER ME1 ;
  RECT 1291.200 0.000 1292.000 1.000 ;
 END
 ANTENNAPARTIALMETALAREA                  4.164 LAYER ME2 ;
 ANTENNADIFFAREA                          5.472 LAYER ME2 ;
 ANTENNADIFFAREA                          5.472 LAYER ME3 ;
 ANTENNADIFFAREA                          5.472 LAYER ME4 ;
END DO62
PIN DI62
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 1276.800 0.000 1277.600 1.000 ;
  LAYER ME3 ;
  RECT 1276.800 0.000 1277.600 1.000 ;
  LAYER ME2 ;
  RECT 1276.800 0.000 1277.600 1.000 ;
  LAYER ME1 ;
  RECT 1276.800 0.000 1277.600 1.000 ;
 END
 ANTENNAPARTIALMETALAREA                  3.138 LAYER ME2 ;
 ANTENNAGATEAREA                          0.086 LAYER ME2 ;
 ANTENNAGATEAREA                          0.086 LAYER ME3 ;
 ANTENNAGATEAREA                          0.086 LAYER ME4 ;
 ANTENNADIFFAREA                          0.160 LAYER ME2 ;
 ANTENNADIFFAREA                          0.160 LAYER ME3 ;
 ANTENNADIFFAREA                          0.160 LAYER ME4 ;
 ANTENNAMAXAREACAR                       48.662 LAYER ME2 ;
 ANTENNAMAXAREACAR                       57.921 LAYER ME3 ;
 ANTENNAMAXAREACAR                       67.181 LAYER ME4 ;
END DI62
PIN DO61
  DIRECTION OUTPUT ;
 PORT
  LAYER ME4 ;
  RECT 1270.400 0.000 1271.200 1.000 ;
  LAYER ME3 ;
  RECT 1270.400 0.000 1271.200 1.000 ;
  LAYER ME2 ;
  RECT 1270.400 0.000 1271.200 1.000 ;
  LAYER ME1 ;
  RECT 1270.400 0.000 1271.200 1.000 ;
 END
 ANTENNAPARTIALMETALAREA                  4.172 LAYER ME2 ;
 ANTENNADIFFAREA                          5.472 LAYER ME2 ;
 ANTENNADIFFAREA                          5.472 LAYER ME3 ;
 ANTENNADIFFAREA                          5.472 LAYER ME4 ;
END DO61
PIN DI61
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 1255.600 0.000 1256.400 1.000 ;
  LAYER ME3 ;
  RECT 1255.600 0.000 1256.400 1.000 ;
  LAYER ME2 ;
  RECT 1255.600 0.000 1256.400 1.000 ;
  LAYER ME1 ;
  RECT 1255.600 0.000 1256.400 1.000 ;
 END
 ANTENNAPARTIALMETALAREA                  3.118 LAYER ME2 ;
 ANTENNAGATEAREA                          0.086 LAYER ME2 ;
 ANTENNAGATEAREA                          0.086 LAYER ME3 ;
 ANTENNAGATEAREA                          0.086 LAYER ME4 ;
 ANTENNADIFFAREA                          0.160 LAYER ME2 ;
 ANTENNADIFFAREA                          0.160 LAYER ME3 ;
 ANTENNADIFFAREA                          0.160 LAYER ME4 ;
 ANTENNAMAXAREACAR                       48.431 LAYER ME2 ;
 ANTENNAMAXAREACAR                       57.690 LAYER ME3 ;
 ANTENNAMAXAREACAR                       66.949 LAYER ME4 ;
END DI61
PIN DO60
  DIRECTION OUTPUT ;
 PORT
  LAYER ME4 ;
  RECT 1250.400 0.000 1251.200 1.000 ;
  LAYER ME3 ;
  RECT 1250.400 0.000 1251.200 1.000 ;
  LAYER ME2 ;
  RECT 1250.400 0.000 1251.200 1.000 ;
  LAYER ME1 ;
  RECT 1250.400 0.000 1251.200 1.000 ;
 END
 ANTENNAPARTIALMETALAREA                  4.140 LAYER ME2 ;
 ANTENNADIFFAREA                          5.472 LAYER ME2 ;
 ANTENNADIFFAREA                          5.472 LAYER ME3 ;
 ANTENNADIFFAREA                          5.472 LAYER ME4 ;
END DO60
PIN DI60
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 1235.600 0.000 1236.400 1.000 ;
  LAYER ME3 ;
  RECT 1235.600 0.000 1236.400 1.000 ;
  LAYER ME2 ;
  RECT 1235.600 0.000 1236.400 1.000 ;
  LAYER ME1 ;
  RECT 1235.600 0.000 1236.400 1.000 ;
 END
 ANTENNAPARTIALMETALAREA                  3.150 LAYER ME2 ;
 ANTENNAGATEAREA                          0.086 LAYER ME2 ;
 ANTENNAGATEAREA                          0.086 LAYER ME3 ;
 ANTENNAGATEAREA                          0.086 LAYER ME4 ;
 ANTENNADIFFAREA                          0.160 LAYER ME2 ;
 ANTENNADIFFAREA                          0.160 LAYER ME3 ;
 ANTENNADIFFAREA                          0.160 LAYER ME4 ;
 ANTENNAMAXAREACAR                       48.801 LAYER ME2 ;
 ANTENNAMAXAREACAR                       58.060 LAYER ME3 ;
 ANTENNAMAXAREACAR                       67.319 LAYER ME4 ;
END DI60
PIN DO59
  DIRECTION OUTPUT ;
 PORT
  LAYER ME4 ;
  RECT 1229.200 0.000 1230.000 1.000 ;
  LAYER ME3 ;
  RECT 1229.200 0.000 1230.000 1.000 ;
  LAYER ME2 ;
  RECT 1229.200 0.000 1230.000 1.000 ;
  LAYER ME1 ;
  RECT 1229.200 0.000 1230.000 1.000 ;
 END
 ANTENNAPARTIALMETALAREA                  4.164 LAYER ME2 ;
 ANTENNADIFFAREA                          5.472 LAYER ME2 ;
 ANTENNADIFFAREA                          5.472 LAYER ME3 ;
 ANTENNADIFFAREA                          5.472 LAYER ME4 ;
END DO59
PIN DI59
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 1214.800 0.000 1215.600 1.000 ;
  LAYER ME3 ;
  RECT 1214.800 0.000 1215.600 1.000 ;
  LAYER ME2 ;
  RECT 1214.800 0.000 1215.600 1.000 ;
  LAYER ME1 ;
  RECT 1214.800 0.000 1215.600 1.000 ;
 END
 ANTENNAPARTIALMETALAREA                  3.138 LAYER ME2 ;
 ANTENNAGATEAREA                          0.086 LAYER ME2 ;
 ANTENNAGATEAREA                          0.086 LAYER ME3 ;
 ANTENNAGATEAREA                          0.086 LAYER ME4 ;
 ANTENNADIFFAREA                          0.160 LAYER ME2 ;
 ANTENNADIFFAREA                          0.160 LAYER ME3 ;
 ANTENNADIFFAREA                          0.160 LAYER ME4 ;
 ANTENNAMAXAREACAR                       48.662 LAYER ME2 ;
 ANTENNAMAXAREACAR                       57.921 LAYER ME3 ;
 ANTENNAMAXAREACAR                       67.181 LAYER ME4 ;
END DI59
PIN DO58
  DIRECTION OUTPUT ;
 PORT
  LAYER ME4 ;
  RECT 1209.600 0.000 1210.400 1.000 ;
  LAYER ME3 ;
  RECT 1209.600 0.000 1210.400 1.000 ;
  LAYER ME2 ;
  RECT 1209.600 0.000 1210.400 1.000 ;
  LAYER ME1 ;
  RECT 1209.600 0.000 1210.400 1.000 ;
 END
 ANTENNAPARTIALMETALAREA                  4.164 LAYER ME2 ;
 ANTENNADIFFAREA                          5.472 LAYER ME2 ;
 ANTENNADIFFAREA                          5.472 LAYER ME3 ;
 ANTENNADIFFAREA                          5.472 LAYER ME4 ;
END DO58
PIN DI58
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 1194.800 0.000 1195.600 1.000 ;
  LAYER ME3 ;
  RECT 1194.800 0.000 1195.600 1.000 ;
  LAYER ME2 ;
  RECT 1194.800 0.000 1195.600 1.000 ;
  LAYER ME1 ;
  RECT 1194.800 0.000 1195.600 1.000 ;
 END
 ANTENNAPARTIALMETALAREA                  3.126 LAYER ME2 ;
 ANTENNAGATEAREA                          0.086 LAYER ME2 ;
 ANTENNAGATEAREA                          0.086 LAYER ME3 ;
 ANTENNAGATEAREA                          0.086 LAYER ME4 ;
 ANTENNADIFFAREA                          0.160 LAYER ME2 ;
 ANTENNADIFFAREA                          0.160 LAYER ME3 ;
 ANTENNADIFFAREA                          0.160 LAYER ME4 ;
 ANTENNAMAXAREACAR                       48.523 LAYER ME2 ;
 ANTENNAMAXAREACAR                       57.782 LAYER ME3 ;
 ANTENNAMAXAREACAR                       67.042 LAYER ME4 ;
END DI58
PIN DO57
  DIRECTION OUTPUT ;
 PORT
  LAYER ME4 ;
  RECT 1188.400 0.000 1189.200 1.000 ;
  LAYER ME3 ;
  RECT 1188.400 0.000 1189.200 1.000 ;
  LAYER ME2 ;
  RECT 1188.400 0.000 1189.200 1.000 ;
  LAYER ME1 ;
  RECT 1188.400 0.000 1189.200 1.000 ;
 END
 ANTENNAPARTIALMETALAREA                  4.140 LAYER ME2 ;
 ANTENNADIFFAREA                          5.472 LAYER ME2 ;
 ANTENNADIFFAREA                          5.472 LAYER ME3 ;
 ANTENNADIFFAREA                          5.472 LAYER ME4 ;
END DO57
PIN DI57
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 1173.600 0.000 1174.400 1.000 ;
  LAYER ME3 ;
  RECT 1173.600 0.000 1174.400 1.000 ;
  LAYER ME2 ;
  RECT 1173.600 0.000 1174.400 1.000 ;
  LAYER ME1 ;
  RECT 1173.600 0.000 1174.400 1.000 ;
 END
 ANTENNAPARTIALMETALAREA                  3.150 LAYER ME2 ;
 ANTENNAGATEAREA                          0.086 LAYER ME2 ;
 ANTENNAGATEAREA                          0.086 LAYER ME3 ;
 ANTENNAGATEAREA                          0.086 LAYER ME4 ;
 ANTENNADIFFAREA                          0.160 LAYER ME2 ;
 ANTENNADIFFAREA                          0.160 LAYER ME3 ;
 ANTENNADIFFAREA                          0.160 LAYER ME4 ;
 ANTENNAMAXAREACAR                       48.801 LAYER ME2 ;
 ANTENNAMAXAREACAR                       58.060 LAYER ME3 ;
 ANTENNAMAXAREACAR                       67.319 LAYER ME4 ;
END DI57
PIN DO56
  DIRECTION OUTPUT ;
 PORT
  LAYER ME4 ;
  RECT 1168.400 0.000 1169.200 1.000 ;
  LAYER ME3 ;
  RECT 1168.400 0.000 1169.200 1.000 ;
  LAYER ME2 ;
  RECT 1168.400 0.000 1169.200 1.000 ;
  LAYER ME1 ;
  RECT 1168.400 0.000 1169.200 1.000 ;
 END
 ANTENNAPARTIALMETALAREA                  4.172 LAYER ME2 ;
 ANTENNADIFFAREA                          5.472 LAYER ME2 ;
 ANTENNADIFFAREA                          5.472 LAYER ME3 ;
 ANTENNADIFFAREA                          5.472 LAYER ME4 ;
END DO56
PIN DI56
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 1154.000 0.000 1154.800 1.000 ;
  LAYER ME3 ;
  RECT 1154.000 0.000 1154.800 1.000 ;
  LAYER ME2 ;
  RECT 1154.000 0.000 1154.800 1.000 ;
  LAYER ME1 ;
  RECT 1154.000 0.000 1154.800 1.000 ;
 END
 ANTENNAPARTIALMETALAREA                  3.130 LAYER ME2 ;
 ANTENNAGATEAREA                          0.086 LAYER ME2 ;
 ANTENNAGATEAREA                          0.086 LAYER ME3 ;
 ANTENNAGATEAREA                          0.086 LAYER ME4 ;
 ANTENNADIFFAREA                          0.160 LAYER ME2 ;
 ANTENNADIFFAREA                          0.160 LAYER ME3 ;
 ANTENNADIFFAREA                          0.160 LAYER ME4 ;
 ANTENNAMAXAREACAR                       48.569 LAYER ME2 ;
 ANTENNAMAXAREACAR                       57.829 LAYER ME3 ;
 ANTENNAMAXAREACAR                       67.088 LAYER ME4 ;
END DI56
PIN DO55
  DIRECTION OUTPUT ;
 PORT
  LAYER ME4 ;
  RECT 1147.600 0.000 1148.400 1.000 ;
  LAYER ME3 ;
  RECT 1147.600 0.000 1148.400 1.000 ;
  LAYER ME2 ;
  RECT 1147.600 0.000 1148.400 1.000 ;
  LAYER ME1 ;
  RECT 1147.600 0.000 1148.400 1.000 ;
 END
 ANTENNAPARTIALMETALAREA                  4.164 LAYER ME2 ;
 ANTENNADIFFAREA                          5.472 LAYER ME2 ;
 ANTENNADIFFAREA                          5.472 LAYER ME3 ;
 ANTENNADIFFAREA                          5.472 LAYER ME4 ;
END DO55
PIN DI55
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 1132.800 0.000 1133.600 1.000 ;
  LAYER ME3 ;
  RECT 1132.800 0.000 1133.600 1.000 ;
  LAYER ME2 ;
  RECT 1132.800 0.000 1133.600 1.000 ;
  LAYER ME1 ;
  RECT 1132.800 0.000 1133.600 1.000 ;
 END
 ANTENNAPARTIALMETALAREA                  3.126 LAYER ME2 ;
 ANTENNAGATEAREA                          0.086 LAYER ME2 ;
 ANTENNAGATEAREA                          0.086 LAYER ME3 ;
 ANTENNAGATEAREA                          0.086 LAYER ME4 ;
 ANTENNADIFFAREA                          0.160 LAYER ME2 ;
 ANTENNADIFFAREA                          0.160 LAYER ME3 ;
 ANTENNADIFFAREA                          0.160 LAYER ME4 ;
 ANTENNAMAXAREACAR                       48.523 LAYER ME2 ;
 ANTENNAMAXAREACAR                       57.782 LAYER ME3 ;
 ANTENNAMAXAREACAR                       67.042 LAYER ME4 ;
END DI55
PIN DO54
  DIRECTION OUTPUT ;
 PORT
  LAYER ME4 ;
  RECT 1127.600 0.000 1128.400 1.000 ;
  LAYER ME3 ;
  RECT 1127.600 0.000 1128.400 1.000 ;
  LAYER ME2 ;
  RECT 1127.600 0.000 1128.400 1.000 ;
  LAYER ME1 ;
  RECT 1127.600 0.000 1128.400 1.000 ;
 END
 ANTENNAPARTIALMETALAREA                  4.148 LAYER ME2 ;
 ANTENNADIFFAREA                          5.472 LAYER ME2 ;
 ANTENNADIFFAREA                          5.472 LAYER ME3 ;
 ANTENNADIFFAREA                          5.472 LAYER ME4 ;
END DO54
PIN DI54
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 1113.200 0.000 1114.000 1.000 ;
  LAYER ME3 ;
  RECT 1113.200 0.000 1114.000 1.000 ;
  LAYER ME2 ;
  RECT 1113.200 0.000 1114.000 1.000 ;
  LAYER ME1 ;
  RECT 1113.200 0.000 1114.000 1.000 ;
 END
 ANTENNAPARTIALMETALAREA                  3.154 LAYER ME2 ;
 ANTENNAGATEAREA                          0.086 LAYER ME2 ;
 ANTENNAGATEAREA                          0.086 LAYER ME3 ;
 ANTENNAGATEAREA                          0.086 LAYER ME4 ;
 ANTENNADIFFAREA                          0.160 LAYER ME2 ;
 ANTENNADIFFAREA                          0.160 LAYER ME3 ;
 ANTENNADIFFAREA                          0.160 LAYER ME4 ;
 ANTENNAMAXAREACAR                       48.847 LAYER ME2 ;
 ANTENNAMAXAREACAR                       58.106 LAYER ME3 ;
 ANTENNAMAXAREACAR                       67.366 LAYER ME4 ;
END DI54
PIN DO53
  DIRECTION OUTPUT ;
 PORT
  LAYER ME4 ;
  RECT 1106.400 0.000 1107.200 1.000 ;
  LAYER ME3 ;
  RECT 1106.400 0.000 1107.200 1.000 ;
  LAYER ME2 ;
  RECT 1106.400 0.000 1107.200 1.000 ;
  LAYER ME1 ;
  RECT 1106.400 0.000 1107.200 1.000 ;
 END
 ANTENNAPARTIALMETALAREA                  4.172 LAYER ME2 ;
 ANTENNADIFFAREA                          5.472 LAYER ME2 ;
 ANTENNADIFFAREA                          5.472 LAYER ME3 ;
 ANTENNADIFFAREA                          5.472 LAYER ME4 ;
END DO53
PIN DI53
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 1092.000 0.000 1092.800 1.000 ;
  LAYER ME3 ;
  RECT 1092.000 0.000 1092.800 1.000 ;
  LAYER ME2 ;
  RECT 1092.000 0.000 1092.800 1.000 ;
  LAYER ME1 ;
  RECT 1092.000 0.000 1092.800 1.000 ;
 END
 ANTENNAPARTIALMETALAREA                  3.130 LAYER ME2 ;
 ANTENNAGATEAREA                          0.086 LAYER ME2 ;
 ANTENNAGATEAREA                          0.086 LAYER ME3 ;
 ANTENNAGATEAREA                          0.086 LAYER ME4 ;
 ANTENNADIFFAREA                          0.160 LAYER ME2 ;
 ANTENNADIFFAREA                          0.160 LAYER ME3 ;
 ANTENNADIFFAREA                          0.160 LAYER ME4 ;
 ANTENNAMAXAREACAR                       48.569 LAYER ME2 ;
 ANTENNAMAXAREACAR                       57.829 LAYER ME3 ;
 ANTENNAMAXAREACAR                       67.088 LAYER ME4 ;
END DI53
PIN DO52
  DIRECTION OUTPUT ;
 PORT
  LAYER ME4 ;
  RECT 1086.800 0.000 1087.600 1.000 ;
  LAYER ME3 ;
  RECT 1086.800 0.000 1087.600 1.000 ;
  LAYER ME2 ;
  RECT 1086.800 0.000 1087.600 1.000 ;
  LAYER ME1 ;
  RECT 1086.800 0.000 1087.600 1.000 ;
 END
 ANTENNAPARTIALMETALAREA                  4.156 LAYER ME2 ;
 ANTENNADIFFAREA                          5.472 LAYER ME2 ;
 ANTENNADIFFAREA                          5.472 LAYER ME3 ;
 ANTENNADIFFAREA                          5.472 LAYER ME4 ;
END DO52
PIN DI52
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 1072.000 0.000 1072.800 1.000 ;
  LAYER ME3 ;
  RECT 1072.000 0.000 1072.800 1.000 ;
  LAYER ME2 ;
  RECT 1072.000 0.000 1072.800 1.000 ;
  LAYER ME1 ;
  RECT 1072.000 0.000 1072.800 1.000 ;
 END
 ANTENNAPARTIALMETALAREA                  3.134 LAYER ME2 ;
 ANTENNAGATEAREA                          0.086 LAYER ME2 ;
 ANTENNAGATEAREA                          0.086 LAYER ME3 ;
 ANTENNAGATEAREA                          0.086 LAYER ME4 ;
 ANTENNADIFFAREA                          0.160 LAYER ME2 ;
 ANTENNADIFFAREA                          0.160 LAYER ME3 ;
 ANTENNADIFFAREA                          0.160 LAYER ME4 ;
 ANTENNAMAXAREACAR                       48.616 LAYER ME2 ;
 ANTENNAMAXAREACAR                       57.875 LAYER ME3 ;
 ANTENNAMAXAREACAR                       67.134 LAYER ME4 ;
END DI52
PIN DO51
  DIRECTION OUTPUT ;
 PORT
  LAYER ME4 ;
  RECT 1065.600 0.000 1066.400 1.000 ;
  LAYER ME3 ;
  RECT 1065.600 0.000 1066.400 1.000 ;
  LAYER ME2 ;
  RECT 1065.600 0.000 1066.400 1.000 ;
  LAYER ME1 ;
  RECT 1065.600 0.000 1066.400 1.000 ;
 END
 ANTENNAPARTIALMETALAREA                  4.148 LAYER ME2 ;
 ANTENNADIFFAREA                          5.472 LAYER ME2 ;
 ANTENNADIFFAREA                          5.472 LAYER ME3 ;
 ANTENNADIFFAREA                          5.472 LAYER ME4 ;
END DO51
PIN DI51
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 1051.200 0.000 1052.000 1.000 ;
  LAYER ME3 ;
  RECT 1051.200 0.000 1052.000 1.000 ;
  LAYER ME2 ;
  RECT 1051.200 0.000 1052.000 1.000 ;
  LAYER ME1 ;
  RECT 1051.200 0.000 1052.000 1.000 ;
 END
 ANTENNAPARTIALMETALAREA                  3.154 LAYER ME2 ;
 ANTENNAGATEAREA                          0.086 LAYER ME2 ;
 ANTENNAGATEAREA                          0.086 LAYER ME3 ;
 ANTENNAGATEAREA                          0.086 LAYER ME4 ;
 ANTENNADIFFAREA                          0.160 LAYER ME2 ;
 ANTENNADIFFAREA                          0.160 LAYER ME3 ;
 ANTENNADIFFAREA                          0.160 LAYER ME4 ;
 ANTENNAMAXAREACAR                       48.847 LAYER ME2 ;
 ANTENNAMAXAREACAR                       58.106 LAYER ME3 ;
 ANTENNAMAXAREACAR                       67.366 LAYER ME4 ;
END DI51
PIN DO50
  DIRECTION OUTPUT ;
 PORT
  LAYER ME4 ;
  RECT 1045.600 0.000 1046.400 1.000 ;
  LAYER ME3 ;
  RECT 1045.600 0.000 1046.400 1.000 ;
  LAYER ME2 ;
  RECT 1045.600 0.000 1046.400 1.000 ;
  LAYER ME1 ;
  RECT 1045.600 0.000 1046.400 1.000 ;
 END
 ANTENNAPARTIALMETALAREA                  4.180 LAYER ME2 ;
 ANTENNADIFFAREA                          5.472 LAYER ME2 ;
 ANTENNADIFFAREA                          5.472 LAYER ME3 ;
 ANTENNADIFFAREA                          5.472 LAYER ME4 ;
END DO50
PIN DI50
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 1031.200 0.000 1032.000 1.000 ;
  LAYER ME3 ;
  RECT 1031.200 0.000 1032.000 1.000 ;
  LAYER ME2 ;
  RECT 1031.200 0.000 1032.000 1.000 ;
  LAYER ME1 ;
  RECT 1031.200 0.000 1032.000 1.000 ;
 END
 ANTENNAPARTIALMETALAREA                  3.122 LAYER ME2 ;
 ANTENNAGATEAREA                          0.086 LAYER ME2 ;
 ANTENNAGATEAREA                          0.086 LAYER ME3 ;
 ANTENNAGATEAREA                          0.086 LAYER ME4 ;
 ANTENNADIFFAREA                          0.160 LAYER ME2 ;
 ANTENNADIFFAREA                          0.160 LAYER ME3 ;
 ANTENNADIFFAREA                          0.160 LAYER ME4 ;
 ANTENNAMAXAREACAR                       48.477 LAYER ME2 ;
 ANTENNAMAXAREACAR                       57.736 LAYER ME3 ;
 ANTENNAMAXAREACAR                       66.995 LAYER ME4 ;
END DI50
PIN DO49
  DIRECTION OUTPUT ;
 PORT
  LAYER ME4 ;
  RECT 1024.800 0.000 1025.600 1.000 ;
  LAYER ME3 ;
  RECT 1024.800 0.000 1025.600 1.000 ;
  LAYER ME2 ;
  RECT 1024.800 0.000 1025.600 1.000 ;
  LAYER ME1 ;
  RECT 1024.800 0.000 1025.600 1.000 ;
 END
 ANTENNAPARTIALMETALAREA                  4.156 LAYER ME2 ;
 ANTENNADIFFAREA                          5.472 LAYER ME2 ;
 ANTENNADIFFAREA                          5.472 LAYER ME3 ;
 ANTENNADIFFAREA                          5.472 LAYER ME4 ;
END DO49
PIN DI49
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 1010.000 0.000 1010.800 1.000 ;
  LAYER ME3 ;
  RECT 1010.000 0.000 1010.800 1.000 ;
  LAYER ME2 ;
  RECT 1010.000 0.000 1010.800 1.000 ;
  LAYER ME1 ;
  RECT 1010.000 0.000 1010.800 1.000 ;
 END
 ANTENNAPARTIALMETALAREA                  3.134 LAYER ME2 ;
 ANTENNAGATEAREA                          0.086 LAYER ME2 ;
 ANTENNAGATEAREA                          0.086 LAYER ME3 ;
 ANTENNAGATEAREA                          0.086 LAYER ME4 ;
 ANTENNADIFFAREA                          0.160 LAYER ME2 ;
 ANTENNADIFFAREA                          0.160 LAYER ME3 ;
 ANTENNADIFFAREA                          0.160 LAYER ME4 ;
 ANTENNAMAXAREACAR                       48.616 LAYER ME2 ;
 ANTENNAMAXAREACAR                       57.875 LAYER ME3 ;
 ANTENNAMAXAREACAR                       67.134 LAYER ME4 ;
END DI49
PIN DO48
  DIRECTION OUTPUT ;
 PORT
  LAYER ME4 ;
  RECT 1004.800 0.000 1005.600 1.000 ;
  LAYER ME3 ;
  RECT 1004.800 0.000 1005.600 1.000 ;
  LAYER ME2 ;
  RECT 1004.800 0.000 1005.600 1.000 ;
  LAYER ME1 ;
  RECT 1004.800 0.000 1005.600 1.000 ;
 END
 ANTENNAPARTIALMETALAREA                  4.156 LAYER ME2 ;
 ANTENNADIFFAREA                          5.472 LAYER ME2 ;
 ANTENNADIFFAREA                          5.472 LAYER ME3 ;
 ANTENNADIFFAREA                          5.472 LAYER ME4 ;
END DO48
PIN WEB3
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 992.000 0.000 992.800 1.000 ;
  LAYER ME3 ;
  RECT 992.000 0.000 992.800 1.000 ;
  LAYER ME2 ;
  RECT 992.000 0.000 992.800 1.000 ;
  LAYER ME1 ;
  RECT 992.000 0.000 992.800 1.000 ;
 END
 ANTENNAPARTIALMETALAREA                  2.836 LAYER ME2 ;
 ANTENNAGATEAREA                          0.072 LAYER ME2 ;
 ANTENNAGATEAREA                          0.072 LAYER ME3 ;
 ANTENNAGATEAREA                          0.072 LAYER ME4 ;
 ANTENNADIFFAREA                          0.160 LAYER ME2 ;
 ANTENNADIFFAREA                          0.160 LAYER ME3 ;
 ANTENNADIFFAREA                          0.160 LAYER ME4 ;
 ANTENNAMAXAREACAR                       54.400 LAYER ME2 ;
 ANTENNAMAXAREACAR                       65.511 LAYER ME3 ;
 ANTENNAMAXAREACAR                       76.622 LAYER ME4 ;
END WEB3
PIN DI48
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 990.400 0.000 991.200 1.000 ;
  LAYER ME3 ;
  RECT 990.400 0.000 991.200 1.000 ;
  LAYER ME2 ;
  RECT 990.400 0.000 991.200 1.000 ;
  LAYER ME1 ;
  RECT 990.400 0.000 991.200 1.000 ;
 END
 ANTENNAPARTIALMETALAREA                  3.146 LAYER ME2 ;
 ANTENNAGATEAREA                          0.086 LAYER ME2 ;
 ANTENNAGATEAREA                          0.086 LAYER ME3 ;
 ANTENNAGATEAREA                          0.086 LAYER ME4 ;
 ANTENNADIFFAREA                          0.160 LAYER ME2 ;
 ANTENNADIFFAREA                          0.160 LAYER ME3 ;
 ANTENNADIFFAREA                          0.160 LAYER ME4 ;
 ANTENNAMAXAREACAR                       48.755 LAYER ME2 ;
 ANTENNAMAXAREACAR                       58.014 LAYER ME3 ;
 ANTENNAMAXAREACAR                       67.273 LAYER ME4 ;
END DI48
PIN DO47
  DIRECTION OUTPUT ;
 PORT
  LAYER ME4 ;
  RECT 983.600 0.000 984.400 1.000 ;
  LAYER ME3 ;
  RECT 983.600 0.000 984.400 1.000 ;
  LAYER ME2 ;
  RECT 983.600 0.000 984.400 1.000 ;
  LAYER ME1 ;
  RECT 983.600 0.000 984.400 1.000 ;
 END
 ANTENNAPARTIALMETALAREA                  4.180 LAYER ME2 ;
 ANTENNADIFFAREA                          5.472 LAYER ME2 ;
 ANTENNADIFFAREA                          5.472 LAYER ME3 ;
 ANTENNADIFFAREA                          5.472 LAYER ME4 ;
END DO47
PIN DI47
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 969.200 0.000 970.000 1.000 ;
  LAYER ME3 ;
  RECT 969.200 0.000 970.000 1.000 ;
  LAYER ME2 ;
  RECT 969.200 0.000 970.000 1.000 ;
  LAYER ME1 ;
  RECT 969.200 0.000 970.000 1.000 ;
 END
 ANTENNAPARTIALMETALAREA                  3.122 LAYER ME2 ;
 ANTENNAGATEAREA                          0.086 LAYER ME2 ;
 ANTENNAGATEAREA                          0.086 LAYER ME3 ;
 ANTENNAGATEAREA                          0.086 LAYER ME4 ;
 ANTENNADIFFAREA                          0.160 LAYER ME2 ;
 ANTENNADIFFAREA                          0.160 LAYER ME3 ;
 ANTENNADIFFAREA                          0.160 LAYER ME4 ;
 ANTENNAMAXAREACAR                       48.477 LAYER ME2 ;
 ANTENNAMAXAREACAR                       57.736 LAYER ME3 ;
 ANTENNAMAXAREACAR                       66.995 LAYER ME4 ;
END DI47
PIN DO46
  DIRECTION OUTPUT ;
 PORT
  LAYER ME4 ;
  RECT 964.000 0.000 964.800 1.000 ;
  LAYER ME3 ;
  RECT 964.000 0.000 964.800 1.000 ;
  LAYER ME2 ;
  RECT 964.000 0.000 964.800 1.000 ;
  LAYER ME1 ;
  RECT 964.000 0.000 964.800 1.000 ;
 END
 ANTENNAPARTIALMETALAREA                  4.148 LAYER ME2 ;
 ANTENNADIFFAREA                          5.472 LAYER ME2 ;
 ANTENNADIFFAREA                          5.472 LAYER ME3 ;
 ANTENNADIFFAREA                          5.472 LAYER ME4 ;
END DO46
PIN DI46
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 949.200 0.000 950.000 1.000 ;
  LAYER ME3 ;
  RECT 949.200 0.000 950.000 1.000 ;
  LAYER ME2 ;
  RECT 949.200 0.000 950.000 1.000 ;
  LAYER ME1 ;
  RECT 949.200 0.000 950.000 1.000 ;
 END
 ANTENNAPARTIALMETALAREA                  3.142 LAYER ME2 ;
 ANTENNAGATEAREA                          0.086 LAYER ME2 ;
 ANTENNAGATEAREA                          0.086 LAYER ME3 ;
 ANTENNAGATEAREA                          0.086 LAYER ME4 ;
 ANTENNADIFFAREA                          0.160 LAYER ME2 ;
 ANTENNADIFFAREA                          0.160 LAYER ME3 ;
 ANTENNADIFFAREA                          0.160 LAYER ME4 ;
 ANTENNAMAXAREACAR                       48.708 LAYER ME2 ;
 ANTENNAMAXAREACAR                       57.968 LAYER ME3 ;
 ANTENNAMAXAREACAR                       67.227 LAYER ME4 ;
END DI46
PIN DO45
  DIRECTION OUTPUT ;
 PORT
  LAYER ME4 ;
  RECT 942.800 0.000 943.600 1.000 ;
  LAYER ME3 ;
  RECT 942.800 0.000 943.600 1.000 ;
  LAYER ME2 ;
  RECT 942.800 0.000 943.600 1.000 ;
  LAYER ME1 ;
  RECT 942.800 0.000 943.600 1.000 ;
 END
 ANTENNAPARTIALMETALAREA                  4.156 LAYER ME2 ;
 ANTENNADIFFAREA                          5.472 LAYER ME2 ;
 ANTENNADIFFAREA                          5.472 LAYER ME3 ;
 ANTENNADIFFAREA                          5.472 LAYER ME4 ;
END DO45
PIN DI45
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 928.400 0.000 929.200 1.000 ;
  LAYER ME3 ;
  RECT 928.400 0.000 929.200 1.000 ;
  LAYER ME2 ;
  RECT 928.400 0.000 929.200 1.000 ;
  LAYER ME1 ;
  RECT 928.400 0.000 929.200 1.000 ;
 END
 ANTENNAPARTIALMETALAREA                  3.146 LAYER ME2 ;
 ANTENNAGATEAREA                          0.086 LAYER ME2 ;
 ANTENNAGATEAREA                          0.086 LAYER ME3 ;
 ANTENNAGATEAREA                          0.086 LAYER ME4 ;
 ANTENNADIFFAREA                          0.160 LAYER ME2 ;
 ANTENNADIFFAREA                          0.160 LAYER ME3 ;
 ANTENNADIFFAREA                          0.160 LAYER ME4 ;
 ANTENNAMAXAREACAR                       48.755 LAYER ME2 ;
 ANTENNAMAXAREACAR                       58.014 LAYER ME3 ;
 ANTENNAMAXAREACAR                       67.273 LAYER ME4 ;
END DI45
PIN DO44
  DIRECTION OUTPUT ;
 PORT
  LAYER ME4 ;
  RECT 923.200 0.000 924.000 1.000 ;
  LAYER ME3 ;
  RECT 923.200 0.000 924.000 1.000 ;
  LAYER ME2 ;
  RECT 923.200 0.000 924.000 1.000 ;
  LAYER ME1 ;
  RECT 923.200 0.000 924.000 1.000 ;
 END
 ANTENNAPARTIALMETALAREA                  4.172 LAYER ME2 ;
 ANTENNADIFFAREA                          5.472 LAYER ME2 ;
 ANTENNADIFFAREA                          5.472 LAYER ME3 ;
 ANTENNADIFFAREA                          5.472 LAYER ME4 ;
END DO44
PIN DI44
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 908.400 0.000 909.200 1.000 ;
  LAYER ME3 ;
  RECT 908.400 0.000 909.200 1.000 ;
  LAYER ME2 ;
  RECT 908.400 0.000 909.200 1.000 ;
  LAYER ME1 ;
  RECT 908.400 0.000 909.200 1.000 ;
 END
 ANTENNAPARTIALMETALAREA                  3.118 LAYER ME2 ;
 ANTENNAGATEAREA                          0.086 LAYER ME2 ;
 ANTENNAGATEAREA                          0.086 LAYER ME3 ;
 ANTENNAGATEAREA                          0.086 LAYER ME4 ;
 ANTENNADIFFAREA                          0.160 LAYER ME2 ;
 ANTENNADIFFAREA                          0.160 LAYER ME3 ;
 ANTENNADIFFAREA                          0.160 LAYER ME4 ;
 ANTENNAMAXAREACAR                       48.431 LAYER ME2 ;
 ANTENNAMAXAREACAR                       57.690 LAYER ME3 ;
 ANTENNAMAXAREACAR                       66.949 LAYER ME4 ;
END DI44
PIN DO43
  DIRECTION OUTPUT ;
 PORT
  LAYER ME4 ;
  RECT 902.000 0.000 902.800 1.000 ;
  LAYER ME3 ;
  RECT 902.000 0.000 902.800 1.000 ;
  LAYER ME2 ;
  RECT 902.000 0.000 902.800 1.000 ;
  LAYER ME1 ;
  RECT 902.000 0.000 902.800 1.000 ;
 END
 ANTENNAPARTIALMETALAREA                  4.148 LAYER ME2 ;
 ANTENNADIFFAREA                          5.472 LAYER ME2 ;
 ANTENNADIFFAREA                          5.472 LAYER ME3 ;
 ANTENNADIFFAREA                          5.472 LAYER ME4 ;
END DO43
PIN DI43
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 887.200 0.000 888.000 1.000 ;
  LAYER ME3 ;
  RECT 887.200 0.000 888.000 1.000 ;
  LAYER ME2 ;
  RECT 887.200 0.000 888.000 1.000 ;
  LAYER ME1 ;
  RECT 887.200 0.000 888.000 1.000 ;
 END
 ANTENNAPARTIALMETALAREA                  3.142 LAYER ME2 ;
 ANTENNAGATEAREA                          0.086 LAYER ME2 ;
 ANTENNAGATEAREA                          0.086 LAYER ME3 ;
 ANTENNAGATEAREA                          0.086 LAYER ME4 ;
 ANTENNADIFFAREA                          0.160 LAYER ME2 ;
 ANTENNADIFFAREA                          0.160 LAYER ME3 ;
 ANTENNADIFFAREA                          0.160 LAYER ME4 ;
 ANTENNAMAXAREACAR                       48.708 LAYER ME2 ;
 ANTENNAMAXAREACAR                       57.968 LAYER ME3 ;
 ANTENNAMAXAREACAR                       67.227 LAYER ME4 ;
END DI43
PIN DO42
  DIRECTION OUTPUT ;
 PORT
  LAYER ME4 ;
  RECT 882.000 0.000 882.800 1.000 ;
  LAYER ME3 ;
  RECT 882.000 0.000 882.800 1.000 ;
  LAYER ME2 ;
  RECT 882.000 0.000 882.800 1.000 ;
  LAYER ME1 ;
  RECT 882.000 0.000 882.800 1.000 ;
 END
 ANTENNAPARTIALMETALAREA                  4.164 LAYER ME2 ;
 ANTENNADIFFAREA                          5.472 LAYER ME2 ;
 ANTENNADIFFAREA                          5.472 LAYER ME3 ;
 ANTENNADIFFAREA                          5.472 LAYER ME4 ;
END DO42
PIN DI42
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 867.600 0.000 868.400 1.000 ;
  LAYER ME3 ;
  RECT 867.600 0.000 868.400 1.000 ;
  LAYER ME2 ;
  RECT 867.600 0.000 868.400 1.000 ;
  LAYER ME1 ;
  RECT 867.600 0.000 868.400 1.000 ;
 END
 ANTENNAPARTIALMETALAREA                  3.138 LAYER ME2 ;
 ANTENNAGATEAREA                          0.086 LAYER ME2 ;
 ANTENNAGATEAREA                          0.086 LAYER ME3 ;
 ANTENNAGATEAREA                          0.086 LAYER ME4 ;
 ANTENNADIFFAREA                          0.160 LAYER ME2 ;
 ANTENNADIFFAREA                          0.160 LAYER ME3 ;
 ANTENNADIFFAREA                          0.160 LAYER ME4 ;
 ANTENNAMAXAREACAR                       48.662 LAYER ME2 ;
 ANTENNAMAXAREACAR                       57.921 LAYER ME3 ;
 ANTENNAMAXAREACAR                       67.181 LAYER ME4 ;
END DI42
PIN DO41
  DIRECTION OUTPUT ;
 PORT
  LAYER ME4 ;
  RECT 861.200 0.000 862.000 1.000 ;
  LAYER ME3 ;
  RECT 861.200 0.000 862.000 1.000 ;
  LAYER ME2 ;
  RECT 861.200 0.000 862.000 1.000 ;
  LAYER ME1 ;
  RECT 861.200 0.000 862.000 1.000 ;
 END
 ANTENNAPARTIALMETALAREA                  4.172 LAYER ME2 ;
 ANTENNADIFFAREA                          5.472 LAYER ME2 ;
 ANTENNADIFFAREA                          5.472 LAYER ME3 ;
 ANTENNADIFFAREA                          5.472 LAYER ME4 ;
END DO41
PIN DI41
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 846.400 0.000 847.200 1.000 ;
  LAYER ME3 ;
  RECT 846.400 0.000 847.200 1.000 ;
  LAYER ME2 ;
  RECT 846.400 0.000 847.200 1.000 ;
  LAYER ME1 ;
  RECT 846.400 0.000 847.200 1.000 ;
 END
 ANTENNAPARTIALMETALAREA                  3.118 LAYER ME2 ;
 ANTENNAGATEAREA                          0.086 LAYER ME2 ;
 ANTENNAGATEAREA                          0.086 LAYER ME3 ;
 ANTENNAGATEAREA                          0.086 LAYER ME4 ;
 ANTENNADIFFAREA                          0.160 LAYER ME2 ;
 ANTENNADIFFAREA                          0.160 LAYER ME3 ;
 ANTENNADIFFAREA                          0.160 LAYER ME4 ;
 ANTENNAMAXAREACAR                       48.431 LAYER ME2 ;
 ANTENNAMAXAREACAR                       57.690 LAYER ME3 ;
 ANTENNAMAXAREACAR                       66.949 LAYER ME4 ;
END DI41
PIN DO40
  DIRECTION OUTPUT ;
 PORT
  LAYER ME4 ;
  RECT 841.200 0.000 842.000 1.000 ;
  LAYER ME3 ;
  RECT 841.200 0.000 842.000 1.000 ;
  LAYER ME2 ;
  RECT 841.200 0.000 842.000 1.000 ;
  LAYER ME1 ;
  RECT 841.200 0.000 842.000 1.000 ;
 END
 ANTENNAPARTIALMETALAREA                  4.140 LAYER ME2 ;
 ANTENNADIFFAREA                          5.472 LAYER ME2 ;
 ANTENNADIFFAREA                          5.472 LAYER ME3 ;
 ANTENNADIFFAREA                          5.472 LAYER ME4 ;
END DO40
PIN DI40
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 826.400 0.000 827.200 1.000 ;
  LAYER ME3 ;
  RECT 826.400 0.000 827.200 1.000 ;
  LAYER ME2 ;
  RECT 826.400 0.000 827.200 1.000 ;
  LAYER ME1 ;
  RECT 826.400 0.000 827.200 1.000 ;
 END
 ANTENNAPARTIALMETALAREA                  3.150 LAYER ME2 ;
 ANTENNAGATEAREA                          0.086 LAYER ME2 ;
 ANTENNAGATEAREA                          0.086 LAYER ME3 ;
 ANTENNAGATEAREA                          0.086 LAYER ME4 ;
 ANTENNADIFFAREA                          0.160 LAYER ME2 ;
 ANTENNADIFFAREA                          0.160 LAYER ME3 ;
 ANTENNADIFFAREA                          0.160 LAYER ME4 ;
 ANTENNAMAXAREACAR                       48.801 LAYER ME2 ;
 ANTENNAMAXAREACAR                       58.060 LAYER ME3 ;
 ANTENNAMAXAREACAR                       67.319 LAYER ME4 ;
END DI40
PIN DO39
  DIRECTION OUTPUT ;
 PORT
  LAYER ME4 ;
  RECT 820.000 0.000 820.800 1.000 ;
  LAYER ME3 ;
  RECT 820.000 0.000 820.800 1.000 ;
  LAYER ME2 ;
  RECT 820.000 0.000 820.800 1.000 ;
  LAYER ME1 ;
  RECT 820.000 0.000 820.800 1.000 ;
 END
 ANTENNAPARTIALMETALAREA                  4.164 LAYER ME2 ;
 ANTENNADIFFAREA                          5.472 LAYER ME2 ;
 ANTENNADIFFAREA                          5.472 LAYER ME3 ;
 ANTENNADIFFAREA                          5.472 LAYER ME4 ;
END DO39
PIN DI39
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 805.600 0.000 806.400 1.000 ;
  LAYER ME3 ;
  RECT 805.600 0.000 806.400 1.000 ;
  LAYER ME2 ;
  RECT 805.600 0.000 806.400 1.000 ;
  LAYER ME1 ;
  RECT 805.600 0.000 806.400 1.000 ;
 END
 ANTENNAPARTIALMETALAREA                  3.138 LAYER ME2 ;
 ANTENNAGATEAREA                          0.086 LAYER ME2 ;
 ANTENNAGATEAREA                          0.086 LAYER ME3 ;
 ANTENNAGATEAREA                          0.086 LAYER ME4 ;
 ANTENNADIFFAREA                          0.160 LAYER ME2 ;
 ANTENNADIFFAREA                          0.160 LAYER ME3 ;
 ANTENNADIFFAREA                          0.160 LAYER ME4 ;
 ANTENNAMAXAREACAR                       48.662 LAYER ME2 ;
 ANTENNAMAXAREACAR                       57.921 LAYER ME3 ;
 ANTENNAMAXAREACAR                       67.181 LAYER ME4 ;
END DI39
PIN DO38
  DIRECTION OUTPUT ;
 PORT
  LAYER ME4 ;
  RECT 800.400 0.000 801.200 1.000 ;
  LAYER ME3 ;
  RECT 800.400 0.000 801.200 1.000 ;
  LAYER ME2 ;
  RECT 800.400 0.000 801.200 1.000 ;
  LAYER ME1 ;
  RECT 800.400 0.000 801.200 1.000 ;
 END
 ANTENNAPARTIALMETALAREA                  4.164 LAYER ME2 ;
 ANTENNADIFFAREA                          5.472 LAYER ME2 ;
 ANTENNADIFFAREA                          5.472 LAYER ME3 ;
 ANTENNADIFFAREA                          5.472 LAYER ME4 ;
END DO38
PIN DI38
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 785.600 0.000 786.400 1.000 ;
  LAYER ME3 ;
  RECT 785.600 0.000 786.400 1.000 ;
  LAYER ME2 ;
  RECT 785.600 0.000 786.400 1.000 ;
  LAYER ME1 ;
  RECT 785.600 0.000 786.400 1.000 ;
 END
 ANTENNAPARTIALMETALAREA                  3.126 LAYER ME2 ;
 ANTENNAGATEAREA                          0.086 LAYER ME2 ;
 ANTENNAGATEAREA                          0.086 LAYER ME3 ;
 ANTENNAGATEAREA                          0.086 LAYER ME4 ;
 ANTENNADIFFAREA                          0.160 LAYER ME2 ;
 ANTENNADIFFAREA                          0.160 LAYER ME3 ;
 ANTENNADIFFAREA                          0.160 LAYER ME4 ;
 ANTENNAMAXAREACAR                       48.523 LAYER ME2 ;
 ANTENNAMAXAREACAR                       57.782 LAYER ME3 ;
 ANTENNAMAXAREACAR                       67.042 LAYER ME4 ;
END DI38
PIN DO37
  DIRECTION OUTPUT ;
 PORT
  LAYER ME4 ;
  RECT 779.200 0.000 780.000 1.000 ;
  LAYER ME3 ;
  RECT 779.200 0.000 780.000 1.000 ;
  LAYER ME2 ;
  RECT 779.200 0.000 780.000 1.000 ;
  LAYER ME1 ;
  RECT 779.200 0.000 780.000 1.000 ;
 END
 ANTENNAPARTIALMETALAREA                  4.140 LAYER ME2 ;
 ANTENNADIFFAREA                          5.472 LAYER ME2 ;
 ANTENNADIFFAREA                          5.472 LAYER ME3 ;
 ANTENNADIFFAREA                          5.472 LAYER ME4 ;
END DO37
PIN DI37
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 764.400 0.000 765.200 1.000 ;
  LAYER ME3 ;
  RECT 764.400 0.000 765.200 1.000 ;
  LAYER ME2 ;
  RECT 764.400 0.000 765.200 1.000 ;
  LAYER ME1 ;
  RECT 764.400 0.000 765.200 1.000 ;
 END
 ANTENNAPARTIALMETALAREA                  3.150 LAYER ME2 ;
 ANTENNAGATEAREA                          0.086 LAYER ME2 ;
 ANTENNAGATEAREA                          0.086 LAYER ME3 ;
 ANTENNAGATEAREA                          0.086 LAYER ME4 ;
 ANTENNADIFFAREA                          0.160 LAYER ME2 ;
 ANTENNADIFFAREA                          0.160 LAYER ME3 ;
 ANTENNADIFFAREA                          0.160 LAYER ME4 ;
 ANTENNAMAXAREACAR                       48.801 LAYER ME2 ;
 ANTENNAMAXAREACAR                       58.060 LAYER ME3 ;
 ANTENNAMAXAREACAR                       67.319 LAYER ME4 ;
END DI37
PIN DO36
  DIRECTION OUTPUT ;
 PORT
  LAYER ME4 ;
  RECT 759.200 0.000 760.000 1.000 ;
  LAYER ME3 ;
  RECT 759.200 0.000 760.000 1.000 ;
  LAYER ME2 ;
  RECT 759.200 0.000 760.000 1.000 ;
  LAYER ME1 ;
  RECT 759.200 0.000 760.000 1.000 ;
 END
 ANTENNAPARTIALMETALAREA                  4.172 LAYER ME2 ;
 ANTENNADIFFAREA                          5.472 LAYER ME2 ;
 ANTENNADIFFAREA                          5.472 LAYER ME3 ;
 ANTENNADIFFAREA                          5.472 LAYER ME4 ;
END DO36
PIN DI36
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 744.800 0.000 745.600 1.000 ;
  LAYER ME3 ;
  RECT 744.800 0.000 745.600 1.000 ;
  LAYER ME2 ;
  RECT 744.800 0.000 745.600 1.000 ;
  LAYER ME1 ;
  RECT 744.800 0.000 745.600 1.000 ;
 END
 ANTENNAPARTIALMETALAREA                  3.130 LAYER ME2 ;
 ANTENNAGATEAREA                          0.086 LAYER ME2 ;
 ANTENNAGATEAREA                          0.086 LAYER ME3 ;
 ANTENNAGATEAREA                          0.086 LAYER ME4 ;
 ANTENNADIFFAREA                          0.160 LAYER ME2 ;
 ANTENNADIFFAREA                          0.160 LAYER ME3 ;
 ANTENNADIFFAREA                          0.160 LAYER ME4 ;
 ANTENNAMAXAREACAR                       48.569 LAYER ME2 ;
 ANTENNAMAXAREACAR                       57.829 LAYER ME3 ;
 ANTENNAMAXAREACAR                       67.088 LAYER ME4 ;
END DI36
PIN DO35
  DIRECTION OUTPUT ;
 PORT
  LAYER ME4 ;
  RECT 738.400 0.000 739.200 1.000 ;
  LAYER ME3 ;
  RECT 738.400 0.000 739.200 1.000 ;
  LAYER ME2 ;
  RECT 738.400 0.000 739.200 1.000 ;
  LAYER ME1 ;
  RECT 738.400 0.000 739.200 1.000 ;
 END
 ANTENNAPARTIALMETALAREA                  4.164 LAYER ME2 ;
 ANTENNADIFFAREA                          5.472 LAYER ME2 ;
 ANTENNADIFFAREA                          5.472 LAYER ME3 ;
 ANTENNADIFFAREA                          5.472 LAYER ME4 ;
END DO35
PIN DI35
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 723.600 0.000 724.400 1.000 ;
  LAYER ME3 ;
  RECT 723.600 0.000 724.400 1.000 ;
  LAYER ME2 ;
  RECT 723.600 0.000 724.400 1.000 ;
  LAYER ME1 ;
  RECT 723.600 0.000 724.400 1.000 ;
 END
 ANTENNAPARTIALMETALAREA                  3.126 LAYER ME2 ;
 ANTENNAGATEAREA                          0.086 LAYER ME2 ;
 ANTENNAGATEAREA                          0.086 LAYER ME3 ;
 ANTENNAGATEAREA                          0.086 LAYER ME4 ;
 ANTENNADIFFAREA                          0.160 LAYER ME2 ;
 ANTENNADIFFAREA                          0.160 LAYER ME3 ;
 ANTENNADIFFAREA                          0.160 LAYER ME4 ;
 ANTENNAMAXAREACAR                       48.523 LAYER ME2 ;
 ANTENNAMAXAREACAR                       57.782 LAYER ME3 ;
 ANTENNAMAXAREACAR                       67.042 LAYER ME4 ;
END DI35
PIN DO34
  DIRECTION OUTPUT ;
 PORT
  LAYER ME4 ;
  RECT 718.400 0.000 719.200 1.000 ;
  LAYER ME3 ;
  RECT 718.400 0.000 719.200 1.000 ;
  LAYER ME2 ;
  RECT 718.400 0.000 719.200 1.000 ;
  LAYER ME1 ;
  RECT 718.400 0.000 719.200 1.000 ;
 END
 ANTENNAPARTIALMETALAREA                  4.148 LAYER ME2 ;
 ANTENNADIFFAREA                          5.472 LAYER ME2 ;
 ANTENNADIFFAREA                          5.472 LAYER ME3 ;
 ANTENNADIFFAREA                          5.472 LAYER ME4 ;
END DO34
PIN DI34
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 704.000 0.000 704.800 1.000 ;
  LAYER ME3 ;
  RECT 704.000 0.000 704.800 1.000 ;
  LAYER ME2 ;
  RECT 704.000 0.000 704.800 1.000 ;
  LAYER ME1 ;
  RECT 704.000 0.000 704.800 1.000 ;
 END
 ANTENNAPARTIALMETALAREA                  3.154 LAYER ME2 ;
 ANTENNAGATEAREA                          0.086 LAYER ME2 ;
 ANTENNAGATEAREA                          0.086 LAYER ME3 ;
 ANTENNAGATEAREA                          0.086 LAYER ME4 ;
 ANTENNADIFFAREA                          0.160 LAYER ME2 ;
 ANTENNADIFFAREA                          0.160 LAYER ME3 ;
 ANTENNADIFFAREA                          0.160 LAYER ME4 ;
 ANTENNAMAXAREACAR                       48.847 LAYER ME2 ;
 ANTENNAMAXAREACAR                       58.106 LAYER ME3 ;
 ANTENNAMAXAREACAR                       67.366 LAYER ME4 ;
END DI34
PIN DO33
  DIRECTION OUTPUT ;
 PORT
  LAYER ME4 ;
  RECT 697.200 0.000 698.000 1.000 ;
  LAYER ME3 ;
  RECT 697.200 0.000 698.000 1.000 ;
  LAYER ME2 ;
  RECT 697.200 0.000 698.000 1.000 ;
  LAYER ME1 ;
  RECT 697.200 0.000 698.000 1.000 ;
 END
 ANTENNAPARTIALMETALAREA                  4.172 LAYER ME2 ;
 ANTENNADIFFAREA                          5.472 LAYER ME2 ;
 ANTENNADIFFAREA                          5.472 LAYER ME3 ;
 ANTENNADIFFAREA                          5.472 LAYER ME4 ;
END DO33
PIN DI33
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 682.800 0.000 683.600 1.000 ;
  LAYER ME3 ;
  RECT 682.800 0.000 683.600 1.000 ;
  LAYER ME2 ;
  RECT 682.800 0.000 683.600 1.000 ;
  LAYER ME1 ;
  RECT 682.800 0.000 683.600 1.000 ;
 END
 ANTENNAPARTIALMETALAREA                  3.130 LAYER ME2 ;
 ANTENNAGATEAREA                          0.086 LAYER ME2 ;
 ANTENNAGATEAREA                          0.086 LAYER ME3 ;
 ANTENNAGATEAREA                          0.086 LAYER ME4 ;
 ANTENNADIFFAREA                          0.160 LAYER ME2 ;
 ANTENNADIFFAREA                          0.160 LAYER ME3 ;
 ANTENNADIFFAREA                          0.160 LAYER ME4 ;
 ANTENNAMAXAREACAR                       48.569 LAYER ME2 ;
 ANTENNAMAXAREACAR                       57.829 LAYER ME3 ;
 ANTENNAMAXAREACAR                       67.088 LAYER ME4 ;
END DI33
PIN DO32
  DIRECTION OUTPUT ;
 PORT
  LAYER ME4 ;
  RECT 677.600 0.000 678.400 1.000 ;
  LAYER ME3 ;
  RECT 677.600 0.000 678.400 1.000 ;
  LAYER ME2 ;
  RECT 677.600 0.000 678.400 1.000 ;
  LAYER ME1 ;
  RECT 677.600 0.000 678.400 1.000 ;
 END
 ANTENNAPARTIALMETALAREA                  4.156 LAYER ME2 ;
 ANTENNADIFFAREA                          5.472 LAYER ME2 ;
 ANTENNADIFFAREA                          5.472 LAYER ME3 ;
 ANTENNADIFFAREA                          5.472 LAYER ME4 ;
END DO32
PIN WEB2
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 664.800 0.000 665.600 1.000 ;
  LAYER ME3 ;
  RECT 664.800 0.000 665.600 1.000 ;
  LAYER ME2 ;
  RECT 664.800 0.000 665.600 1.000 ;
  LAYER ME1 ;
  RECT 664.800 0.000 665.600 1.000 ;
 END
 ANTENNAPARTIALMETALAREA                  2.868 LAYER ME2 ;
 ANTENNAGATEAREA                          0.072 LAYER ME2 ;
 ANTENNAGATEAREA                          0.072 LAYER ME3 ;
 ANTENNAGATEAREA                          0.072 LAYER ME4 ;
 ANTENNADIFFAREA                          0.160 LAYER ME2 ;
 ANTENNADIFFAREA                          0.160 LAYER ME3 ;
 ANTENNADIFFAREA                          0.160 LAYER ME4 ;
 ANTENNAMAXAREACAR                       54.844 LAYER ME2 ;
 ANTENNAMAXAREACAR                       65.956 LAYER ME3 ;
 ANTENNAMAXAREACAR                       77.067 LAYER ME4 ;
END WEB2
PIN DI32
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 662.800 0.000 663.600 1.000 ;
  LAYER ME3 ;
  RECT 662.800 0.000 663.600 1.000 ;
  LAYER ME2 ;
  RECT 662.800 0.000 663.600 1.000 ;
  LAYER ME1 ;
  RECT 662.800 0.000 663.600 1.000 ;
 END
 ANTENNAPARTIALMETALAREA                  3.134 LAYER ME2 ;
 ANTENNAGATEAREA                          0.086 LAYER ME2 ;
 ANTENNAGATEAREA                          0.086 LAYER ME3 ;
 ANTENNAGATEAREA                          0.086 LAYER ME4 ;
 ANTENNADIFFAREA                          0.160 LAYER ME2 ;
 ANTENNADIFFAREA                          0.160 LAYER ME3 ;
 ANTENNADIFFAREA                          0.160 LAYER ME4 ;
 ANTENNAMAXAREACAR                       48.616 LAYER ME2 ;
 ANTENNAMAXAREACAR                       57.875 LAYER ME3 ;
 ANTENNAMAXAREACAR                       67.134 LAYER ME4 ;
END DI32
PIN DO31
  DIRECTION OUTPUT ;
 PORT
  LAYER ME4 ;
  RECT 656.400 0.000 657.200 1.000 ;
  LAYER ME3 ;
  RECT 656.400 0.000 657.200 1.000 ;
  LAYER ME2 ;
  RECT 656.400 0.000 657.200 1.000 ;
  LAYER ME1 ;
  RECT 656.400 0.000 657.200 1.000 ;
 END
 ANTENNAPARTIALMETALAREA                  4.148 LAYER ME2 ;
 ANTENNADIFFAREA                          5.472 LAYER ME2 ;
 ANTENNADIFFAREA                          5.472 LAYER ME3 ;
 ANTENNADIFFAREA                          5.472 LAYER ME4 ;
END DO31
PIN DI31
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 642.000 0.000 642.800 1.000 ;
  LAYER ME3 ;
  RECT 642.000 0.000 642.800 1.000 ;
  LAYER ME2 ;
  RECT 642.000 0.000 642.800 1.000 ;
  LAYER ME1 ;
  RECT 642.000 0.000 642.800 1.000 ;
 END
 ANTENNAPARTIALMETALAREA                  3.154 LAYER ME2 ;
 ANTENNAGATEAREA                          0.086 LAYER ME2 ;
 ANTENNAGATEAREA                          0.086 LAYER ME3 ;
 ANTENNAGATEAREA                          0.086 LAYER ME4 ;
 ANTENNADIFFAREA                          0.160 LAYER ME2 ;
 ANTENNADIFFAREA                          0.160 LAYER ME3 ;
 ANTENNADIFFAREA                          0.160 LAYER ME4 ;
 ANTENNAMAXAREACAR                       48.847 LAYER ME2 ;
 ANTENNAMAXAREACAR                       58.106 LAYER ME3 ;
 ANTENNAMAXAREACAR                       67.366 LAYER ME4 ;
END DI31
PIN DO30
  DIRECTION OUTPUT ;
 PORT
  LAYER ME4 ;
  RECT 636.400 0.000 637.200 1.000 ;
  LAYER ME3 ;
  RECT 636.400 0.000 637.200 1.000 ;
  LAYER ME2 ;
  RECT 636.400 0.000 637.200 1.000 ;
  LAYER ME1 ;
  RECT 636.400 0.000 637.200 1.000 ;
 END
 ANTENNAPARTIALMETALAREA                  4.180 LAYER ME2 ;
 ANTENNADIFFAREA                          5.472 LAYER ME2 ;
 ANTENNADIFFAREA                          5.472 LAYER ME3 ;
 ANTENNADIFFAREA                          5.472 LAYER ME4 ;
END DO30
PIN DI30
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 622.000 0.000 622.800 1.000 ;
  LAYER ME3 ;
  RECT 622.000 0.000 622.800 1.000 ;
  LAYER ME2 ;
  RECT 622.000 0.000 622.800 1.000 ;
  LAYER ME1 ;
  RECT 622.000 0.000 622.800 1.000 ;
 END
 ANTENNAPARTIALMETALAREA                  3.122 LAYER ME2 ;
 ANTENNAGATEAREA                          0.086 LAYER ME2 ;
 ANTENNAGATEAREA                          0.086 LAYER ME3 ;
 ANTENNAGATEAREA                          0.086 LAYER ME4 ;
 ANTENNADIFFAREA                          0.160 LAYER ME2 ;
 ANTENNADIFFAREA                          0.160 LAYER ME3 ;
 ANTENNADIFFAREA                          0.160 LAYER ME4 ;
 ANTENNAMAXAREACAR                       48.477 LAYER ME2 ;
 ANTENNAMAXAREACAR                       57.736 LAYER ME3 ;
 ANTENNAMAXAREACAR                       66.995 LAYER ME4 ;
END DI30
PIN DO29
  DIRECTION OUTPUT ;
 PORT
  LAYER ME4 ;
  RECT 615.600 0.000 616.400 1.000 ;
  LAYER ME3 ;
  RECT 615.600 0.000 616.400 1.000 ;
  LAYER ME2 ;
  RECT 615.600 0.000 616.400 1.000 ;
  LAYER ME1 ;
  RECT 615.600 0.000 616.400 1.000 ;
 END
 ANTENNAPARTIALMETALAREA                  4.156 LAYER ME2 ;
 ANTENNADIFFAREA                          5.472 LAYER ME2 ;
 ANTENNADIFFAREA                          5.472 LAYER ME3 ;
 ANTENNADIFFAREA                          5.472 LAYER ME4 ;
END DO29
PIN DI29
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 600.800 0.000 601.600 1.000 ;
  LAYER ME3 ;
  RECT 600.800 0.000 601.600 1.000 ;
  LAYER ME2 ;
  RECT 600.800 0.000 601.600 1.000 ;
  LAYER ME1 ;
  RECT 600.800 0.000 601.600 1.000 ;
 END
 ANTENNAPARTIALMETALAREA                  3.134 LAYER ME2 ;
 ANTENNAGATEAREA                          0.086 LAYER ME2 ;
 ANTENNAGATEAREA                          0.086 LAYER ME3 ;
 ANTENNAGATEAREA                          0.086 LAYER ME4 ;
 ANTENNADIFFAREA                          0.160 LAYER ME2 ;
 ANTENNADIFFAREA                          0.160 LAYER ME3 ;
 ANTENNADIFFAREA                          0.160 LAYER ME4 ;
 ANTENNAMAXAREACAR                       48.616 LAYER ME2 ;
 ANTENNAMAXAREACAR                       57.875 LAYER ME3 ;
 ANTENNAMAXAREACAR                       67.134 LAYER ME4 ;
END DI29
PIN DO28
  DIRECTION OUTPUT ;
 PORT
  LAYER ME4 ;
  RECT 595.600 0.000 596.400 1.000 ;
  LAYER ME3 ;
  RECT 595.600 0.000 596.400 1.000 ;
  LAYER ME2 ;
  RECT 595.600 0.000 596.400 1.000 ;
  LAYER ME1 ;
  RECT 595.600 0.000 596.400 1.000 ;
 END
 ANTENNAPARTIALMETALAREA                  4.156 LAYER ME2 ;
 ANTENNADIFFAREA                          5.472 LAYER ME2 ;
 ANTENNADIFFAREA                          5.472 LAYER ME3 ;
 ANTENNADIFFAREA                          5.472 LAYER ME4 ;
END DO28
PIN DI28
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 581.200 0.000 582.000 1.000 ;
  LAYER ME3 ;
  RECT 581.200 0.000 582.000 1.000 ;
  LAYER ME2 ;
  RECT 581.200 0.000 582.000 1.000 ;
  LAYER ME1 ;
  RECT 581.200 0.000 582.000 1.000 ;
 END
 ANTENNAPARTIALMETALAREA                  3.146 LAYER ME2 ;
 ANTENNAGATEAREA                          0.086 LAYER ME2 ;
 ANTENNAGATEAREA                          0.086 LAYER ME3 ;
 ANTENNAGATEAREA                          0.086 LAYER ME4 ;
 ANTENNADIFFAREA                          0.160 LAYER ME2 ;
 ANTENNADIFFAREA                          0.160 LAYER ME3 ;
 ANTENNADIFFAREA                          0.160 LAYER ME4 ;
 ANTENNAMAXAREACAR                       48.755 LAYER ME2 ;
 ANTENNAMAXAREACAR                       58.014 LAYER ME3 ;
 ANTENNAMAXAREACAR                       67.273 LAYER ME4 ;
END DI28
PIN DO27
  DIRECTION OUTPUT ;
 PORT
  LAYER ME4 ;
  RECT 574.400 0.000 575.200 1.000 ;
  LAYER ME3 ;
  RECT 574.400 0.000 575.200 1.000 ;
  LAYER ME2 ;
  RECT 574.400 0.000 575.200 1.000 ;
  LAYER ME1 ;
  RECT 574.400 0.000 575.200 1.000 ;
 END
 ANTENNAPARTIALMETALAREA                  4.180 LAYER ME2 ;
 ANTENNADIFFAREA                          5.472 LAYER ME2 ;
 ANTENNADIFFAREA                          5.472 LAYER ME3 ;
 ANTENNADIFFAREA                          5.472 LAYER ME4 ;
END DO27
PIN DI27
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 560.000 0.000 560.800 1.000 ;
  LAYER ME3 ;
  RECT 560.000 0.000 560.800 1.000 ;
  LAYER ME2 ;
  RECT 560.000 0.000 560.800 1.000 ;
  LAYER ME1 ;
  RECT 560.000 0.000 560.800 1.000 ;
 END
 ANTENNAPARTIALMETALAREA                  3.122 LAYER ME2 ;
 ANTENNAGATEAREA                          0.086 LAYER ME2 ;
 ANTENNAGATEAREA                          0.086 LAYER ME3 ;
 ANTENNAGATEAREA                          0.086 LAYER ME4 ;
 ANTENNADIFFAREA                          0.160 LAYER ME2 ;
 ANTENNADIFFAREA                          0.160 LAYER ME3 ;
 ANTENNADIFFAREA                          0.160 LAYER ME4 ;
 ANTENNAMAXAREACAR                       48.477 LAYER ME2 ;
 ANTENNAMAXAREACAR                       57.736 LAYER ME3 ;
 ANTENNAMAXAREACAR                       66.995 LAYER ME4 ;
END DI27
PIN DO26
  DIRECTION OUTPUT ;
 PORT
  LAYER ME4 ;
  RECT 554.800 0.000 555.600 1.000 ;
  LAYER ME3 ;
  RECT 554.800 0.000 555.600 1.000 ;
  LAYER ME2 ;
  RECT 554.800 0.000 555.600 1.000 ;
  LAYER ME1 ;
  RECT 554.800 0.000 555.600 1.000 ;
 END
 ANTENNAPARTIALMETALAREA                  4.148 LAYER ME2 ;
 ANTENNADIFFAREA                          5.472 LAYER ME2 ;
 ANTENNADIFFAREA                          5.472 LAYER ME3 ;
 ANTENNADIFFAREA                          5.472 LAYER ME4 ;
END DO26
PIN DI26
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 540.000 0.000 540.800 1.000 ;
  LAYER ME3 ;
  RECT 540.000 0.000 540.800 1.000 ;
  LAYER ME2 ;
  RECT 540.000 0.000 540.800 1.000 ;
  LAYER ME1 ;
  RECT 540.000 0.000 540.800 1.000 ;
 END
 ANTENNAPARTIALMETALAREA                  3.142 LAYER ME2 ;
 ANTENNAGATEAREA                          0.086 LAYER ME2 ;
 ANTENNAGATEAREA                          0.086 LAYER ME3 ;
 ANTENNAGATEAREA                          0.086 LAYER ME4 ;
 ANTENNADIFFAREA                          0.160 LAYER ME2 ;
 ANTENNADIFFAREA                          0.160 LAYER ME3 ;
 ANTENNADIFFAREA                          0.160 LAYER ME4 ;
 ANTENNAMAXAREACAR                       48.708 LAYER ME2 ;
 ANTENNAMAXAREACAR                       57.968 LAYER ME3 ;
 ANTENNAMAXAREACAR                       67.227 LAYER ME4 ;
END DI26
PIN DO25
  DIRECTION OUTPUT ;
 PORT
  LAYER ME4 ;
  RECT 533.600 0.000 534.400 1.000 ;
  LAYER ME3 ;
  RECT 533.600 0.000 534.400 1.000 ;
  LAYER ME2 ;
  RECT 533.600 0.000 534.400 1.000 ;
  LAYER ME1 ;
  RECT 533.600 0.000 534.400 1.000 ;
 END
 ANTENNAPARTIALMETALAREA                  4.156 LAYER ME2 ;
 ANTENNADIFFAREA                          5.472 LAYER ME2 ;
 ANTENNADIFFAREA                          5.472 LAYER ME3 ;
 ANTENNADIFFAREA                          5.472 LAYER ME4 ;
END DO25
PIN DI25
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 519.200 0.000 520.000 1.000 ;
  LAYER ME3 ;
  RECT 519.200 0.000 520.000 1.000 ;
  LAYER ME2 ;
  RECT 519.200 0.000 520.000 1.000 ;
  LAYER ME1 ;
  RECT 519.200 0.000 520.000 1.000 ;
 END
 ANTENNAPARTIALMETALAREA                  3.146 LAYER ME2 ;
 ANTENNAGATEAREA                          0.086 LAYER ME2 ;
 ANTENNAGATEAREA                          0.086 LAYER ME3 ;
 ANTENNAGATEAREA                          0.086 LAYER ME4 ;
 ANTENNADIFFAREA                          0.160 LAYER ME2 ;
 ANTENNADIFFAREA                          0.160 LAYER ME3 ;
 ANTENNADIFFAREA                          0.160 LAYER ME4 ;
 ANTENNAMAXAREACAR                       48.755 LAYER ME2 ;
 ANTENNAMAXAREACAR                       58.014 LAYER ME3 ;
 ANTENNAMAXAREACAR                       67.273 LAYER ME4 ;
END DI25
PIN DO24
  DIRECTION OUTPUT ;
 PORT
  LAYER ME4 ;
  RECT 514.000 0.000 514.800 1.000 ;
  LAYER ME3 ;
  RECT 514.000 0.000 514.800 1.000 ;
  LAYER ME2 ;
  RECT 514.000 0.000 514.800 1.000 ;
  LAYER ME1 ;
  RECT 514.000 0.000 514.800 1.000 ;
 END
 ANTENNAPARTIALMETALAREA                  4.172 LAYER ME2 ;
 ANTENNADIFFAREA                          5.472 LAYER ME2 ;
 ANTENNADIFFAREA                          5.472 LAYER ME3 ;
 ANTENNADIFFAREA                          5.472 LAYER ME4 ;
END DO24
PIN DI24
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 499.200 0.000 500.000 1.000 ;
  LAYER ME3 ;
  RECT 499.200 0.000 500.000 1.000 ;
  LAYER ME2 ;
  RECT 499.200 0.000 500.000 1.000 ;
  LAYER ME1 ;
  RECT 499.200 0.000 500.000 1.000 ;
 END
 ANTENNAPARTIALMETALAREA                  3.118 LAYER ME2 ;
 ANTENNAGATEAREA                          0.086 LAYER ME2 ;
 ANTENNAGATEAREA                          0.086 LAYER ME3 ;
 ANTENNAGATEAREA                          0.086 LAYER ME4 ;
 ANTENNADIFFAREA                          0.160 LAYER ME2 ;
 ANTENNADIFFAREA                          0.160 LAYER ME3 ;
 ANTENNADIFFAREA                          0.160 LAYER ME4 ;
 ANTENNAMAXAREACAR                       48.431 LAYER ME2 ;
 ANTENNAMAXAREACAR                       57.690 LAYER ME3 ;
 ANTENNAMAXAREACAR                       66.949 LAYER ME4 ;
END DI24
PIN DO23
  DIRECTION OUTPUT ;
 PORT
  LAYER ME4 ;
  RECT 492.800 0.000 493.600 1.000 ;
  LAYER ME3 ;
  RECT 492.800 0.000 493.600 1.000 ;
  LAYER ME2 ;
  RECT 492.800 0.000 493.600 1.000 ;
  LAYER ME1 ;
  RECT 492.800 0.000 493.600 1.000 ;
 END
 ANTENNAPARTIALMETALAREA                  4.148 LAYER ME2 ;
 ANTENNADIFFAREA                          5.472 LAYER ME2 ;
 ANTENNADIFFAREA                          5.472 LAYER ME3 ;
 ANTENNADIFFAREA                          5.472 LAYER ME4 ;
END DO23
PIN DI23
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 478.000 0.000 478.800 1.000 ;
  LAYER ME3 ;
  RECT 478.000 0.000 478.800 1.000 ;
  LAYER ME2 ;
  RECT 478.000 0.000 478.800 1.000 ;
  LAYER ME1 ;
  RECT 478.000 0.000 478.800 1.000 ;
 END
 ANTENNAPARTIALMETALAREA                  3.142 LAYER ME2 ;
 ANTENNAGATEAREA                          0.086 LAYER ME2 ;
 ANTENNAGATEAREA                          0.086 LAYER ME3 ;
 ANTENNAGATEAREA                          0.086 LAYER ME4 ;
 ANTENNADIFFAREA                          0.160 LAYER ME2 ;
 ANTENNADIFFAREA                          0.160 LAYER ME3 ;
 ANTENNADIFFAREA                          0.160 LAYER ME4 ;
 ANTENNAMAXAREACAR                       48.708 LAYER ME2 ;
 ANTENNAMAXAREACAR                       57.968 LAYER ME3 ;
 ANTENNAMAXAREACAR                       67.227 LAYER ME4 ;
END DI23
PIN DO22
  DIRECTION OUTPUT ;
 PORT
  LAYER ME4 ;
  RECT 472.800 0.000 473.600 1.000 ;
  LAYER ME3 ;
  RECT 472.800 0.000 473.600 1.000 ;
  LAYER ME2 ;
  RECT 472.800 0.000 473.600 1.000 ;
  LAYER ME1 ;
  RECT 472.800 0.000 473.600 1.000 ;
 END
 ANTENNAPARTIALMETALAREA                  4.164 LAYER ME2 ;
 ANTENNADIFFAREA                          5.472 LAYER ME2 ;
 ANTENNADIFFAREA                          5.472 LAYER ME3 ;
 ANTENNADIFFAREA                          5.472 LAYER ME4 ;
END DO22
PIN DI22
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 458.400 0.000 459.200 1.000 ;
  LAYER ME3 ;
  RECT 458.400 0.000 459.200 1.000 ;
  LAYER ME2 ;
  RECT 458.400 0.000 459.200 1.000 ;
  LAYER ME1 ;
  RECT 458.400 0.000 459.200 1.000 ;
 END
 ANTENNAPARTIALMETALAREA                  3.138 LAYER ME2 ;
 ANTENNAGATEAREA                          0.086 LAYER ME2 ;
 ANTENNAGATEAREA                          0.086 LAYER ME3 ;
 ANTENNAGATEAREA                          0.086 LAYER ME4 ;
 ANTENNADIFFAREA                          0.160 LAYER ME2 ;
 ANTENNADIFFAREA                          0.160 LAYER ME3 ;
 ANTENNADIFFAREA                          0.160 LAYER ME4 ;
 ANTENNAMAXAREACAR                       48.662 LAYER ME2 ;
 ANTENNAMAXAREACAR                       57.921 LAYER ME3 ;
 ANTENNAMAXAREACAR                       67.181 LAYER ME4 ;
END DI22
PIN DO21
  DIRECTION OUTPUT ;
 PORT
  LAYER ME4 ;
  RECT 452.000 0.000 452.800 1.000 ;
  LAYER ME3 ;
  RECT 452.000 0.000 452.800 1.000 ;
  LAYER ME2 ;
  RECT 452.000 0.000 452.800 1.000 ;
  LAYER ME1 ;
  RECT 452.000 0.000 452.800 1.000 ;
 END
 ANTENNAPARTIALMETALAREA                  4.172 LAYER ME2 ;
 ANTENNADIFFAREA                          5.472 LAYER ME2 ;
 ANTENNADIFFAREA                          5.472 LAYER ME3 ;
 ANTENNADIFFAREA                          5.472 LAYER ME4 ;
END DO21
PIN DI21
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 437.200 0.000 438.000 1.000 ;
  LAYER ME3 ;
  RECT 437.200 0.000 438.000 1.000 ;
  LAYER ME2 ;
  RECT 437.200 0.000 438.000 1.000 ;
  LAYER ME1 ;
  RECT 437.200 0.000 438.000 1.000 ;
 END
 ANTENNAPARTIALMETALAREA                  3.118 LAYER ME2 ;
 ANTENNAGATEAREA                          0.086 LAYER ME2 ;
 ANTENNAGATEAREA                          0.086 LAYER ME3 ;
 ANTENNAGATEAREA                          0.086 LAYER ME4 ;
 ANTENNADIFFAREA                          0.160 LAYER ME2 ;
 ANTENNADIFFAREA                          0.160 LAYER ME3 ;
 ANTENNADIFFAREA                          0.160 LAYER ME4 ;
 ANTENNAMAXAREACAR                       48.431 LAYER ME2 ;
 ANTENNAMAXAREACAR                       57.690 LAYER ME3 ;
 ANTENNAMAXAREACAR                       66.949 LAYER ME4 ;
END DI21
PIN DO20
  DIRECTION OUTPUT ;
 PORT
  LAYER ME4 ;
  RECT 432.000 0.000 432.800 1.000 ;
  LAYER ME3 ;
  RECT 432.000 0.000 432.800 1.000 ;
  LAYER ME2 ;
  RECT 432.000 0.000 432.800 1.000 ;
  LAYER ME1 ;
  RECT 432.000 0.000 432.800 1.000 ;
 END
 ANTENNAPARTIALMETALAREA                  4.140 LAYER ME2 ;
 ANTENNADIFFAREA                          5.472 LAYER ME2 ;
 ANTENNADIFFAREA                          5.472 LAYER ME3 ;
 ANTENNADIFFAREA                          5.472 LAYER ME4 ;
END DO20
PIN DI20
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 417.200 0.000 418.000 1.000 ;
  LAYER ME3 ;
  RECT 417.200 0.000 418.000 1.000 ;
  LAYER ME2 ;
  RECT 417.200 0.000 418.000 1.000 ;
  LAYER ME1 ;
  RECT 417.200 0.000 418.000 1.000 ;
 END
 ANTENNAPARTIALMETALAREA                  3.150 LAYER ME2 ;
 ANTENNAGATEAREA                          0.086 LAYER ME2 ;
 ANTENNAGATEAREA                          0.086 LAYER ME3 ;
 ANTENNAGATEAREA                          0.086 LAYER ME4 ;
 ANTENNADIFFAREA                          0.160 LAYER ME2 ;
 ANTENNADIFFAREA                          0.160 LAYER ME3 ;
 ANTENNADIFFAREA                          0.160 LAYER ME4 ;
 ANTENNAMAXAREACAR                       48.801 LAYER ME2 ;
 ANTENNAMAXAREACAR                       58.060 LAYER ME3 ;
 ANTENNAMAXAREACAR                       67.319 LAYER ME4 ;
END DI20
PIN DO19
  DIRECTION OUTPUT ;
 PORT
  LAYER ME4 ;
  RECT 410.800 0.000 411.600 1.000 ;
  LAYER ME3 ;
  RECT 410.800 0.000 411.600 1.000 ;
  LAYER ME2 ;
  RECT 410.800 0.000 411.600 1.000 ;
  LAYER ME1 ;
  RECT 410.800 0.000 411.600 1.000 ;
 END
 ANTENNAPARTIALMETALAREA                  4.164 LAYER ME2 ;
 ANTENNADIFFAREA                          5.472 LAYER ME2 ;
 ANTENNADIFFAREA                          5.472 LAYER ME3 ;
 ANTENNADIFFAREA                          5.472 LAYER ME4 ;
END DO19
PIN DI19
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 396.400 0.000 397.200 1.000 ;
  LAYER ME3 ;
  RECT 396.400 0.000 397.200 1.000 ;
  LAYER ME2 ;
  RECT 396.400 0.000 397.200 1.000 ;
  LAYER ME1 ;
  RECT 396.400 0.000 397.200 1.000 ;
 END
 ANTENNAPARTIALMETALAREA                  3.138 LAYER ME2 ;
 ANTENNAGATEAREA                          0.086 LAYER ME2 ;
 ANTENNAGATEAREA                          0.086 LAYER ME3 ;
 ANTENNAGATEAREA                          0.086 LAYER ME4 ;
 ANTENNADIFFAREA                          0.160 LAYER ME2 ;
 ANTENNADIFFAREA                          0.160 LAYER ME3 ;
 ANTENNADIFFAREA                          0.160 LAYER ME4 ;
 ANTENNAMAXAREACAR                       48.662 LAYER ME2 ;
 ANTENNAMAXAREACAR                       57.921 LAYER ME3 ;
 ANTENNAMAXAREACAR                       67.181 LAYER ME4 ;
END DI19
PIN DO18
  DIRECTION OUTPUT ;
 PORT
  LAYER ME4 ;
  RECT 391.200 0.000 392.000 1.000 ;
  LAYER ME3 ;
  RECT 391.200 0.000 392.000 1.000 ;
  LAYER ME2 ;
  RECT 391.200 0.000 392.000 1.000 ;
  LAYER ME1 ;
  RECT 391.200 0.000 392.000 1.000 ;
 END
 ANTENNAPARTIALMETALAREA                  4.164 LAYER ME2 ;
 ANTENNADIFFAREA                          5.472 LAYER ME2 ;
 ANTENNADIFFAREA                          5.472 LAYER ME3 ;
 ANTENNADIFFAREA                          5.472 LAYER ME4 ;
END DO18
PIN DI18
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 376.400 0.000 377.200 1.000 ;
  LAYER ME3 ;
  RECT 376.400 0.000 377.200 1.000 ;
  LAYER ME2 ;
  RECT 376.400 0.000 377.200 1.000 ;
  LAYER ME1 ;
  RECT 376.400 0.000 377.200 1.000 ;
 END
 ANTENNAPARTIALMETALAREA                  3.126 LAYER ME2 ;
 ANTENNAGATEAREA                          0.086 LAYER ME2 ;
 ANTENNAGATEAREA                          0.086 LAYER ME3 ;
 ANTENNAGATEAREA                          0.086 LAYER ME4 ;
 ANTENNADIFFAREA                          0.160 LAYER ME2 ;
 ANTENNADIFFAREA                          0.160 LAYER ME3 ;
 ANTENNADIFFAREA                          0.160 LAYER ME4 ;
 ANTENNAMAXAREACAR                       48.523 LAYER ME2 ;
 ANTENNAMAXAREACAR                       57.782 LAYER ME3 ;
 ANTENNAMAXAREACAR                       67.042 LAYER ME4 ;
END DI18
PIN DO17
  DIRECTION OUTPUT ;
 PORT
  LAYER ME4 ;
  RECT 370.000 0.000 370.800 1.000 ;
  LAYER ME3 ;
  RECT 370.000 0.000 370.800 1.000 ;
  LAYER ME2 ;
  RECT 370.000 0.000 370.800 1.000 ;
  LAYER ME1 ;
  RECT 370.000 0.000 370.800 1.000 ;
 END
 ANTENNAPARTIALMETALAREA                  4.140 LAYER ME2 ;
 ANTENNADIFFAREA                          5.472 LAYER ME2 ;
 ANTENNADIFFAREA                          5.472 LAYER ME3 ;
 ANTENNADIFFAREA                          5.472 LAYER ME4 ;
END DO17
PIN DI17
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 355.200 0.000 356.000 1.000 ;
  LAYER ME3 ;
  RECT 355.200 0.000 356.000 1.000 ;
  LAYER ME2 ;
  RECT 355.200 0.000 356.000 1.000 ;
  LAYER ME1 ;
  RECT 355.200 0.000 356.000 1.000 ;
 END
 ANTENNAPARTIALMETALAREA                  3.150 LAYER ME2 ;
 ANTENNAGATEAREA                          0.086 LAYER ME2 ;
 ANTENNAGATEAREA                          0.086 LAYER ME3 ;
 ANTENNAGATEAREA                          0.086 LAYER ME4 ;
 ANTENNADIFFAREA                          0.160 LAYER ME2 ;
 ANTENNADIFFAREA                          0.160 LAYER ME3 ;
 ANTENNADIFFAREA                          0.160 LAYER ME4 ;
 ANTENNAMAXAREACAR                       48.801 LAYER ME2 ;
 ANTENNAMAXAREACAR                       58.060 LAYER ME3 ;
 ANTENNAMAXAREACAR                       67.319 LAYER ME4 ;
END DI17
PIN DO16
  DIRECTION OUTPUT ;
 PORT
  LAYER ME4 ;
  RECT 350.000 0.000 350.800 1.000 ;
  LAYER ME3 ;
  RECT 350.000 0.000 350.800 1.000 ;
  LAYER ME2 ;
  RECT 350.000 0.000 350.800 1.000 ;
  LAYER ME1 ;
  RECT 350.000 0.000 350.800 1.000 ;
 END
 ANTENNAPARTIALMETALAREA                  4.172 LAYER ME2 ;
 ANTENNADIFFAREA                          5.472 LAYER ME2 ;
 ANTENNADIFFAREA                          5.472 LAYER ME3 ;
 ANTENNADIFFAREA                          5.472 LAYER ME4 ;
END DO16
PIN WEB1
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 337.200 0.000 338.000 1.000 ;
  LAYER ME3 ;
  RECT 337.200 0.000 338.000 1.000 ;
  LAYER ME2 ;
  RECT 337.200 0.000 338.000 1.000 ;
  LAYER ME1 ;
  RECT 337.200 0.000 338.000 1.000 ;
 END
 ANTENNAPARTIALMETALAREA                  2.840 LAYER ME2 ;
 ANTENNAGATEAREA                          0.072 LAYER ME2 ;
 ANTENNAGATEAREA                          0.072 LAYER ME3 ;
 ANTENNAGATEAREA                          0.072 LAYER ME4 ;
 ANTENNADIFFAREA                          0.160 LAYER ME2 ;
 ANTENNADIFFAREA                          0.160 LAYER ME3 ;
 ANTENNADIFFAREA                          0.160 LAYER ME4 ;
 ANTENNAMAXAREACAR                       54.456 LAYER ME2 ;
 ANTENNAMAXAREACAR                       65.567 LAYER ME3 ;
 ANTENNAMAXAREACAR                       76.678 LAYER ME4 ;
END WEB1
PIN DI16
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 335.600 0.000 336.400 1.000 ;
  LAYER ME3 ;
  RECT 335.600 0.000 336.400 1.000 ;
  LAYER ME2 ;
  RECT 335.600 0.000 336.400 1.000 ;
  LAYER ME1 ;
  RECT 335.600 0.000 336.400 1.000 ;
 END
 ANTENNAPARTIALMETALAREA                  3.130 LAYER ME2 ;
 ANTENNAGATEAREA                          0.086 LAYER ME2 ;
 ANTENNAGATEAREA                          0.086 LAYER ME3 ;
 ANTENNAGATEAREA                          0.086 LAYER ME4 ;
 ANTENNADIFFAREA                          0.160 LAYER ME2 ;
 ANTENNADIFFAREA                          0.160 LAYER ME3 ;
 ANTENNADIFFAREA                          0.160 LAYER ME4 ;
 ANTENNAMAXAREACAR                       48.569 LAYER ME2 ;
 ANTENNAMAXAREACAR                       57.829 LAYER ME3 ;
 ANTENNAMAXAREACAR                       67.088 LAYER ME4 ;
END DI16
PIN DO15
  DIRECTION OUTPUT ;
 PORT
  LAYER ME4 ;
  RECT 329.200 0.000 330.000 1.000 ;
  LAYER ME3 ;
  RECT 329.200 0.000 330.000 1.000 ;
  LAYER ME2 ;
  RECT 329.200 0.000 330.000 1.000 ;
  LAYER ME1 ;
  RECT 329.200 0.000 330.000 1.000 ;
 END
 ANTENNAPARTIALMETALAREA                  4.164 LAYER ME2 ;
 ANTENNADIFFAREA                          5.472 LAYER ME2 ;
 ANTENNADIFFAREA                          5.472 LAYER ME3 ;
 ANTENNADIFFAREA                          5.472 LAYER ME4 ;
END DO15
PIN DI15
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 314.400 0.000 315.200 1.000 ;
  LAYER ME3 ;
  RECT 314.400 0.000 315.200 1.000 ;
  LAYER ME2 ;
  RECT 314.400 0.000 315.200 1.000 ;
  LAYER ME1 ;
  RECT 314.400 0.000 315.200 1.000 ;
 END
 ANTENNAPARTIALMETALAREA                  3.126 LAYER ME2 ;
 ANTENNAGATEAREA                          0.086 LAYER ME2 ;
 ANTENNAGATEAREA                          0.086 LAYER ME3 ;
 ANTENNAGATEAREA                          0.086 LAYER ME4 ;
 ANTENNADIFFAREA                          0.160 LAYER ME2 ;
 ANTENNADIFFAREA                          0.160 LAYER ME3 ;
 ANTENNADIFFAREA                          0.160 LAYER ME4 ;
 ANTENNAMAXAREACAR                       48.523 LAYER ME2 ;
 ANTENNAMAXAREACAR                       57.782 LAYER ME3 ;
 ANTENNAMAXAREACAR                       67.042 LAYER ME4 ;
END DI15
PIN DO14
  DIRECTION OUTPUT ;
 PORT
  LAYER ME4 ;
  RECT 309.200 0.000 310.000 1.000 ;
  LAYER ME3 ;
  RECT 309.200 0.000 310.000 1.000 ;
  LAYER ME2 ;
  RECT 309.200 0.000 310.000 1.000 ;
  LAYER ME1 ;
  RECT 309.200 0.000 310.000 1.000 ;
 END
 ANTENNAPARTIALMETALAREA                  4.148 LAYER ME2 ;
 ANTENNADIFFAREA                          5.472 LAYER ME2 ;
 ANTENNADIFFAREA                          5.472 LAYER ME3 ;
 ANTENNADIFFAREA                          5.472 LAYER ME4 ;
END DO14
PIN DI14
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 294.800 0.000 295.600 1.000 ;
  LAYER ME3 ;
  RECT 294.800 0.000 295.600 1.000 ;
  LAYER ME2 ;
  RECT 294.800 0.000 295.600 1.000 ;
  LAYER ME1 ;
  RECT 294.800 0.000 295.600 1.000 ;
 END
 ANTENNAPARTIALMETALAREA                  3.154 LAYER ME2 ;
 ANTENNAGATEAREA                          0.086 LAYER ME2 ;
 ANTENNAGATEAREA                          0.086 LAYER ME3 ;
 ANTENNAGATEAREA                          0.086 LAYER ME4 ;
 ANTENNADIFFAREA                          0.160 LAYER ME2 ;
 ANTENNADIFFAREA                          0.160 LAYER ME3 ;
 ANTENNADIFFAREA                          0.160 LAYER ME4 ;
 ANTENNAMAXAREACAR                       48.847 LAYER ME2 ;
 ANTENNAMAXAREACAR                       58.106 LAYER ME3 ;
 ANTENNAMAXAREACAR                       67.366 LAYER ME4 ;
END DI14
PIN DO13
  DIRECTION OUTPUT ;
 PORT
  LAYER ME4 ;
  RECT 288.000 0.000 288.800 1.000 ;
  LAYER ME3 ;
  RECT 288.000 0.000 288.800 1.000 ;
  LAYER ME2 ;
  RECT 288.000 0.000 288.800 1.000 ;
  LAYER ME1 ;
  RECT 288.000 0.000 288.800 1.000 ;
 END
 ANTENNAPARTIALMETALAREA                  4.172 LAYER ME2 ;
 ANTENNADIFFAREA                          5.472 LAYER ME2 ;
 ANTENNADIFFAREA                          5.472 LAYER ME3 ;
 ANTENNADIFFAREA                          5.472 LAYER ME4 ;
END DO13
PIN DI13
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 273.600 0.000 274.400 1.000 ;
  LAYER ME3 ;
  RECT 273.600 0.000 274.400 1.000 ;
  LAYER ME2 ;
  RECT 273.600 0.000 274.400 1.000 ;
  LAYER ME1 ;
  RECT 273.600 0.000 274.400 1.000 ;
 END
 ANTENNAPARTIALMETALAREA                  3.130 LAYER ME2 ;
 ANTENNAGATEAREA                          0.086 LAYER ME2 ;
 ANTENNAGATEAREA                          0.086 LAYER ME3 ;
 ANTENNAGATEAREA                          0.086 LAYER ME4 ;
 ANTENNADIFFAREA                          0.160 LAYER ME2 ;
 ANTENNADIFFAREA                          0.160 LAYER ME3 ;
 ANTENNADIFFAREA                          0.160 LAYER ME4 ;
 ANTENNAMAXAREACAR                       48.569 LAYER ME2 ;
 ANTENNAMAXAREACAR                       57.829 LAYER ME3 ;
 ANTENNAMAXAREACAR                       67.088 LAYER ME4 ;
END DI13
PIN DO12
  DIRECTION OUTPUT ;
 PORT
  LAYER ME4 ;
  RECT 268.400 0.000 269.200 1.000 ;
  LAYER ME3 ;
  RECT 268.400 0.000 269.200 1.000 ;
  LAYER ME2 ;
  RECT 268.400 0.000 269.200 1.000 ;
  LAYER ME1 ;
  RECT 268.400 0.000 269.200 1.000 ;
 END
 ANTENNAPARTIALMETALAREA                  4.156 LAYER ME2 ;
 ANTENNADIFFAREA                          5.472 LAYER ME2 ;
 ANTENNADIFFAREA                          5.472 LAYER ME3 ;
 ANTENNADIFFAREA                          5.472 LAYER ME4 ;
END DO12
PIN DI12
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 253.600 0.000 254.400 1.000 ;
  LAYER ME3 ;
  RECT 253.600 0.000 254.400 1.000 ;
  LAYER ME2 ;
  RECT 253.600 0.000 254.400 1.000 ;
  LAYER ME1 ;
  RECT 253.600 0.000 254.400 1.000 ;
 END
 ANTENNAPARTIALMETALAREA                  3.134 LAYER ME2 ;
 ANTENNAGATEAREA                          0.086 LAYER ME2 ;
 ANTENNAGATEAREA                          0.086 LAYER ME3 ;
 ANTENNAGATEAREA                          0.086 LAYER ME4 ;
 ANTENNADIFFAREA                          0.160 LAYER ME2 ;
 ANTENNADIFFAREA                          0.160 LAYER ME3 ;
 ANTENNADIFFAREA                          0.160 LAYER ME4 ;
 ANTENNAMAXAREACAR                       48.616 LAYER ME2 ;
 ANTENNAMAXAREACAR                       57.875 LAYER ME3 ;
 ANTENNAMAXAREACAR                       67.134 LAYER ME4 ;
END DI12
PIN DO11
  DIRECTION OUTPUT ;
 PORT
  LAYER ME4 ;
  RECT 247.200 0.000 248.000 1.000 ;
  LAYER ME3 ;
  RECT 247.200 0.000 248.000 1.000 ;
  LAYER ME2 ;
  RECT 247.200 0.000 248.000 1.000 ;
  LAYER ME1 ;
  RECT 247.200 0.000 248.000 1.000 ;
 END
 ANTENNAPARTIALMETALAREA                  4.148 LAYER ME2 ;
 ANTENNADIFFAREA                          5.472 LAYER ME2 ;
 ANTENNADIFFAREA                          5.472 LAYER ME3 ;
 ANTENNADIFFAREA                          5.472 LAYER ME4 ;
END DO11
PIN DI11
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 232.800 0.000 233.600 1.000 ;
  LAYER ME3 ;
  RECT 232.800 0.000 233.600 1.000 ;
  LAYER ME2 ;
  RECT 232.800 0.000 233.600 1.000 ;
  LAYER ME1 ;
  RECT 232.800 0.000 233.600 1.000 ;
 END
 ANTENNAPARTIALMETALAREA                  3.154 LAYER ME2 ;
 ANTENNAGATEAREA                          0.086 LAYER ME2 ;
 ANTENNAGATEAREA                          0.086 LAYER ME3 ;
 ANTENNAGATEAREA                          0.086 LAYER ME4 ;
 ANTENNADIFFAREA                          0.160 LAYER ME2 ;
 ANTENNADIFFAREA                          0.160 LAYER ME3 ;
 ANTENNADIFFAREA                          0.160 LAYER ME4 ;
 ANTENNAMAXAREACAR                       48.847 LAYER ME2 ;
 ANTENNAMAXAREACAR                       58.106 LAYER ME3 ;
 ANTENNAMAXAREACAR                       67.366 LAYER ME4 ;
END DI11
PIN DO10
  DIRECTION OUTPUT ;
 PORT
  LAYER ME4 ;
  RECT 227.200 0.000 228.000 1.000 ;
  LAYER ME3 ;
  RECT 227.200 0.000 228.000 1.000 ;
  LAYER ME2 ;
  RECT 227.200 0.000 228.000 1.000 ;
  LAYER ME1 ;
  RECT 227.200 0.000 228.000 1.000 ;
 END
 ANTENNAPARTIALMETALAREA                  4.180 LAYER ME2 ;
 ANTENNADIFFAREA                          5.472 LAYER ME2 ;
 ANTENNADIFFAREA                          5.472 LAYER ME3 ;
 ANTENNADIFFAREA                          5.472 LAYER ME4 ;
END DO10
PIN DI10
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 212.800 0.000 213.600 1.000 ;
  LAYER ME3 ;
  RECT 212.800 0.000 213.600 1.000 ;
  LAYER ME2 ;
  RECT 212.800 0.000 213.600 1.000 ;
  LAYER ME1 ;
  RECT 212.800 0.000 213.600 1.000 ;
 END
 ANTENNAPARTIALMETALAREA                  3.122 LAYER ME2 ;
 ANTENNAGATEAREA                          0.086 LAYER ME2 ;
 ANTENNAGATEAREA                          0.086 LAYER ME3 ;
 ANTENNAGATEAREA                          0.086 LAYER ME4 ;
 ANTENNADIFFAREA                          0.160 LAYER ME2 ;
 ANTENNADIFFAREA                          0.160 LAYER ME3 ;
 ANTENNADIFFAREA                          0.160 LAYER ME4 ;
 ANTENNAMAXAREACAR                       48.477 LAYER ME2 ;
 ANTENNAMAXAREACAR                       57.736 LAYER ME3 ;
 ANTENNAMAXAREACAR                       66.995 LAYER ME4 ;
END DI10
PIN DO9
  DIRECTION OUTPUT ;
 PORT
  LAYER ME4 ;
  RECT 206.400 0.000 207.200 1.000 ;
  LAYER ME3 ;
  RECT 206.400 0.000 207.200 1.000 ;
  LAYER ME2 ;
  RECT 206.400 0.000 207.200 1.000 ;
  LAYER ME1 ;
  RECT 206.400 0.000 207.200 1.000 ;
 END
 ANTENNAPARTIALMETALAREA                  4.156 LAYER ME2 ;
 ANTENNADIFFAREA                          5.472 LAYER ME2 ;
 ANTENNADIFFAREA                          5.472 LAYER ME3 ;
 ANTENNADIFFAREA                          5.472 LAYER ME4 ;
END DO9
PIN DI9
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 191.600 0.000 192.400 1.000 ;
  LAYER ME3 ;
  RECT 191.600 0.000 192.400 1.000 ;
  LAYER ME2 ;
  RECT 191.600 0.000 192.400 1.000 ;
  LAYER ME1 ;
  RECT 191.600 0.000 192.400 1.000 ;
 END
 ANTENNAPARTIALMETALAREA                  3.134 LAYER ME2 ;
 ANTENNAGATEAREA                          0.086 LAYER ME2 ;
 ANTENNAGATEAREA                          0.086 LAYER ME3 ;
 ANTENNAGATEAREA                          0.086 LAYER ME4 ;
 ANTENNADIFFAREA                          0.160 LAYER ME2 ;
 ANTENNADIFFAREA                          0.160 LAYER ME3 ;
 ANTENNADIFFAREA                          0.160 LAYER ME4 ;
 ANTENNAMAXAREACAR                       48.616 LAYER ME2 ;
 ANTENNAMAXAREACAR                       57.875 LAYER ME3 ;
 ANTENNAMAXAREACAR                       67.134 LAYER ME4 ;
END DI9
PIN DO8
  DIRECTION OUTPUT ;
 PORT
  LAYER ME4 ;
  RECT 186.400 0.000 187.200 1.000 ;
  LAYER ME3 ;
  RECT 186.400 0.000 187.200 1.000 ;
  LAYER ME2 ;
  RECT 186.400 0.000 187.200 1.000 ;
  LAYER ME1 ;
  RECT 186.400 0.000 187.200 1.000 ;
 END
 ANTENNAPARTIALMETALAREA                  4.156 LAYER ME2 ;
 ANTENNADIFFAREA                          5.472 LAYER ME2 ;
 ANTENNADIFFAREA                          5.472 LAYER ME3 ;
 ANTENNADIFFAREA                          5.472 LAYER ME4 ;
END DO8
PIN DI8
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 172.000 0.000 172.800 1.000 ;
  LAYER ME3 ;
  RECT 172.000 0.000 172.800 1.000 ;
  LAYER ME2 ;
  RECT 172.000 0.000 172.800 1.000 ;
  LAYER ME1 ;
  RECT 172.000 0.000 172.800 1.000 ;
 END
 ANTENNAPARTIALMETALAREA                  3.146 LAYER ME2 ;
 ANTENNAGATEAREA                          0.086 LAYER ME2 ;
 ANTENNAGATEAREA                          0.086 LAYER ME3 ;
 ANTENNAGATEAREA                          0.086 LAYER ME4 ;
 ANTENNADIFFAREA                          0.160 LAYER ME2 ;
 ANTENNADIFFAREA                          0.160 LAYER ME3 ;
 ANTENNADIFFAREA                          0.160 LAYER ME4 ;
 ANTENNAMAXAREACAR                       48.755 LAYER ME2 ;
 ANTENNAMAXAREACAR                       58.014 LAYER ME3 ;
 ANTENNAMAXAREACAR                       67.273 LAYER ME4 ;
END DI8
PIN DO7
  DIRECTION OUTPUT ;
 PORT
  LAYER ME4 ;
  RECT 165.200 0.000 166.000 1.000 ;
  LAYER ME3 ;
  RECT 165.200 0.000 166.000 1.000 ;
  LAYER ME2 ;
  RECT 165.200 0.000 166.000 1.000 ;
  LAYER ME1 ;
  RECT 165.200 0.000 166.000 1.000 ;
 END
 ANTENNAPARTIALMETALAREA                  4.180 LAYER ME2 ;
 ANTENNADIFFAREA                          5.472 LAYER ME2 ;
 ANTENNADIFFAREA                          5.472 LAYER ME3 ;
 ANTENNADIFFAREA                          5.472 LAYER ME4 ;
END DO7
PIN DI7
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 150.800 0.000 151.600 1.000 ;
  LAYER ME3 ;
  RECT 150.800 0.000 151.600 1.000 ;
  LAYER ME2 ;
  RECT 150.800 0.000 151.600 1.000 ;
  LAYER ME1 ;
  RECT 150.800 0.000 151.600 1.000 ;
 END
 ANTENNAPARTIALMETALAREA                  3.122 LAYER ME2 ;
 ANTENNAGATEAREA                          0.086 LAYER ME2 ;
 ANTENNAGATEAREA                          0.086 LAYER ME3 ;
 ANTENNAGATEAREA                          0.086 LAYER ME4 ;
 ANTENNADIFFAREA                          0.160 LAYER ME2 ;
 ANTENNADIFFAREA                          0.160 LAYER ME3 ;
 ANTENNADIFFAREA                          0.160 LAYER ME4 ;
 ANTENNAMAXAREACAR                       48.477 LAYER ME2 ;
 ANTENNAMAXAREACAR                       57.736 LAYER ME3 ;
 ANTENNAMAXAREACAR                       66.995 LAYER ME4 ;
END DI7
PIN DO6
  DIRECTION OUTPUT ;
 PORT
  LAYER ME4 ;
  RECT 145.600 0.000 146.400 1.000 ;
  LAYER ME3 ;
  RECT 145.600 0.000 146.400 1.000 ;
  LAYER ME2 ;
  RECT 145.600 0.000 146.400 1.000 ;
  LAYER ME1 ;
  RECT 145.600 0.000 146.400 1.000 ;
 END
 ANTENNAPARTIALMETALAREA                  4.148 LAYER ME2 ;
 ANTENNADIFFAREA                          5.472 LAYER ME2 ;
 ANTENNADIFFAREA                          5.472 LAYER ME3 ;
 ANTENNADIFFAREA                          5.472 LAYER ME4 ;
END DO6
PIN DI6
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 130.800 0.000 131.600 1.000 ;
  LAYER ME3 ;
  RECT 130.800 0.000 131.600 1.000 ;
  LAYER ME2 ;
  RECT 130.800 0.000 131.600 1.000 ;
  LAYER ME1 ;
  RECT 130.800 0.000 131.600 1.000 ;
 END
 ANTENNAPARTIALMETALAREA                  3.142 LAYER ME2 ;
 ANTENNAGATEAREA                          0.086 LAYER ME2 ;
 ANTENNAGATEAREA                          0.086 LAYER ME3 ;
 ANTENNAGATEAREA                          0.086 LAYER ME4 ;
 ANTENNADIFFAREA                          0.160 LAYER ME2 ;
 ANTENNADIFFAREA                          0.160 LAYER ME3 ;
 ANTENNADIFFAREA                          0.160 LAYER ME4 ;
 ANTENNAMAXAREACAR                       48.708 LAYER ME2 ;
 ANTENNAMAXAREACAR                       57.968 LAYER ME3 ;
 ANTENNAMAXAREACAR                       67.227 LAYER ME4 ;
END DI6
PIN DO5
  DIRECTION OUTPUT ;
 PORT
  LAYER ME4 ;
  RECT 124.400 0.000 125.200 1.000 ;
  LAYER ME3 ;
  RECT 124.400 0.000 125.200 1.000 ;
  LAYER ME2 ;
  RECT 124.400 0.000 125.200 1.000 ;
  LAYER ME1 ;
  RECT 124.400 0.000 125.200 1.000 ;
 END
 ANTENNAPARTIALMETALAREA                  4.156 LAYER ME2 ;
 ANTENNADIFFAREA                          5.472 LAYER ME2 ;
 ANTENNADIFFAREA                          5.472 LAYER ME3 ;
 ANTENNADIFFAREA                          5.472 LAYER ME4 ;
END DO5
PIN DI5
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 110.000 0.000 110.800 1.000 ;
  LAYER ME3 ;
  RECT 110.000 0.000 110.800 1.000 ;
  LAYER ME2 ;
  RECT 110.000 0.000 110.800 1.000 ;
  LAYER ME1 ;
  RECT 110.000 0.000 110.800 1.000 ;
 END
 ANTENNAPARTIALMETALAREA                  3.146 LAYER ME2 ;
 ANTENNAGATEAREA                          0.086 LAYER ME2 ;
 ANTENNAGATEAREA                          0.086 LAYER ME3 ;
 ANTENNAGATEAREA                          0.086 LAYER ME4 ;
 ANTENNADIFFAREA                          0.160 LAYER ME2 ;
 ANTENNADIFFAREA                          0.160 LAYER ME3 ;
 ANTENNADIFFAREA                          0.160 LAYER ME4 ;
 ANTENNAMAXAREACAR                       48.755 LAYER ME2 ;
 ANTENNAMAXAREACAR                       58.014 LAYER ME3 ;
 ANTENNAMAXAREACAR                       67.273 LAYER ME4 ;
END DI5
PIN DO4
  DIRECTION OUTPUT ;
 PORT
  LAYER ME4 ;
  RECT 104.800 0.000 105.600 1.000 ;
  LAYER ME3 ;
  RECT 104.800 0.000 105.600 1.000 ;
  LAYER ME2 ;
  RECT 104.800 0.000 105.600 1.000 ;
  LAYER ME1 ;
  RECT 104.800 0.000 105.600 1.000 ;
 END
 ANTENNAPARTIALMETALAREA                  4.172 LAYER ME2 ;
 ANTENNADIFFAREA                          5.472 LAYER ME2 ;
 ANTENNADIFFAREA                          5.472 LAYER ME3 ;
 ANTENNADIFFAREA                          5.472 LAYER ME4 ;
END DO4
PIN DI4
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 90.000 0.000 90.800 1.000 ;
  LAYER ME3 ;
  RECT 90.000 0.000 90.800 1.000 ;
  LAYER ME2 ;
  RECT 90.000 0.000 90.800 1.000 ;
  LAYER ME1 ;
  RECT 90.000 0.000 90.800 1.000 ;
 END
 ANTENNAPARTIALMETALAREA                  3.118 LAYER ME2 ;
 ANTENNAGATEAREA                          0.086 LAYER ME2 ;
 ANTENNAGATEAREA                          0.086 LAYER ME3 ;
 ANTENNAGATEAREA                          0.086 LAYER ME4 ;
 ANTENNADIFFAREA                          0.160 LAYER ME2 ;
 ANTENNADIFFAREA                          0.160 LAYER ME3 ;
 ANTENNADIFFAREA                          0.160 LAYER ME4 ;
 ANTENNAMAXAREACAR                       48.431 LAYER ME2 ;
 ANTENNAMAXAREACAR                       57.690 LAYER ME3 ;
 ANTENNAMAXAREACAR                       66.949 LAYER ME4 ;
END DI4
PIN DO3
  DIRECTION OUTPUT ;
 PORT
  LAYER ME4 ;
  RECT 83.600 0.000 84.400 1.000 ;
  LAYER ME3 ;
  RECT 83.600 0.000 84.400 1.000 ;
  LAYER ME2 ;
  RECT 83.600 0.000 84.400 1.000 ;
  LAYER ME1 ;
  RECT 83.600 0.000 84.400 1.000 ;
 END
 ANTENNAPARTIALMETALAREA                  4.148 LAYER ME2 ;
 ANTENNADIFFAREA                          5.472 LAYER ME2 ;
 ANTENNADIFFAREA                          5.472 LAYER ME3 ;
 ANTENNADIFFAREA                          5.472 LAYER ME4 ;
END DO3
PIN DI3
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 68.800 0.000 69.600 1.000 ;
  LAYER ME3 ;
  RECT 68.800 0.000 69.600 1.000 ;
  LAYER ME2 ;
  RECT 68.800 0.000 69.600 1.000 ;
  LAYER ME1 ;
  RECT 68.800 0.000 69.600 1.000 ;
 END
 ANTENNAPARTIALMETALAREA                  3.142 LAYER ME2 ;
 ANTENNAGATEAREA                          0.086 LAYER ME2 ;
 ANTENNAGATEAREA                          0.086 LAYER ME3 ;
 ANTENNAGATEAREA                          0.086 LAYER ME4 ;
 ANTENNADIFFAREA                          0.160 LAYER ME2 ;
 ANTENNADIFFAREA                          0.160 LAYER ME3 ;
 ANTENNADIFFAREA                          0.160 LAYER ME4 ;
 ANTENNAMAXAREACAR                       48.708 LAYER ME2 ;
 ANTENNAMAXAREACAR                       57.968 LAYER ME3 ;
 ANTENNAMAXAREACAR                       67.227 LAYER ME4 ;
END DI3
PIN DO2
  DIRECTION OUTPUT ;
 PORT
  LAYER ME4 ;
  RECT 63.600 0.000 64.400 1.000 ;
  LAYER ME3 ;
  RECT 63.600 0.000 64.400 1.000 ;
  LAYER ME2 ;
  RECT 63.600 0.000 64.400 1.000 ;
  LAYER ME1 ;
  RECT 63.600 0.000 64.400 1.000 ;
 END
 ANTENNAPARTIALMETALAREA                  4.164 LAYER ME2 ;
 ANTENNADIFFAREA                          5.472 LAYER ME2 ;
 ANTENNADIFFAREA                          5.472 LAYER ME3 ;
 ANTENNADIFFAREA                          5.472 LAYER ME4 ;
END DO2
PIN DI2
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 49.200 0.000 50.000 1.000 ;
  LAYER ME3 ;
  RECT 49.200 0.000 50.000 1.000 ;
  LAYER ME2 ;
  RECT 49.200 0.000 50.000 1.000 ;
  LAYER ME1 ;
  RECT 49.200 0.000 50.000 1.000 ;
 END
 ANTENNAPARTIALMETALAREA                  3.138 LAYER ME2 ;
 ANTENNAGATEAREA                          0.086 LAYER ME2 ;
 ANTENNAGATEAREA                          0.086 LAYER ME3 ;
 ANTENNAGATEAREA                          0.086 LAYER ME4 ;
 ANTENNADIFFAREA                          0.160 LAYER ME2 ;
 ANTENNADIFFAREA                          0.160 LAYER ME3 ;
 ANTENNADIFFAREA                          0.160 LAYER ME4 ;
 ANTENNAMAXAREACAR                       48.662 LAYER ME2 ;
 ANTENNAMAXAREACAR                       57.921 LAYER ME3 ;
 ANTENNAMAXAREACAR                       67.181 LAYER ME4 ;
END DI2
PIN DO1
  DIRECTION OUTPUT ;
 PORT
  LAYER ME4 ;
  RECT 42.800 0.000 43.600 1.000 ;
  LAYER ME3 ;
  RECT 42.800 0.000 43.600 1.000 ;
  LAYER ME2 ;
  RECT 42.800 0.000 43.600 1.000 ;
  LAYER ME1 ;
  RECT 42.800 0.000 43.600 1.000 ;
 END
 ANTENNAPARTIALMETALAREA                  4.172 LAYER ME2 ;
 ANTENNADIFFAREA                          5.472 LAYER ME2 ;
 ANTENNADIFFAREA                          5.472 LAYER ME3 ;
 ANTENNADIFFAREA                          5.472 LAYER ME4 ;
END DO1
PIN DI1
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 28.000 0.000 28.800 1.000 ;
  LAYER ME3 ;
  RECT 28.000 0.000 28.800 1.000 ;
  LAYER ME2 ;
  RECT 28.000 0.000 28.800 1.000 ;
  LAYER ME1 ;
  RECT 28.000 0.000 28.800 1.000 ;
 END
 ANTENNAPARTIALMETALAREA                  3.118 LAYER ME2 ;
 ANTENNAGATEAREA                          0.086 LAYER ME2 ;
 ANTENNAGATEAREA                          0.086 LAYER ME3 ;
 ANTENNAGATEAREA                          0.086 LAYER ME4 ;
 ANTENNADIFFAREA                          0.160 LAYER ME2 ;
 ANTENNADIFFAREA                          0.160 LAYER ME3 ;
 ANTENNADIFFAREA                          0.160 LAYER ME4 ;
 ANTENNAMAXAREACAR                       48.431 LAYER ME2 ;
 ANTENNAMAXAREACAR                       57.690 LAYER ME3 ;
 ANTENNAMAXAREACAR                       66.949 LAYER ME4 ;
END DI1
PIN DO0
  DIRECTION OUTPUT ;
 PORT
  LAYER ME4 ;
  RECT 22.800 0.000 23.600 1.000 ;
  LAYER ME3 ;
  RECT 22.800 0.000 23.600 1.000 ;
  LAYER ME2 ;
  RECT 22.800 0.000 23.600 1.000 ;
  LAYER ME1 ;
  RECT 22.800 0.000 23.600 1.000 ;
 END
 ANTENNAPARTIALMETALAREA                  4.140 LAYER ME2 ;
 ANTENNADIFFAREA                          5.472 LAYER ME2 ;
 ANTENNADIFFAREA                          5.472 LAYER ME3 ;
 ANTENNADIFFAREA                          5.472 LAYER ME4 ;
END DO0
PIN WEB0
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 10.000 0.000 10.800 1.000 ;
  LAYER ME3 ;
  RECT 10.000 0.000 10.800 1.000 ;
  LAYER ME2 ;
  RECT 10.000 0.000 10.800 1.000 ;
  LAYER ME1 ;
  RECT 10.000 0.000 10.800 1.000 ;
 END
 ANTENNAPARTIALMETALAREA                  2.852 LAYER ME2 ;
 ANTENNAGATEAREA                          0.072 LAYER ME2 ;
 ANTENNAGATEAREA                          0.072 LAYER ME3 ;
 ANTENNAGATEAREA                          0.072 LAYER ME4 ;
 ANTENNADIFFAREA                          0.160 LAYER ME2 ;
 ANTENNADIFFAREA                          0.160 LAYER ME3 ;
 ANTENNADIFFAREA                          0.160 LAYER ME4 ;
 ANTENNAMAXAREACAR                       54.622 LAYER ME2 ;
 ANTENNAMAXAREACAR                       65.733 LAYER ME3 ;
 ANTENNAMAXAREACAR                       76.844 LAYER ME4 ;
END WEB0
PIN DI0
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 8.000 0.000 8.800 1.000 ;
  LAYER ME3 ;
  RECT 8.000 0.000 8.800 1.000 ;
  LAYER ME2 ;
  RECT 8.000 0.000 8.800 1.000 ;
  LAYER ME1 ;
  RECT 8.000 0.000 8.800 1.000 ;
 END
 ANTENNAPARTIALMETALAREA                  3.150 LAYER ME2 ;
 ANTENNAGATEAREA                          0.086 LAYER ME2 ;
 ANTENNAGATEAREA                          0.086 LAYER ME3 ;
 ANTENNAGATEAREA                          0.086 LAYER ME4 ;
 ANTENNADIFFAREA                          0.160 LAYER ME2 ;
 ANTENNADIFFAREA                          0.160 LAYER ME3 ;
 ANTENNADIFFAREA                          0.160 LAYER ME4 ;
 ANTENNAMAXAREACAR                       48.801 LAYER ME2 ;
 ANTENNAMAXAREACAR                       58.060 LAYER ME3 ;
 ANTENNAMAXAREACAR                       67.319 LAYER ME4 ;
END DI0
PIN VCC
  DIRECTION INOUT ;
  USE POWER ;
  SHAPE RING ;
 PORT
  LAYER ME4 ;
  RECT 2.000 193.930 2682.940 195.930 ;
  RECT 2.000 3.600 2682.940 5.600 ;
  RECT 2680.940 3.600 2682.940 195.930 ;
  RECT 2.000 3.600 4.000 195.930 ;
 END
END VCC
PIN GND
  DIRECTION INOUT ;
  USE GROUND ;
  SHAPE RING ;
 PORT
  LAYER ME3 ;
  RECT 0.000 195.930 2684.940 197.930 ;
  RECT 0.000 1.600 2684.940 3.600 ;
  RECT 2682.940 1.600 2684.940 197.930 ;
  RECT 0.000 1.600 2.000 197.930 ;
 END
END GND
OBS
  LAYER ME4 ;
  RECT 5.420 7.020 2679.520 192.510 ;
  RECT 2680.940 5.600 2682.940 193.930 ;
  RECT 2.000 5.600 4.000 193.930 ;
  RECT 4.000 193.930 2680.940 195.930 ;
  RECT 4.000 3.600 2680.940 5.600 ;
  RECT 2.000 193.930 4.000 195.930 ;
  RECT 2680.940 3.600 2682.940 5.600 ;
  RECT 2680.940 193.930 2682.940 195.930 ;
  RECT 2.000 3.600 4.000 5.600 ;
  RECT 2672.800 0.000 2673.600 1.000 ;
  RECT 2658.400 0.000 2659.200 1.000 ;
  RECT 2653.200 0.000 2654.000 1.000 ;
  RECT 2638.400 0.000 2639.200 1.000 ;
  RECT 2632.000 0.000 2632.800 1.000 ;
  RECT 2617.600 0.000 2618.400 1.000 ;
  RECT 2612.400 0.000 2613.200 1.000 ;
  RECT 2597.600 0.000 2598.400 1.000 ;
  RECT 2591.200 0.000 2592.000 1.000 ;
  RECT 2576.400 0.000 2577.200 1.000 ;
  RECT 2571.200 0.000 2572.000 1.000 ;
  RECT 2556.800 0.000 2557.600 1.000 ;
  RECT 2550.400 0.000 2551.200 1.000 ;
  RECT 2535.600 0.000 2536.400 1.000 ;
  RECT 2530.400 0.000 2531.200 1.000 ;
  RECT 2515.600 0.000 2516.400 1.000 ;
  RECT 2509.200 0.000 2510.000 1.000 ;
  RECT 2494.800 0.000 2495.600 1.000 ;
  RECT 2489.600 0.000 2490.400 1.000 ;
  RECT 2474.800 0.000 2475.600 1.000 ;
  RECT 2468.400 0.000 2469.200 1.000 ;
  RECT 2453.600 0.000 2454.400 1.000 ;
  RECT 2448.400 0.000 2449.200 1.000 ;
  RECT 2434.000 0.000 2434.800 1.000 ;
  RECT 2427.600 0.000 2428.400 1.000 ;
  RECT 2412.800 0.000 2413.600 1.000 ;
  RECT 2407.600 0.000 2408.400 1.000 ;
  RECT 2392.800 0.000 2393.600 1.000 ;
  RECT 2386.400 0.000 2387.200 1.000 ;
  RECT 2372.000 0.000 2372.800 1.000 ;
  RECT 2366.800 0.000 2367.600 1.000 ;
  RECT 2353.600 0.000 2354.400 1.000 ;
  RECT 2352.000 0.000 2352.800 1.000 ;
  RECT 2345.600 0.000 2346.400 1.000 ;
  RECT 2330.800 0.000 2331.600 1.000 ;
  RECT 2325.600 0.000 2326.400 1.000 ;
  RECT 2311.200 0.000 2312.000 1.000 ;
  RECT 2304.800 0.000 2305.600 1.000 ;
  RECT 2290.000 0.000 2290.800 1.000 ;
  RECT 2284.800 0.000 2285.600 1.000 ;
  RECT 2270.400 0.000 2271.200 1.000 ;
  RECT 2263.600 0.000 2264.400 1.000 ;
  RECT 2249.200 0.000 2250.000 1.000 ;
  RECT 2244.000 0.000 2244.800 1.000 ;
  RECT 2229.200 0.000 2230.000 1.000 ;
  RECT 2222.800 0.000 2223.600 1.000 ;
  RECT 2208.400 0.000 2209.200 1.000 ;
  RECT 2203.200 0.000 2204.000 1.000 ;
  RECT 2188.400 0.000 2189.200 1.000 ;
  RECT 2182.000 0.000 2182.800 1.000 ;
  RECT 2167.200 0.000 2168.000 1.000 ;
  RECT 2162.000 0.000 2162.800 1.000 ;
  RECT 2147.600 0.000 2148.400 1.000 ;
  RECT 2141.200 0.000 2142.000 1.000 ;
  RECT 2126.400 0.000 2127.200 1.000 ;
  RECT 2121.200 0.000 2122.000 1.000 ;
  RECT 2106.400 0.000 2107.200 1.000 ;
  RECT 2100.000 0.000 2100.800 1.000 ;
  RECT 2085.600 0.000 2086.400 1.000 ;
  RECT 2080.400 0.000 2081.200 1.000 ;
  RECT 2065.600 0.000 2066.400 1.000 ;
  RECT 2059.200 0.000 2060.000 1.000 ;
  RECT 2044.400 0.000 2045.200 1.000 ;
  RECT 2039.200 0.000 2040.000 1.000 ;
  RECT 2026.400 0.000 2027.200 1.000 ;
  RECT 2024.800 0.000 2025.600 1.000 ;
  RECT 2018.400 0.000 2019.200 1.000 ;
  RECT 2003.600 0.000 2004.400 1.000 ;
  RECT 1998.400 0.000 1999.200 1.000 ;
  RECT 1983.600 0.000 1984.400 1.000 ;
  RECT 1977.200 0.000 1978.000 1.000 ;
  RECT 1962.800 0.000 1963.600 1.000 ;
  RECT 1957.600 0.000 1958.400 1.000 ;
  RECT 1942.800 0.000 1943.600 1.000 ;
  RECT 1936.400 0.000 1937.200 1.000 ;
  RECT 1921.600 0.000 1922.400 1.000 ;
  RECT 1916.400 0.000 1917.200 1.000 ;
  RECT 1902.000 0.000 1902.800 1.000 ;
  RECT 1895.600 0.000 1896.400 1.000 ;
  RECT 1880.800 0.000 1881.600 1.000 ;
  RECT 1875.600 0.000 1876.400 1.000 ;
  RECT 1861.200 0.000 1862.000 1.000 ;
  RECT 1854.400 0.000 1855.200 1.000 ;
  RECT 1840.000 0.000 1840.800 1.000 ;
  RECT 1834.800 0.000 1835.600 1.000 ;
  RECT 1820.000 0.000 1820.800 1.000 ;
  RECT 1813.600 0.000 1814.400 1.000 ;
  RECT 1799.200 0.000 1800.000 1.000 ;
  RECT 1794.000 0.000 1794.800 1.000 ;
  RECT 1779.200 0.000 1780.000 1.000 ;
  RECT 1772.800 0.000 1773.600 1.000 ;
  RECT 1758.000 0.000 1758.800 1.000 ;
  RECT 1752.800 0.000 1753.600 1.000 ;
  RECT 1738.400 0.000 1739.200 1.000 ;
  RECT 1732.000 0.000 1732.800 1.000 ;
  RECT 1717.200 0.000 1718.000 1.000 ;
  RECT 1712.000 0.000 1712.800 1.000 ;
  RECT 1699.200 0.000 1700.000 1.000 ;
  RECT 1697.200 0.000 1698.000 1.000 ;
  RECT 1690.800 0.000 1691.600 1.000 ;
  RECT 1676.400 0.000 1677.200 1.000 ;
  RECT 1671.200 0.000 1672.000 1.000 ;
  RECT 1656.400 0.000 1657.200 1.000 ;
  RECT 1650.000 0.000 1650.800 1.000 ;
  RECT 1635.200 0.000 1636.000 1.000 ;
  RECT 1630.000 0.000 1630.800 1.000 ;
  RECT 1615.600 0.000 1616.400 1.000 ;
  RECT 1609.200 0.000 1610.000 1.000 ;
  RECT 1594.400 0.000 1595.200 1.000 ;
  RECT 1589.200 0.000 1590.000 1.000 ;
  RECT 1574.400 0.000 1575.200 1.000 ;
  RECT 1568.000 0.000 1568.800 1.000 ;
  RECT 1553.600 0.000 1554.400 1.000 ;
  RECT 1548.400 0.000 1549.200 1.000 ;
  RECT 1533.600 0.000 1534.400 1.000 ;
  RECT 1527.200 0.000 1528.000 1.000 ;
  RECT 1512.400 0.000 1513.200 1.000 ;
  RECT 1507.200 0.000 1508.000 1.000 ;
  RECT 1492.800 0.000 1493.600 1.000 ;
  RECT 1486.400 0.000 1487.200 1.000 ;
  RECT 1471.600 0.000 1472.400 1.000 ;
  RECT 1466.400 0.000 1467.200 1.000 ;
  RECT 1452.000 0.000 1452.800 1.000 ;
  RECT 1445.200 0.000 1446.000 1.000 ;
  RECT 1430.800 0.000 1431.600 1.000 ;
  RECT 1425.600 0.000 1426.400 1.000 ;
  RECT 1410.800 0.000 1411.600 1.000 ;
  RECT 1404.400 0.000 1405.200 1.000 ;
  RECT 1390.000 0.000 1390.800 1.000 ;
  RECT 1384.800 0.000 1385.600 1.000 ;
  RECT 1371.600 0.000 1372.400 1.000 ;
  RECT 1370.000 0.000 1370.800 1.000 ;
  RECT 1349.200 0.000 1350.000 1.000 ;
  RECT 1348.000 0.000 1348.800 1.000 ;
  RECT 1346.800 0.000 1347.600 1.000 ;
  RECT 1345.600 0.000 1346.400 1.000 ;
  RECT 1344.400 0.000 1345.200 1.000 ;
  RECT 1343.200 0.000 1344.000 1.000 ;
  RECT 1337.200 0.000 1338.000 1.000 ;
  RECT 1330.000 0.000 1330.800 1.000 ;
  RECT 1327.200 0.000 1328.000 1.000 ;
  RECT 1324.400 0.000 1325.200 1.000 ;
  RECT 1322.000 0.000 1322.800 1.000 ;
  RECT 1320.400 0.000 1321.200 1.000 ;
  RECT 1318.000 0.000 1318.800 1.000 ;
  RECT 1311.200 0.000 1312.000 1.000 ;
  RECT 1296.400 0.000 1297.200 1.000 ;
  RECT 1291.200 0.000 1292.000 1.000 ;
  RECT 1276.800 0.000 1277.600 1.000 ;
  RECT 1270.400 0.000 1271.200 1.000 ;
  RECT 1255.600 0.000 1256.400 1.000 ;
  RECT 1250.400 0.000 1251.200 1.000 ;
  RECT 1235.600 0.000 1236.400 1.000 ;
  RECT 1229.200 0.000 1230.000 1.000 ;
  RECT 1214.800 0.000 1215.600 1.000 ;
  RECT 1209.600 0.000 1210.400 1.000 ;
  RECT 1194.800 0.000 1195.600 1.000 ;
  RECT 1188.400 0.000 1189.200 1.000 ;
  RECT 1173.600 0.000 1174.400 1.000 ;
  RECT 1168.400 0.000 1169.200 1.000 ;
  RECT 1154.000 0.000 1154.800 1.000 ;
  RECT 1147.600 0.000 1148.400 1.000 ;
  RECT 1132.800 0.000 1133.600 1.000 ;
  RECT 1127.600 0.000 1128.400 1.000 ;
  RECT 1113.200 0.000 1114.000 1.000 ;
  RECT 1106.400 0.000 1107.200 1.000 ;
  RECT 1092.000 0.000 1092.800 1.000 ;
  RECT 1086.800 0.000 1087.600 1.000 ;
  RECT 1072.000 0.000 1072.800 1.000 ;
  RECT 1065.600 0.000 1066.400 1.000 ;
  RECT 1051.200 0.000 1052.000 1.000 ;
  RECT 1045.600 0.000 1046.400 1.000 ;
  RECT 1031.200 0.000 1032.000 1.000 ;
  RECT 1024.800 0.000 1025.600 1.000 ;
  RECT 1010.000 0.000 1010.800 1.000 ;
  RECT 1004.800 0.000 1005.600 1.000 ;
  RECT 992.000 0.000 992.800 1.000 ;
  RECT 990.400 0.000 991.200 1.000 ;
  RECT 983.600 0.000 984.400 1.000 ;
  RECT 969.200 0.000 970.000 1.000 ;
  RECT 964.000 0.000 964.800 1.000 ;
  RECT 949.200 0.000 950.000 1.000 ;
  RECT 942.800 0.000 943.600 1.000 ;
  RECT 928.400 0.000 929.200 1.000 ;
  RECT 923.200 0.000 924.000 1.000 ;
  RECT 908.400 0.000 909.200 1.000 ;
  RECT 902.000 0.000 902.800 1.000 ;
  RECT 887.200 0.000 888.000 1.000 ;
  RECT 882.000 0.000 882.800 1.000 ;
  RECT 867.600 0.000 868.400 1.000 ;
  RECT 861.200 0.000 862.000 1.000 ;
  RECT 846.400 0.000 847.200 1.000 ;
  RECT 841.200 0.000 842.000 1.000 ;
  RECT 826.400 0.000 827.200 1.000 ;
  RECT 820.000 0.000 820.800 1.000 ;
  RECT 805.600 0.000 806.400 1.000 ;
  RECT 800.400 0.000 801.200 1.000 ;
  RECT 785.600 0.000 786.400 1.000 ;
  RECT 779.200 0.000 780.000 1.000 ;
  RECT 764.400 0.000 765.200 1.000 ;
  RECT 759.200 0.000 760.000 1.000 ;
  RECT 744.800 0.000 745.600 1.000 ;
  RECT 738.400 0.000 739.200 1.000 ;
  RECT 723.600 0.000 724.400 1.000 ;
  RECT 718.400 0.000 719.200 1.000 ;
  RECT 704.000 0.000 704.800 1.000 ;
  RECT 697.200 0.000 698.000 1.000 ;
  RECT 682.800 0.000 683.600 1.000 ;
  RECT 677.600 0.000 678.400 1.000 ;
  RECT 664.800 0.000 665.600 1.000 ;
  RECT 662.800 0.000 663.600 1.000 ;
  RECT 656.400 0.000 657.200 1.000 ;
  RECT 642.000 0.000 642.800 1.000 ;
  RECT 636.400 0.000 637.200 1.000 ;
  RECT 622.000 0.000 622.800 1.000 ;
  RECT 615.600 0.000 616.400 1.000 ;
  RECT 600.800 0.000 601.600 1.000 ;
  RECT 595.600 0.000 596.400 1.000 ;
  RECT 581.200 0.000 582.000 1.000 ;
  RECT 574.400 0.000 575.200 1.000 ;
  RECT 560.000 0.000 560.800 1.000 ;
  RECT 554.800 0.000 555.600 1.000 ;
  RECT 540.000 0.000 540.800 1.000 ;
  RECT 533.600 0.000 534.400 1.000 ;
  RECT 519.200 0.000 520.000 1.000 ;
  RECT 514.000 0.000 514.800 1.000 ;
  RECT 499.200 0.000 500.000 1.000 ;
  RECT 492.800 0.000 493.600 1.000 ;
  RECT 478.000 0.000 478.800 1.000 ;
  RECT 472.800 0.000 473.600 1.000 ;
  RECT 458.400 0.000 459.200 1.000 ;
  RECT 452.000 0.000 452.800 1.000 ;
  RECT 437.200 0.000 438.000 1.000 ;
  RECT 432.000 0.000 432.800 1.000 ;
  RECT 417.200 0.000 418.000 1.000 ;
  RECT 410.800 0.000 411.600 1.000 ;
  RECT 396.400 0.000 397.200 1.000 ;
  RECT 391.200 0.000 392.000 1.000 ;
  RECT 376.400 0.000 377.200 1.000 ;
  RECT 370.000 0.000 370.800 1.000 ;
  RECT 355.200 0.000 356.000 1.000 ;
  RECT 350.000 0.000 350.800 1.000 ;
  RECT 337.200 0.000 338.000 1.000 ;
  RECT 335.600 0.000 336.400 1.000 ;
  RECT 329.200 0.000 330.000 1.000 ;
  RECT 314.400 0.000 315.200 1.000 ;
  RECT 309.200 0.000 310.000 1.000 ;
  RECT 294.800 0.000 295.600 1.000 ;
  RECT 288.000 0.000 288.800 1.000 ;
  RECT 273.600 0.000 274.400 1.000 ;
  RECT 268.400 0.000 269.200 1.000 ;
  RECT 253.600 0.000 254.400 1.000 ;
  RECT 247.200 0.000 248.000 1.000 ;
  RECT 232.800 0.000 233.600 1.000 ;
  RECT 227.200 0.000 228.000 1.000 ;
  RECT 212.800 0.000 213.600 1.000 ;
  RECT 206.400 0.000 207.200 1.000 ;
  RECT 191.600 0.000 192.400 1.000 ;
  RECT 186.400 0.000 187.200 1.000 ;
  RECT 172.000 0.000 172.800 1.000 ;
  RECT 165.200 0.000 166.000 1.000 ;
  RECT 150.800 0.000 151.600 1.000 ;
  RECT 145.600 0.000 146.400 1.000 ;
  RECT 130.800 0.000 131.600 1.000 ;
  RECT 124.400 0.000 125.200 1.000 ;
  RECT 110.000 0.000 110.800 1.000 ;
  RECT 104.800 0.000 105.600 1.000 ;
  RECT 90.000 0.000 90.800 1.000 ;
  RECT 83.600 0.000 84.400 1.000 ;
  RECT 68.800 0.000 69.600 1.000 ;
  RECT 63.600 0.000 64.400 1.000 ;
  RECT 49.200 0.000 50.000 1.000 ;
  RECT 42.800 0.000 43.600 1.000 ;
  RECT 28.000 0.000 28.800 1.000 ;
  RECT 22.800 0.000 23.600 1.000 ;
  RECT 10.000 0.000 10.800 1.000 ;
  RECT 8.000 0.000 8.800 1.000 ;
  RECT 2679.800 9.570 2680.940 11.170 ;
  RECT 2679.800 14.200 2680.940 15.200 ;
  RECT 2679.800 18.730 2680.940 19.730 ;
  RECT 2679.800 21.230 2680.940 22.070 ;
  RECT 2679.800 24.170 2680.940 25.170 ;
  RECT 2679.800 36.320 2680.940 37.320 ;
  RECT 2679.800 39.480 2680.940 40.080 ;
  RECT 2679.800 45.560 2680.940 46.160 ;
  RECT 2679.800 57.100 2680.940 61.420 ;
  RECT 2678.380 5.880 2679.520 7.020 ;
  RECT 1380.220 5.600 1388.220 7.020 ;
  RECT 1370.180 5.880 1378.180 7.020 ;
  RECT 1390.020 5.880 1398.020 7.020 ;
  RECT 1400.060 5.600 1408.060 7.020 ;
  RECT 1411.100 5.880 1419.100 7.020 ;
  RECT 1421.140 5.600 1429.140 7.020 ;
  RECT 1430.940 5.880 1438.940 7.020 ;
  RECT 1440.980 5.600 1448.980 7.020 ;
  RECT 1452.020 5.880 1460.020 7.020 ;
  RECT 1462.060 5.600 1470.060 7.020 ;
  RECT 1471.860 5.880 1479.860 7.020 ;
  RECT 1481.900 5.600 1489.900 7.020 ;
  RECT 1492.940 5.880 1500.940 7.020 ;
  RECT 1502.980 5.600 1510.980 7.020 ;
  RECT 1512.780 5.880 1520.780 7.020 ;
  RECT 1522.820 5.600 1530.820 7.020 ;
  RECT 1533.860 5.880 1541.860 7.020 ;
  RECT 1543.900 5.600 1551.900 7.020 ;
  RECT 1553.700 5.880 1561.700 7.020 ;
  RECT 1563.740 5.600 1571.740 7.020 ;
  RECT 1574.780 5.880 1582.780 7.020 ;
  RECT 1584.820 5.600 1592.820 7.020 ;
  RECT 1594.620 5.880 1602.620 7.020 ;
  RECT 1604.660 5.600 1612.660 7.020 ;
  RECT 1615.700 5.880 1623.700 7.020 ;
  RECT 1625.740 5.600 1633.740 7.020 ;
  RECT 1635.540 5.880 1643.540 7.020 ;
  RECT 1645.580 5.600 1653.580 7.020 ;
  RECT 1656.620 5.880 1664.620 7.020 ;
  RECT 1666.660 5.600 1674.660 7.020 ;
  RECT 1676.460 5.880 1684.460 7.020 ;
  RECT 1686.500 5.600 1694.500 7.020 ;
  RECT 1707.580 5.600 1715.580 7.020 ;
  RECT 1697.540 5.880 1705.540 7.020 ;
  RECT 1717.380 5.880 1725.380 7.020 ;
  RECT 1727.420 5.600 1735.420 7.020 ;
  RECT 1738.460 5.880 1746.460 7.020 ;
  RECT 1748.500 5.600 1756.500 7.020 ;
  RECT 1758.300 5.880 1766.300 7.020 ;
  RECT 1768.340 5.600 1776.340 7.020 ;
  RECT 1779.380 5.880 1787.380 7.020 ;
  RECT 1789.420 5.600 1797.420 7.020 ;
  RECT 1799.220 5.880 1807.220 7.020 ;
  RECT 1809.260 5.600 1817.260 7.020 ;
  RECT 1820.300 5.880 1828.300 7.020 ;
  RECT 1830.340 5.600 1838.340 7.020 ;
  RECT 1840.140 5.880 1848.140 7.020 ;
  RECT 1850.180 5.600 1858.180 7.020 ;
  RECT 1861.220 5.880 1869.220 7.020 ;
  RECT 1871.260 5.600 1879.260 7.020 ;
  RECT 1881.060 5.880 1889.060 7.020 ;
  RECT 1891.100 5.600 1899.100 7.020 ;
  RECT 1902.140 5.880 1910.140 7.020 ;
  RECT 1912.180 5.600 1920.180 7.020 ;
  RECT 1921.980 5.880 1929.980 7.020 ;
  RECT 1932.020 5.600 1940.020 7.020 ;
  RECT 1943.060 5.880 1951.060 7.020 ;
  RECT 1953.100 5.600 1961.100 7.020 ;
  RECT 1962.900 5.880 1970.900 7.020 ;
  RECT 1972.940 5.600 1980.940 7.020 ;
  RECT 1983.980 5.880 1991.980 7.020 ;
  RECT 1994.020 5.600 2002.020 7.020 ;
  RECT 2003.820 5.880 2011.820 7.020 ;
  RECT 2013.860 5.600 2021.860 7.020 ;
  RECT 2034.940 5.600 2042.940 7.020 ;
  RECT 2024.900 5.880 2032.900 7.020 ;
  RECT 2044.740 5.880 2052.740 7.020 ;
  RECT 2054.780 5.600 2062.780 7.020 ;
  RECT 2065.820 5.880 2073.820 7.020 ;
  RECT 2075.860 5.600 2083.860 7.020 ;
  RECT 2085.660 5.880 2093.660 7.020 ;
  RECT 2095.700 5.600 2103.700 7.020 ;
  RECT 2106.740 5.880 2114.740 7.020 ;
  RECT 2116.780 5.600 2124.780 7.020 ;
  RECT 2126.580 5.880 2134.580 7.020 ;
  RECT 2136.620 5.600 2144.620 7.020 ;
  RECT 2147.660 5.880 2155.660 7.020 ;
  RECT 2157.700 5.600 2165.700 7.020 ;
  RECT 2167.500 5.880 2175.500 7.020 ;
  RECT 2177.540 5.600 2185.540 7.020 ;
  RECT 2188.580 5.880 2196.580 7.020 ;
  RECT 2198.620 5.600 2206.620 7.020 ;
  RECT 2208.420 5.880 2216.420 7.020 ;
  RECT 2218.460 5.600 2226.460 7.020 ;
  RECT 2229.500 5.880 2237.500 7.020 ;
  RECT 2239.540 5.600 2247.540 7.020 ;
  RECT 2249.340 5.880 2257.340 7.020 ;
  RECT 2259.380 5.600 2267.380 7.020 ;
  RECT 2270.420 5.880 2278.420 7.020 ;
  RECT 2280.460 5.600 2288.460 7.020 ;
  RECT 2290.260 5.880 2298.260 7.020 ;
  RECT 2300.300 5.600 2308.300 7.020 ;
  RECT 2311.340 5.880 2319.340 7.020 ;
  RECT 2321.380 5.600 2329.380 7.020 ;
  RECT 2331.180 5.880 2339.180 7.020 ;
  RECT 2341.220 5.600 2349.220 7.020 ;
  RECT 2362.300 5.600 2370.300 7.020 ;
  RECT 2352.260 5.880 2360.260 7.020 ;
  RECT 2372.100 5.880 2380.100 7.020 ;
  RECT 2382.140 5.600 2390.140 7.020 ;
  RECT 2393.180 5.880 2401.180 7.020 ;
  RECT 2403.220 5.600 2411.220 7.020 ;
  RECT 2413.020 5.880 2421.020 7.020 ;
  RECT 2423.060 5.600 2431.060 7.020 ;
  RECT 2434.100 5.880 2442.100 7.020 ;
  RECT 2444.140 5.600 2452.140 7.020 ;
  RECT 2453.940 5.880 2461.940 7.020 ;
  RECT 2463.980 5.600 2471.980 7.020 ;
  RECT 2475.020 5.880 2483.020 7.020 ;
  RECT 2485.060 5.600 2493.060 7.020 ;
  RECT 2494.860 5.880 2502.860 7.020 ;
  RECT 2504.900 5.600 2512.900 7.020 ;
  RECT 2515.940 5.880 2523.940 7.020 ;
  RECT 2525.980 5.600 2533.980 7.020 ;
  RECT 2535.780 5.880 2543.780 7.020 ;
  RECT 2545.820 5.600 2553.820 7.020 ;
  RECT 2556.860 5.880 2564.860 7.020 ;
  RECT 2566.900 5.600 2574.900 7.020 ;
  RECT 2576.700 5.880 2584.700 7.020 ;
  RECT 2586.740 5.600 2594.740 7.020 ;
  RECT 2597.780 5.880 2605.780 7.020 ;
  RECT 2607.820 5.600 2615.820 7.020 ;
  RECT 2617.620 5.880 2625.620 7.020 ;
  RECT 2627.660 5.600 2635.660 7.020 ;
  RECT 2638.700 5.880 2646.700 7.020 ;
  RECT 2648.740 5.600 2656.740 7.020 ;
  RECT 2658.540 5.880 2666.540 7.020 ;
  RECT 2668.580 5.600 2676.580 7.020 ;
  RECT 1331.880 5.600 1334.940 7.020 ;
  RECT 1335.440 5.880 1338.890 7.020 ;
  RECT 1339.390 5.600 1343.140 7.020 ;
  RECT 1344.290 5.880 1350.210 7.020 ;
  RECT 1351.360 5.600 1355.110 7.020 ;
  RECT 1355.610 5.600 1359.360 7.020 ;
  RECT 1359.860 5.600 1363.610 7.020 ;
  RECT 1329.160 5.600 1330.920 7.020 ;
  RECT 1327.160 5.880 1328.920 7.020 ;
  RECT 1323.820 5.600 1325.580 7.020 ;
  RECT 1321.820 5.880 1323.580 7.020 ;
  RECT 1319.820 5.600 1321.580 7.020 ;
  RECT 1317.820 5.880 1319.580 7.020 ;
  RECT 4.000 57.100 5.140 61.420 ;
  RECT 4.000 45.560 5.140 46.160 ;
  RECT 4.000 39.480 5.140 40.080 ;
  RECT 4.000 36.320 5.140 37.320 ;
  RECT 4.000 24.170 5.140 25.170 ;
  RECT 4.000 21.230 5.140 22.070 ;
  RECT 4.000 18.730 5.140 19.730 ;
  RECT 4.000 14.200 5.140 15.200 ;
  RECT 4.000 9.570 5.140 11.170 ;
  RECT 5.420 5.880 6.560 7.020 ;
  RECT 18.400 5.600 26.400 7.020 ;
  RECT 8.360 5.880 16.360 7.020 ;
  RECT 28.200 5.880 36.200 7.020 ;
  RECT 38.240 5.600 46.240 7.020 ;
  RECT 49.280 5.880 57.280 7.020 ;
  RECT 59.320 5.600 67.320 7.020 ;
  RECT 69.120 5.880 77.120 7.020 ;
  RECT 79.160 5.600 87.160 7.020 ;
  RECT 90.200 5.880 98.200 7.020 ;
  RECT 100.240 5.600 108.240 7.020 ;
  RECT 110.040 5.880 118.040 7.020 ;
  RECT 120.080 5.600 128.080 7.020 ;
  RECT 131.120 5.880 139.120 7.020 ;
  RECT 141.160 5.600 149.160 7.020 ;
  RECT 150.960 5.880 158.960 7.020 ;
  RECT 161.000 5.600 169.000 7.020 ;
  RECT 172.040 5.880 180.040 7.020 ;
  RECT 182.080 5.600 190.080 7.020 ;
  RECT 191.880 5.880 199.880 7.020 ;
  RECT 201.920 5.600 209.920 7.020 ;
  RECT 212.960 5.880 220.960 7.020 ;
  RECT 223.000 5.600 231.000 7.020 ;
  RECT 232.800 5.880 240.800 7.020 ;
  RECT 242.840 5.600 250.840 7.020 ;
  RECT 253.880 5.880 261.880 7.020 ;
  RECT 263.920 5.600 271.920 7.020 ;
  RECT 273.720 5.880 281.720 7.020 ;
  RECT 283.760 5.600 291.760 7.020 ;
  RECT 294.800 5.880 302.800 7.020 ;
  RECT 304.840 5.600 312.840 7.020 ;
  RECT 314.640 5.880 322.640 7.020 ;
  RECT 324.680 5.600 332.680 7.020 ;
  RECT 345.760 5.600 353.760 7.020 ;
  RECT 335.720 5.880 343.720 7.020 ;
  RECT 355.560 5.880 363.560 7.020 ;
  RECT 365.600 5.600 373.600 7.020 ;
  RECT 376.640 5.880 384.640 7.020 ;
  RECT 386.680 5.600 394.680 7.020 ;
  RECT 396.480 5.880 404.480 7.020 ;
  RECT 406.520 5.600 414.520 7.020 ;
  RECT 417.560 5.880 425.560 7.020 ;
  RECT 427.600 5.600 435.600 7.020 ;
  RECT 437.400 5.880 445.400 7.020 ;
  RECT 447.440 5.600 455.440 7.020 ;
  RECT 458.480 5.880 466.480 7.020 ;
  RECT 468.520 5.600 476.520 7.020 ;
  RECT 478.320 5.880 486.320 7.020 ;
  RECT 488.360 5.600 496.360 7.020 ;
  RECT 499.400 5.880 507.400 7.020 ;
  RECT 509.440 5.600 517.440 7.020 ;
  RECT 519.240 5.880 527.240 7.020 ;
  RECT 529.280 5.600 537.280 7.020 ;
  RECT 540.320 5.880 548.320 7.020 ;
  RECT 550.360 5.600 558.360 7.020 ;
  RECT 560.160 5.880 568.160 7.020 ;
  RECT 570.200 5.600 578.200 7.020 ;
  RECT 581.240 5.880 589.240 7.020 ;
  RECT 591.280 5.600 599.280 7.020 ;
  RECT 601.080 5.880 609.080 7.020 ;
  RECT 611.120 5.600 619.120 7.020 ;
  RECT 622.160 5.880 630.160 7.020 ;
  RECT 632.200 5.600 640.200 7.020 ;
  RECT 642.000 5.880 650.000 7.020 ;
  RECT 652.040 5.600 660.040 7.020 ;
  RECT 673.120 5.600 681.120 7.020 ;
  RECT 663.080 5.880 671.080 7.020 ;
  RECT 682.920 5.880 690.920 7.020 ;
  RECT 692.960 5.600 700.960 7.020 ;
  RECT 704.000 5.880 712.000 7.020 ;
  RECT 714.040 5.600 722.040 7.020 ;
  RECT 723.840 5.880 731.840 7.020 ;
  RECT 733.880 5.600 741.880 7.020 ;
  RECT 744.920 5.880 752.920 7.020 ;
  RECT 754.960 5.600 762.960 7.020 ;
  RECT 764.760 5.880 772.760 7.020 ;
  RECT 774.800 5.600 782.800 7.020 ;
  RECT 785.840 5.880 793.840 7.020 ;
  RECT 795.880 5.600 803.880 7.020 ;
  RECT 805.680 5.880 813.680 7.020 ;
  RECT 815.720 5.600 823.720 7.020 ;
  RECT 826.760 5.880 834.760 7.020 ;
  RECT 836.800 5.600 844.800 7.020 ;
  RECT 846.600 5.880 854.600 7.020 ;
  RECT 856.640 5.600 864.640 7.020 ;
  RECT 867.680 5.880 875.680 7.020 ;
  RECT 877.720 5.600 885.720 7.020 ;
  RECT 887.520 5.880 895.520 7.020 ;
  RECT 897.560 5.600 905.560 7.020 ;
  RECT 908.600 5.880 916.600 7.020 ;
  RECT 918.640 5.600 926.640 7.020 ;
  RECT 928.440 5.880 936.440 7.020 ;
  RECT 938.480 5.600 946.480 7.020 ;
  RECT 949.520 5.880 957.520 7.020 ;
  RECT 959.560 5.600 967.560 7.020 ;
  RECT 969.360 5.880 977.360 7.020 ;
  RECT 979.400 5.600 987.400 7.020 ;
  RECT 1000.480 5.600 1008.480 7.020 ;
  RECT 990.440 5.880 998.440 7.020 ;
  RECT 1010.280 5.880 1018.280 7.020 ;
  RECT 1020.320 5.600 1028.320 7.020 ;
  RECT 1031.360 5.880 1039.360 7.020 ;
  RECT 1041.400 5.600 1049.400 7.020 ;
  RECT 1051.200 5.880 1059.200 7.020 ;
  RECT 1061.240 5.600 1069.240 7.020 ;
  RECT 1072.280 5.880 1080.280 7.020 ;
  RECT 1082.320 5.600 1090.320 7.020 ;
  RECT 1092.120 5.880 1100.120 7.020 ;
  RECT 1102.160 5.600 1110.160 7.020 ;
  RECT 1113.200 5.880 1121.200 7.020 ;
  RECT 1123.240 5.600 1131.240 7.020 ;
  RECT 1133.040 5.880 1141.040 7.020 ;
  RECT 1143.080 5.600 1151.080 7.020 ;
  RECT 1154.120 5.880 1162.120 7.020 ;
  RECT 1164.160 5.600 1172.160 7.020 ;
  RECT 1173.960 5.880 1181.960 7.020 ;
  RECT 1184.000 5.600 1192.000 7.020 ;
  RECT 1195.040 5.880 1203.040 7.020 ;
  RECT 1205.080 5.600 1213.080 7.020 ;
  RECT 1214.880 5.880 1222.880 7.020 ;
  RECT 1224.920 5.600 1232.920 7.020 ;
  RECT 1235.960 5.880 1243.960 7.020 ;
  RECT 1246.000 5.600 1254.000 7.020 ;
  RECT 1255.800 5.880 1263.800 7.020 ;
  RECT 1265.840 5.600 1273.840 7.020 ;
  RECT 1276.880 5.880 1284.880 7.020 ;
  RECT 1286.920 5.600 1294.920 7.020 ;
  RECT 1296.720 5.880 1304.720 7.020 ;
  RECT 1306.760 5.600 1314.760 7.020 ;
  RECT 2679.800 191.940 2680.940 192.320 ;
  RECT 2679.800 184.020 2680.940 184.300 ;
  RECT 2679.800 180.340 2680.940 180.620 ;
  RECT 2679.800 176.660 2680.940 176.940 ;
  RECT 2679.800 172.980 2680.940 173.260 ;
  RECT 2679.800 169.300 2680.940 169.580 ;
  RECT 2679.800 165.620 2680.940 165.900 ;
  RECT 2679.800 161.940 2680.940 162.220 ;
  RECT 2679.800 158.260 2680.940 158.540 ;
  RECT 2679.800 154.580 2680.940 154.860 ;
  RECT 2679.800 150.900 2680.940 151.180 ;
  RECT 2679.800 147.220 2680.940 147.500 ;
  RECT 2679.800 143.540 2680.940 143.820 ;
  RECT 2679.800 139.860 2680.940 140.140 ;
  RECT 2679.800 136.180 2680.940 136.460 ;
  RECT 2679.800 132.500 2680.940 132.780 ;
  RECT 2679.800 128.820 2680.940 129.100 ;
  RECT 2679.800 125.140 2680.940 125.420 ;
  RECT 2679.800 121.460 2680.940 121.740 ;
  RECT 2679.800 117.780 2680.940 118.060 ;
  RECT 2679.800 114.100 2680.940 114.380 ;
  RECT 2679.800 110.420 2680.940 110.700 ;
  RECT 2679.800 106.740 2680.940 107.020 ;
  RECT 2679.800 103.060 2680.940 103.340 ;
  RECT 2679.800 99.380 2680.940 99.660 ;
  RECT 2679.800 95.700 2680.940 95.980 ;
  RECT 2679.800 92.020 2680.940 92.300 ;
  RECT 2679.800 88.340 2680.940 88.620 ;
  RECT 2679.800 84.660 2680.940 84.940 ;
  RECT 2679.800 80.980 2680.940 81.260 ;
  RECT 2679.800 77.300 2680.940 77.580 ;
  RECT 2679.800 73.620 2680.940 73.900 ;
  RECT 2679.800 69.940 2680.940 70.220 ;
  RECT 2679.800 65.600 2680.940 65.980 ;
  RECT 1368.820 192.790 1369.070 193.930 ;
  RECT 1409.740 192.790 1409.990 193.930 ;
  RECT 1450.660 192.790 1450.910 193.930 ;
  RECT 1491.580 192.790 1491.830 193.930 ;
  RECT 1532.500 192.790 1532.750 193.930 ;
  RECT 1573.420 192.790 1573.670 193.930 ;
  RECT 1614.340 192.790 1614.590 193.930 ;
  RECT 1655.260 192.790 1655.510 193.930 ;
  RECT 1696.180 192.790 1696.430 193.930 ;
  RECT 1737.100 192.790 1737.350 193.930 ;
  RECT 1778.020 192.790 1778.270 193.930 ;
  RECT 1818.940 192.790 1819.190 193.930 ;
  RECT 1859.860 192.790 1860.110 193.930 ;
  RECT 1900.780 192.790 1901.030 193.930 ;
  RECT 1941.700 192.790 1941.950 193.930 ;
  RECT 1982.620 192.790 1982.870 193.930 ;
  RECT 2023.540 192.790 2023.790 193.930 ;
  RECT 2064.460 192.790 2064.710 193.930 ;
  RECT 2105.380 192.790 2105.630 193.930 ;
  RECT 2146.300 192.790 2146.550 193.930 ;
  RECT 2187.220 192.790 2187.470 193.930 ;
  RECT 2228.140 192.790 2228.390 193.930 ;
  RECT 2269.060 192.790 2269.310 193.930 ;
  RECT 2309.980 192.790 2310.230 193.930 ;
  RECT 2350.900 192.790 2351.150 193.930 ;
  RECT 2391.820 192.790 2392.070 193.930 ;
  RECT 2432.740 192.790 2432.990 193.930 ;
  RECT 2473.660 192.790 2473.910 193.930 ;
  RECT 2514.580 192.790 2514.830 193.930 ;
  RECT 2555.500 192.790 2555.750 193.930 ;
  RECT 2596.420 192.790 2596.670 193.930 ;
  RECT 2637.340 192.790 2637.590 193.930 ;
  RECT 1351.810 192.790 1354.320 193.930 ;
  RECT 1339.390 192.790 1341.780 193.930 ;
  RECT 1331.880 192.790 1334.940 193.930 ;
  RECT 1356.060 192.790 1358.910 193.930 ;
  RECT 1360.360 192.790 1363.610 193.930 ;
  RECT 1329.160 192.790 1330.920 193.930 ;
  RECT 1319.820 192.790 1321.580 193.930 ;
  RECT 1323.820 192.790 1325.580 193.930 ;
  RECT 4.000 65.600 5.140 65.980 ;
  RECT 4.000 69.940 5.140 70.220 ;
  RECT 4.000 73.620 5.140 73.900 ;
  RECT 4.000 77.300 5.140 77.580 ;
  RECT 4.000 80.980 5.140 81.260 ;
  RECT 4.000 84.660 5.140 84.940 ;
  RECT 4.000 88.340 5.140 88.620 ;
  RECT 4.000 92.020 5.140 92.300 ;
  RECT 4.000 95.700 5.140 95.980 ;
  RECT 4.000 99.380 5.140 99.660 ;
  RECT 4.000 103.060 5.140 103.340 ;
  RECT 4.000 106.740 5.140 107.020 ;
  RECT 4.000 110.420 5.140 110.700 ;
  RECT 4.000 114.100 5.140 114.380 ;
  RECT 4.000 117.780 5.140 118.060 ;
  RECT 4.000 121.460 5.140 121.740 ;
  RECT 4.000 125.140 5.140 125.420 ;
  RECT 4.000 128.820 5.140 129.100 ;
  RECT 4.000 132.500 5.140 132.780 ;
  RECT 4.000 136.180 5.140 136.460 ;
  RECT 4.000 139.860 5.140 140.140 ;
  RECT 4.000 143.540 5.140 143.820 ;
  RECT 4.000 147.220 5.140 147.500 ;
  RECT 4.000 150.900 5.140 151.180 ;
  RECT 4.000 154.580 5.140 154.860 ;
  RECT 4.000 158.260 5.140 158.540 ;
  RECT 4.000 161.940 5.140 162.220 ;
  RECT 4.000 165.620 5.140 165.900 ;
  RECT 4.000 169.300 5.140 169.580 ;
  RECT 4.000 172.980 5.140 173.260 ;
  RECT 4.000 176.660 5.140 176.940 ;
  RECT 4.000 180.340 5.140 180.620 ;
  RECT 4.000 184.020 5.140 184.300 ;
  RECT 4.000 191.940 5.140 192.320 ;
  RECT 47.350 192.790 47.600 193.930 ;
  RECT 88.270 192.790 88.520 193.930 ;
  RECT 129.190 192.790 129.440 193.930 ;
  RECT 170.110 192.790 170.360 193.930 ;
  RECT 211.030 192.790 211.280 193.930 ;
  RECT 251.950 192.790 252.200 193.930 ;
  RECT 292.870 192.790 293.120 193.930 ;
  RECT 333.790 192.790 334.040 193.930 ;
  RECT 374.710 192.790 374.960 193.930 ;
  RECT 415.630 192.790 415.880 193.930 ;
  RECT 456.550 192.790 456.800 193.930 ;
  RECT 497.470 192.790 497.720 193.930 ;
  RECT 538.390 192.790 538.640 193.930 ;
  RECT 579.310 192.790 579.560 193.930 ;
  RECT 620.230 192.790 620.480 193.930 ;
  RECT 661.150 192.790 661.400 193.930 ;
  RECT 702.070 192.790 702.320 193.930 ;
  RECT 742.990 192.790 743.240 193.930 ;
  RECT 783.910 192.790 784.160 193.930 ;
  RECT 824.830 192.790 825.080 193.930 ;
  RECT 865.750 192.790 866.000 193.930 ;
  RECT 906.670 192.790 906.920 193.930 ;
  RECT 947.590 192.790 947.840 193.930 ;
  RECT 988.510 192.790 988.760 193.930 ;
  RECT 1029.430 192.790 1029.680 193.930 ;
  RECT 1070.350 192.790 1070.600 193.930 ;
  RECT 1111.270 192.790 1111.520 193.930 ;
  RECT 1152.190 192.790 1152.440 193.930 ;
  RECT 1193.110 192.790 1193.360 193.930 ;
  RECT 1234.030 192.790 1234.280 193.930 ;
  RECT 1274.950 192.790 1275.200 193.930 ;
  RECT 2.000 193.930 2682.940 195.930 ;
  RECT 2.000 3.600 2682.940 5.600 ;
  RECT 2680.940 3.600 2682.940 195.930 ;
  RECT 2.000 3.600 4.000 195.930 ;
  LAYER ME3 ;
  RECT 5.420 7.020 2679.520 192.510 ;
  RECT 2682.940 3.600 2684.940 195.930 ;
  RECT 0.000 3.600 2.000 195.930 ;
  RECT 2.000 195.930 2682.940 197.930 ;
  RECT 2.000 1.600 2682.940 3.600 ;
  RECT 2680.940 187.000 2682.660 193.930 ;
  RECT 2680.940 64.930 2682.660 67.240 ;
  RECT 2680.940 44.080 2682.660 61.260 ;
  RECT 2680.940 39.620 2682.660 41.480 ;
  RECT 2680.940 29.870 2682.660 33.520 ;
  RECT 2680.940 24.270 2682.660 26.870 ;
  RECT 2680.940 18.130 2682.660 21.270 ;
  RECT 2680.940 5.600 2682.660 11.230 ;
  RECT 2.280 187.000 4.000 193.930 ;
  RECT 2.280 64.930 4.000 67.240 ;
  RECT 2.280 44.080 4.000 61.260 ;
  RECT 2.280 39.620 4.000 41.480 ;
  RECT 2.280 29.870 4.000 33.520 ;
  RECT 2.280 24.270 4.000 26.870 ;
  RECT 2.280 18.130 4.000 21.270 ;
  RECT 2.280 5.600 4.000 11.230 ;
  RECT 2638.020 193.930 2680.940 195.650 ;
  RECT 2597.100 193.930 2635.770 195.650 ;
  RECT 2556.180 193.930 2594.850 195.650 ;
  RECT 2515.260 193.930 2553.930 195.650 ;
  RECT 2474.340 193.930 2513.010 195.650 ;
  RECT 2433.420 193.930 2472.090 195.650 ;
  RECT 2392.500 193.930 2431.170 195.650 ;
  RECT 2351.580 193.930 2390.250 195.650 ;
  RECT 2310.660 193.930 2349.330 195.650 ;
  RECT 2269.740 193.930 2308.410 195.650 ;
  RECT 2228.820 193.930 2267.490 195.650 ;
  RECT 2187.900 193.930 2226.570 195.650 ;
  RECT 2146.980 193.930 2185.650 195.650 ;
  RECT 2106.060 193.930 2144.730 195.650 ;
  RECT 2065.140 193.930 2103.810 195.650 ;
  RECT 2024.220 193.930 2062.890 195.650 ;
  RECT 1983.300 193.930 2021.970 195.650 ;
  RECT 1942.380 193.930 1981.050 195.650 ;
  RECT 1901.460 193.930 1940.130 195.650 ;
  RECT 1860.540 193.930 1899.210 195.650 ;
  RECT 1819.620 193.930 1858.290 195.650 ;
  RECT 1778.700 193.930 1817.370 195.650 ;
  RECT 1737.780 193.930 1776.450 195.650 ;
  RECT 1696.860 193.930 1735.530 195.650 ;
  RECT 1655.940 193.930 1694.610 195.650 ;
  RECT 1615.020 193.930 1653.690 195.650 ;
  RECT 1574.100 193.930 1612.770 195.650 ;
  RECT 1533.180 193.930 1571.850 195.650 ;
  RECT 1492.260 193.930 1530.930 195.650 ;
  RECT 1451.340 193.930 1490.010 195.650 ;
  RECT 1410.420 193.930 1449.090 195.650 ;
  RECT 1369.500 193.930 1408.170 195.650 ;
  RECT 1350.760 193.930 1363.760 195.650 ;
  RECT 1339.630 193.930 1344.440 195.650 ;
  RECT 1329.920 193.930 1334.440 195.650 ;
  RECT 1324.580 193.930 1326.160 195.650 ;
  RECT 1276.770 193.930 1315.800 195.650 ;
  RECT 1235.850 193.930 1274.520 195.650 ;
  RECT 1194.930 193.930 1233.600 195.650 ;
  RECT 1154.010 193.930 1192.680 195.650 ;
  RECT 1113.090 193.930 1151.760 195.650 ;
  RECT 1072.170 193.930 1110.840 195.650 ;
  RECT 1031.250 193.930 1069.920 195.650 ;
  RECT 990.330 193.930 1029.000 195.650 ;
  RECT 949.410 193.930 988.080 195.650 ;
  RECT 908.490 193.930 947.160 195.650 ;
  RECT 867.570 193.930 906.240 195.650 ;
  RECT 826.650 193.930 865.320 195.650 ;
  RECT 785.730 193.930 824.400 195.650 ;
  RECT 744.810 193.930 783.480 195.650 ;
  RECT 703.890 193.930 742.560 195.650 ;
  RECT 662.970 193.930 701.640 195.650 ;
  RECT 622.050 193.930 660.720 195.650 ;
  RECT 581.130 193.930 619.800 195.650 ;
  RECT 540.210 193.930 578.880 195.650 ;
  RECT 499.290 193.930 537.960 195.650 ;
  RECT 458.370 193.930 497.040 195.650 ;
  RECT 417.450 193.930 456.120 195.650 ;
  RECT 376.530 193.930 415.200 195.650 ;
  RECT 335.610 193.930 374.280 195.650 ;
  RECT 294.690 193.930 333.360 195.650 ;
  RECT 253.770 193.930 292.440 195.650 ;
  RECT 212.850 193.930 251.520 195.650 ;
  RECT 171.930 193.930 210.600 195.650 ;
  RECT 131.010 193.930 169.680 195.650 ;
  RECT 90.090 193.930 128.760 195.650 ;
  RECT 49.170 193.930 87.840 195.650 ;
  RECT 4.000 193.930 46.920 195.650 ;
  RECT 2667.540 3.880 2677.380 5.600 ;
  RECT 2647.700 3.880 2657.540 5.600 ;
  RECT 2626.620 3.880 2637.700 5.600 ;
  RECT 2606.780 3.880 2616.620 5.600 ;
  RECT 2585.700 3.880 2596.780 5.600 ;
  RECT 2565.860 3.880 2575.700 5.600 ;
  RECT 2544.780 3.880 2555.860 5.600 ;
  RECT 2524.940 3.880 2534.780 5.600 ;
  RECT 2503.860 3.880 2514.940 5.600 ;
  RECT 2484.020 3.880 2493.860 5.600 ;
  RECT 2462.940 3.880 2474.020 5.600 ;
  RECT 2443.100 3.880 2452.940 5.600 ;
  RECT 2422.020 3.880 2433.100 5.600 ;
  RECT 2402.180 3.880 2412.020 5.600 ;
  RECT 2381.100 3.880 2392.180 5.600 ;
  RECT 2361.260 3.880 2371.100 5.600 ;
  RECT 2340.180 3.880 2351.260 5.600 ;
  RECT 2320.340 3.880 2330.180 5.600 ;
  RECT 2299.260 3.880 2310.340 5.600 ;
  RECT 2279.420 3.880 2289.260 5.600 ;
  RECT 2258.340 3.880 2269.420 5.600 ;
  RECT 2238.500 3.880 2248.340 5.600 ;
  RECT 2217.420 3.880 2228.500 5.600 ;
  RECT 2197.580 3.880 2207.420 5.600 ;
  RECT 2176.500 3.880 2187.580 5.600 ;
  RECT 2156.660 3.880 2166.500 5.600 ;
  RECT 2135.580 3.880 2146.660 5.600 ;
  RECT 2115.740 3.880 2125.580 5.600 ;
  RECT 2094.660 3.880 2105.740 5.600 ;
  RECT 2074.820 3.880 2084.660 5.600 ;
  RECT 2053.740 3.880 2064.820 5.600 ;
  RECT 2033.900 3.880 2043.740 5.600 ;
  RECT 2012.820 3.880 2023.900 5.600 ;
  RECT 1992.980 3.880 2002.820 5.600 ;
  RECT 1971.900 3.880 1982.980 5.600 ;
  RECT 1952.060 3.880 1961.900 5.600 ;
  RECT 1930.980 3.880 1942.060 5.600 ;
  RECT 1911.140 3.880 1920.980 5.600 ;
  RECT 1890.060 3.880 1901.140 5.600 ;
  RECT 1870.220 3.880 1880.060 5.600 ;
  RECT 1849.140 3.880 1860.220 5.600 ;
  RECT 1829.300 3.880 1839.140 5.600 ;
  RECT 1808.220 3.880 1819.300 5.600 ;
  RECT 1788.380 3.880 1798.220 5.600 ;
  RECT 1767.300 3.880 1778.380 5.600 ;
  RECT 1747.460 3.880 1757.300 5.600 ;
  RECT 1726.380 3.880 1737.460 5.600 ;
  RECT 1706.540 3.880 1716.380 5.600 ;
  RECT 1685.460 3.880 1696.540 5.600 ;
  RECT 1665.620 3.880 1675.460 5.600 ;
  RECT 1644.540 3.880 1655.620 5.600 ;
  RECT 1624.700 3.880 1634.540 5.600 ;
  RECT 1603.620 3.880 1614.700 5.600 ;
  RECT 1583.780 3.880 1593.620 5.600 ;
  RECT 1562.700 3.880 1573.780 5.600 ;
  RECT 1542.860 3.880 1552.700 5.600 ;
  RECT 1521.780 3.880 1532.860 5.600 ;
  RECT 1501.940 3.880 1511.780 5.600 ;
  RECT 1480.860 3.880 1491.940 5.600 ;
  RECT 1461.020 3.880 1470.860 5.600 ;
  RECT 1439.940 3.880 1451.020 5.600 ;
  RECT 1420.100 3.880 1429.940 5.600 ;
  RECT 1399.020 3.880 1410.100 5.600 ;
  RECT 1379.180 3.880 1389.020 5.600 ;
  RECT 1351.210 3.880 1369.180 5.600 ;
  RECT 1339.890 3.880 1343.290 5.600 ;
  RECT 1329.920 3.880 1334.440 5.600 ;
  RECT 1324.580 3.880 1326.160 5.600 ;
  RECT 1305.720 3.880 1316.820 5.600 ;
  RECT 1285.880 3.880 1295.720 5.600 ;
  RECT 1264.800 3.880 1275.880 5.600 ;
  RECT 1244.960 3.880 1254.800 5.600 ;
  RECT 1223.880 3.880 1234.960 5.600 ;
  RECT 1204.040 3.880 1213.880 5.600 ;
  RECT 1182.960 3.880 1194.040 5.600 ;
  RECT 1163.120 3.880 1172.960 5.600 ;
  RECT 1142.040 3.880 1153.120 5.600 ;
  RECT 1122.200 3.880 1132.040 5.600 ;
  RECT 1101.120 3.880 1112.200 5.600 ;
  RECT 1081.280 3.880 1091.120 5.600 ;
  RECT 1060.200 3.880 1071.280 5.600 ;
  RECT 1040.360 3.880 1050.200 5.600 ;
  RECT 1019.280 3.880 1030.360 5.600 ;
  RECT 999.440 3.880 1009.280 5.600 ;
  RECT 978.360 3.880 989.440 5.600 ;
  RECT 958.520 3.880 968.360 5.600 ;
  RECT 937.440 3.880 948.520 5.600 ;
  RECT 917.600 3.880 927.440 5.600 ;
  RECT 896.520 3.880 907.600 5.600 ;
  RECT 876.680 3.880 886.520 5.600 ;
  RECT 855.600 3.880 866.680 5.600 ;
  RECT 835.760 3.880 845.600 5.600 ;
  RECT 814.680 3.880 825.760 5.600 ;
  RECT 794.840 3.880 804.680 5.600 ;
  RECT 773.760 3.880 784.840 5.600 ;
  RECT 753.920 3.880 763.760 5.600 ;
  RECT 732.840 3.880 743.920 5.600 ;
  RECT 713.000 3.880 722.840 5.600 ;
  RECT 691.920 3.880 703.000 5.600 ;
  RECT 672.080 3.880 681.920 5.600 ;
  RECT 651.000 3.880 662.080 5.600 ;
  RECT 631.160 3.880 641.000 5.600 ;
  RECT 610.080 3.880 621.160 5.600 ;
  RECT 590.240 3.880 600.080 5.600 ;
  RECT 569.160 3.880 580.240 5.600 ;
  RECT 549.320 3.880 559.160 5.600 ;
  RECT 528.240 3.880 539.320 5.600 ;
  RECT 508.400 3.880 518.240 5.600 ;
  RECT 487.320 3.880 498.400 5.600 ;
  RECT 467.480 3.880 477.320 5.600 ;
  RECT 446.400 3.880 457.480 5.600 ;
  RECT 426.560 3.880 436.400 5.600 ;
  RECT 405.480 3.880 416.560 5.600 ;
  RECT 385.640 3.880 395.480 5.600 ;
  RECT 364.560 3.880 375.640 5.600 ;
  RECT 344.720 3.880 354.560 5.600 ;
  RECT 323.640 3.880 334.720 5.600 ;
  RECT 303.800 3.880 313.640 5.600 ;
  RECT 282.720 3.880 293.800 5.600 ;
  RECT 262.880 3.880 272.720 5.600 ;
  RECT 241.800 3.880 252.880 5.600 ;
  RECT 221.960 3.880 231.800 5.600 ;
  RECT 200.880 3.880 211.960 5.600 ;
  RECT 181.040 3.880 190.880 5.600 ;
  RECT 159.960 3.880 171.040 5.600 ;
  RECT 140.120 3.880 149.960 5.600 ;
  RECT 119.040 3.880 130.120 5.600 ;
  RECT 99.200 3.880 109.040 5.600 ;
  RECT 78.120 3.880 89.200 5.600 ;
  RECT 58.280 3.880 68.120 5.600 ;
  RECT 37.200 3.880 48.280 5.600 ;
  RECT 17.360 3.880 27.200 5.600 ;
  RECT 2.280 193.930 4.000 195.650 ;
  RECT 0.000 195.930 2.000 197.930 ;
  RECT 2680.940 3.880 2682.660 5.600 ;
  RECT 2682.940 1.600 2684.940 3.600 ;
  RECT 2680.940 193.930 2682.660 195.650 ;
  RECT 2682.940 195.930 2684.940 197.930 ;
  RECT 2.280 3.880 4.000 5.600 ;
  RECT 0.000 1.600 2.000 3.600 ;
  RECT 2672.800 0.000 2673.600 1.000 ;
  RECT 2658.400 0.000 2659.200 1.000 ;
  RECT 2653.200 0.000 2654.000 1.000 ;
  RECT 2638.400 0.000 2639.200 1.000 ;
  RECT 2632.000 0.000 2632.800 1.000 ;
  RECT 2617.600 0.000 2618.400 1.000 ;
  RECT 2612.400 0.000 2613.200 1.000 ;
  RECT 2597.600 0.000 2598.400 1.000 ;
  RECT 2591.200 0.000 2592.000 1.000 ;
  RECT 2576.400 0.000 2577.200 1.000 ;
  RECT 2571.200 0.000 2572.000 1.000 ;
  RECT 2556.800 0.000 2557.600 1.000 ;
  RECT 2550.400 0.000 2551.200 1.000 ;
  RECT 2535.600 0.000 2536.400 1.000 ;
  RECT 2530.400 0.000 2531.200 1.000 ;
  RECT 2515.600 0.000 2516.400 1.000 ;
  RECT 2509.200 0.000 2510.000 1.000 ;
  RECT 2494.800 0.000 2495.600 1.000 ;
  RECT 2489.600 0.000 2490.400 1.000 ;
  RECT 2474.800 0.000 2475.600 1.000 ;
  RECT 2468.400 0.000 2469.200 1.000 ;
  RECT 2453.600 0.000 2454.400 1.000 ;
  RECT 2448.400 0.000 2449.200 1.000 ;
  RECT 2434.000 0.000 2434.800 1.000 ;
  RECT 2427.600 0.000 2428.400 1.000 ;
  RECT 2412.800 0.000 2413.600 1.000 ;
  RECT 2407.600 0.000 2408.400 1.000 ;
  RECT 2392.800 0.000 2393.600 1.000 ;
  RECT 2386.400 0.000 2387.200 1.000 ;
  RECT 2372.000 0.000 2372.800 1.000 ;
  RECT 2366.800 0.000 2367.600 1.000 ;
  RECT 2353.600 0.000 2354.400 1.000 ;
  RECT 2352.000 0.000 2352.800 1.000 ;
  RECT 2345.600 0.000 2346.400 1.000 ;
  RECT 2330.800 0.000 2331.600 1.000 ;
  RECT 2325.600 0.000 2326.400 1.000 ;
  RECT 2311.200 0.000 2312.000 1.000 ;
  RECT 2304.800 0.000 2305.600 1.000 ;
  RECT 2290.000 0.000 2290.800 1.000 ;
  RECT 2284.800 0.000 2285.600 1.000 ;
  RECT 2270.400 0.000 2271.200 1.000 ;
  RECT 2263.600 0.000 2264.400 1.000 ;
  RECT 2249.200 0.000 2250.000 1.000 ;
  RECT 2244.000 0.000 2244.800 1.000 ;
  RECT 2229.200 0.000 2230.000 1.000 ;
  RECT 2222.800 0.000 2223.600 1.000 ;
  RECT 2208.400 0.000 2209.200 1.000 ;
  RECT 2203.200 0.000 2204.000 1.000 ;
  RECT 2188.400 0.000 2189.200 1.000 ;
  RECT 2182.000 0.000 2182.800 1.000 ;
  RECT 2167.200 0.000 2168.000 1.000 ;
  RECT 2162.000 0.000 2162.800 1.000 ;
  RECT 2147.600 0.000 2148.400 1.000 ;
  RECT 2141.200 0.000 2142.000 1.000 ;
  RECT 2126.400 0.000 2127.200 1.000 ;
  RECT 2121.200 0.000 2122.000 1.000 ;
  RECT 2106.400 0.000 2107.200 1.000 ;
  RECT 2100.000 0.000 2100.800 1.000 ;
  RECT 2085.600 0.000 2086.400 1.000 ;
  RECT 2080.400 0.000 2081.200 1.000 ;
  RECT 2065.600 0.000 2066.400 1.000 ;
  RECT 2059.200 0.000 2060.000 1.000 ;
  RECT 2044.400 0.000 2045.200 1.000 ;
  RECT 2039.200 0.000 2040.000 1.000 ;
  RECT 2026.400 0.000 2027.200 1.000 ;
  RECT 2024.800 0.000 2025.600 1.000 ;
  RECT 2018.400 0.000 2019.200 1.000 ;
  RECT 2003.600 0.000 2004.400 1.000 ;
  RECT 1998.400 0.000 1999.200 1.000 ;
  RECT 1983.600 0.000 1984.400 1.000 ;
  RECT 1977.200 0.000 1978.000 1.000 ;
  RECT 1962.800 0.000 1963.600 1.000 ;
  RECT 1957.600 0.000 1958.400 1.000 ;
  RECT 1942.800 0.000 1943.600 1.000 ;
  RECT 1936.400 0.000 1937.200 1.000 ;
  RECT 1921.600 0.000 1922.400 1.000 ;
  RECT 1916.400 0.000 1917.200 1.000 ;
  RECT 1902.000 0.000 1902.800 1.000 ;
  RECT 1895.600 0.000 1896.400 1.000 ;
  RECT 1880.800 0.000 1881.600 1.000 ;
  RECT 1875.600 0.000 1876.400 1.000 ;
  RECT 1861.200 0.000 1862.000 1.000 ;
  RECT 1854.400 0.000 1855.200 1.000 ;
  RECT 1840.000 0.000 1840.800 1.000 ;
  RECT 1834.800 0.000 1835.600 1.000 ;
  RECT 1820.000 0.000 1820.800 1.000 ;
  RECT 1813.600 0.000 1814.400 1.000 ;
  RECT 1799.200 0.000 1800.000 1.000 ;
  RECT 1794.000 0.000 1794.800 1.000 ;
  RECT 1779.200 0.000 1780.000 1.000 ;
  RECT 1772.800 0.000 1773.600 1.000 ;
  RECT 1758.000 0.000 1758.800 1.000 ;
  RECT 1752.800 0.000 1753.600 1.000 ;
  RECT 1738.400 0.000 1739.200 1.000 ;
  RECT 1732.000 0.000 1732.800 1.000 ;
  RECT 1717.200 0.000 1718.000 1.000 ;
  RECT 1712.000 0.000 1712.800 1.000 ;
  RECT 1699.200 0.000 1700.000 1.000 ;
  RECT 1697.200 0.000 1698.000 1.000 ;
  RECT 1690.800 0.000 1691.600 1.000 ;
  RECT 1676.400 0.000 1677.200 1.000 ;
  RECT 1671.200 0.000 1672.000 1.000 ;
  RECT 1656.400 0.000 1657.200 1.000 ;
  RECT 1650.000 0.000 1650.800 1.000 ;
  RECT 1635.200 0.000 1636.000 1.000 ;
  RECT 1630.000 0.000 1630.800 1.000 ;
  RECT 1615.600 0.000 1616.400 1.000 ;
  RECT 1609.200 0.000 1610.000 1.000 ;
  RECT 1594.400 0.000 1595.200 1.000 ;
  RECT 1589.200 0.000 1590.000 1.000 ;
  RECT 1574.400 0.000 1575.200 1.000 ;
  RECT 1568.000 0.000 1568.800 1.000 ;
  RECT 1553.600 0.000 1554.400 1.000 ;
  RECT 1548.400 0.000 1549.200 1.000 ;
  RECT 1533.600 0.000 1534.400 1.000 ;
  RECT 1527.200 0.000 1528.000 1.000 ;
  RECT 1512.400 0.000 1513.200 1.000 ;
  RECT 1507.200 0.000 1508.000 1.000 ;
  RECT 1492.800 0.000 1493.600 1.000 ;
  RECT 1486.400 0.000 1487.200 1.000 ;
  RECT 1471.600 0.000 1472.400 1.000 ;
  RECT 1466.400 0.000 1467.200 1.000 ;
  RECT 1452.000 0.000 1452.800 1.000 ;
  RECT 1445.200 0.000 1446.000 1.000 ;
  RECT 1430.800 0.000 1431.600 1.000 ;
  RECT 1425.600 0.000 1426.400 1.000 ;
  RECT 1410.800 0.000 1411.600 1.000 ;
  RECT 1404.400 0.000 1405.200 1.000 ;
  RECT 1390.000 0.000 1390.800 1.000 ;
  RECT 1384.800 0.000 1385.600 1.000 ;
  RECT 1371.600 0.000 1372.400 1.000 ;
  RECT 1370.000 0.000 1370.800 1.000 ;
  RECT 1349.200 0.000 1350.000 1.000 ;
  RECT 1348.000 0.000 1348.800 1.000 ;
  RECT 1346.800 0.000 1347.600 1.000 ;
  RECT 1345.600 0.000 1346.400 1.000 ;
  RECT 1344.400 0.000 1345.200 1.000 ;
  RECT 1343.200 0.000 1344.000 1.000 ;
  RECT 1337.200 0.000 1338.000 1.000 ;
  RECT 1330.000 0.000 1330.800 1.000 ;
  RECT 1327.200 0.000 1328.000 1.000 ;
  RECT 1324.400 0.000 1325.200 1.000 ;
  RECT 1322.000 0.000 1322.800 1.000 ;
  RECT 1320.400 0.000 1321.200 1.000 ;
  RECT 1318.000 0.000 1318.800 1.000 ;
  RECT 1311.200 0.000 1312.000 1.000 ;
  RECT 1296.400 0.000 1297.200 1.000 ;
  RECT 1291.200 0.000 1292.000 1.000 ;
  RECT 1276.800 0.000 1277.600 1.000 ;
  RECT 1270.400 0.000 1271.200 1.000 ;
  RECT 1255.600 0.000 1256.400 1.000 ;
  RECT 1250.400 0.000 1251.200 1.000 ;
  RECT 1235.600 0.000 1236.400 1.000 ;
  RECT 1229.200 0.000 1230.000 1.000 ;
  RECT 1214.800 0.000 1215.600 1.000 ;
  RECT 1209.600 0.000 1210.400 1.000 ;
  RECT 1194.800 0.000 1195.600 1.000 ;
  RECT 1188.400 0.000 1189.200 1.000 ;
  RECT 1173.600 0.000 1174.400 1.000 ;
  RECT 1168.400 0.000 1169.200 1.000 ;
  RECT 1154.000 0.000 1154.800 1.000 ;
  RECT 1147.600 0.000 1148.400 1.000 ;
  RECT 1132.800 0.000 1133.600 1.000 ;
  RECT 1127.600 0.000 1128.400 1.000 ;
  RECT 1113.200 0.000 1114.000 1.000 ;
  RECT 1106.400 0.000 1107.200 1.000 ;
  RECT 1092.000 0.000 1092.800 1.000 ;
  RECT 1086.800 0.000 1087.600 1.000 ;
  RECT 1072.000 0.000 1072.800 1.000 ;
  RECT 1065.600 0.000 1066.400 1.000 ;
  RECT 1051.200 0.000 1052.000 1.000 ;
  RECT 1045.600 0.000 1046.400 1.000 ;
  RECT 1031.200 0.000 1032.000 1.000 ;
  RECT 1024.800 0.000 1025.600 1.000 ;
  RECT 1010.000 0.000 1010.800 1.000 ;
  RECT 1004.800 0.000 1005.600 1.000 ;
  RECT 992.000 0.000 992.800 1.000 ;
  RECT 990.400 0.000 991.200 1.000 ;
  RECT 983.600 0.000 984.400 1.000 ;
  RECT 969.200 0.000 970.000 1.000 ;
  RECT 964.000 0.000 964.800 1.000 ;
  RECT 949.200 0.000 950.000 1.000 ;
  RECT 942.800 0.000 943.600 1.000 ;
  RECT 928.400 0.000 929.200 1.000 ;
  RECT 923.200 0.000 924.000 1.000 ;
  RECT 908.400 0.000 909.200 1.000 ;
  RECT 902.000 0.000 902.800 1.000 ;
  RECT 887.200 0.000 888.000 1.000 ;
  RECT 882.000 0.000 882.800 1.000 ;
  RECT 867.600 0.000 868.400 1.000 ;
  RECT 861.200 0.000 862.000 1.000 ;
  RECT 846.400 0.000 847.200 1.000 ;
  RECT 841.200 0.000 842.000 1.000 ;
  RECT 826.400 0.000 827.200 1.000 ;
  RECT 820.000 0.000 820.800 1.000 ;
  RECT 805.600 0.000 806.400 1.000 ;
  RECT 800.400 0.000 801.200 1.000 ;
  RECT 785.600 0.000 786.400 1.000 ;
  RECT 779.200 0.000 780.000 1.000 ;
  RECT 764.400 0.000 765.200 1.000 ;
  RECT 759.200 0.000 760.000 1.000 ;
  RECT 744.800 0.000 745.600 1.000 ;
  RECT 738.400 0.000 739.200 1.000 ;
  RECT 723.600 0.000 724.400 1.000 ;
  RECT 718.400 0.000 719.200 1.000 ;
  RECT 704.000 0.000 704.800 1.000 ;
  RECT 697.200 0.000 698.000 1.000 ;
  RECT 682.800 0.000 683.600 1.000 ;
  RECT 677.600 0.000 678.400 1.000 ;
  RECT 664.800 0.000 665.600 1.000 ;
  RECT 662.800 0.000 663.600 1.000 ;
  RECT 656.400 0.000 657.200 1.000 ;
  RECT 642.000 0.000 642.800 1.000 ;
  RECT 636.400 0.000 637.200 1.000 ;
  RECT 622.000 0.000 622.800 1.000 ;
  RECT 615.600 0.000 616.400 1.000 ;
  RECT 600.800 0.000 601.600 1.000 ;
  RECT 595.600 0.000 596.400 1.000 ;
  RECT 581.200 0.000 582.000 1.000 ;
  RECT 574.400 0.000 575.200 1.000 ;
  RECT 560.000 0.000 560.800 1.000 ;
  RECT 554.800 0.000 555.600 1.000 ;
  RECT 540.000 0.000 540.800 1.000 ;
  RECT 533.600 0.000 534.400 1.000 ;
  RECT 519.200 0.000 520.000 1.000 ;
  RECT 514.000 0.000 514.800 1.000 ;
  RECT 499.200 0.000 500.000 1.000 ;
  RECT 492.800 0.000 493.600 1.000 ;
  RECT 478.000 0.000 478.800 1.000 ;
  RECT 472.800 0.000 473.600 1.000 ;
  RECT 458.400 0.000 459.200 1.000 ;
  RECT 452.000 0.000 452.800 1.000 ;
  RECT 437.200 0.000 438.000 1.000 ;
  RECT 432.000 0.000 432.800 1.000 ;
  RECT 417.200 0.000 418.000 1.000 ;
  RECT 410.800 0.000 411.600 1.000 ;
  RECT 396.400 0.000 397.200 1.000 ;
  RECT 391.200 0.000 392.000 1.000 ;
  RECT 376.400 0.000 377.200 1.000 ;
  RECT 370.000 0.000 370.800 1.000 ;
  RECT 355.200 0.000 356.000 1.000 ;
  RECT 350.000 0.000 350.800 1.000 ;
  RECT 337.200 0.000 338.000 1.000 ;
  RECT 335.600 0.000 336.400 1.000 ;
  RECT 329.200 0.000 330.000 1.000 ;
  RECT 314.400 0.000 315.200 1.000 ;
  RECT 309.200 0.000 310.000 1.000 ;
  RECT 294.800 0.000 295.600 1.000 ;
  RECT 288.000 0.000 288.800 1.000 ;
  RECT 273.600 0.000 274.400 1.000 ;
  RECT 268.400 0.000 269.200 1.000 ;
  RECT 253.600 0.000 254.400 1.000 ;
  RECT 247.200 0.000 248.000 1.000 ;
  RECT 232.800 0.000 233.600 1.000 ;
  RECT 227.200 0.000 228.000 1.000 ;
  RECT 212.800 0.000 213.600 1.000 ;
  RECT 206.400 0.000 207.200 1.000 ;
  RECT 191.600 0.000 192.400 1.000 ;
  RECT 186.400 0.000 187.200 1.000 ;
  RECT 172.000 0.000 172.800 1.000 ;
  RECT 165.200 0.000 166.000 1.000 ;
  RECT 150.800 0.000 151.600 1.000 ;
  RECT 145.600 0.000 146.400 1.000 ;
  RECT 130.800 0.000 131.600 1.000 ;
  RECT 124.400 0.000 125.200 1.000 ;
  RECT 110.000 0.000 110.800 1.000 ;
  RECT 104.800 0.000 105.600 1.000 ;
  RECT 90.000 0.000 90.800 1.000 ;
  RECT 83.600 0.000 84.400 1.000 ;
  RECT 68.800 0.000 69.600 1.000 ;
  RECT 63.600 0.000 64.400 1.000 ;
  RECT 49.200 0.000 50.000 1.000 ;
  RECT 42.800 0.000 43.600 1.000 ;
  RECT 28.000 0.000 28.800 1.000 ;
  RECT 22.800 0.000 23.600 1.000 ;
  RECT 10.000 0.000 10.800 1.000 ;
  RECT 8.000 0.000 8.800 1.000 ;
  RECT 2679.520 62.260 2682.940 63.930 ;
  RECT 2679.520 22.270 2682.940 23.270 ;
  RECT 2679.520 16.130 2682.940 17.130 ;
  RECT 2679.520 12.230 2682.940 13.230 ;
  RECT 2679.520 27.870 2682.940 28.870 ;
  RECT 2679.520 42.480 2682.940 43.080 ;
  RECT 2679.520 37.620 2682.940 38.620 ;
  RECT 2679.520 34.520 2682.940 36.020 ;
  RECT 2679.800 9.570 2680.660 11.170 ;
  RECT 2679.800 14.200 2680.660 15.200 ;
  RECT 2679.800 18.730 2680.660 19.730 ;
  RECT 2679.800 21.230 2680.660 22.070 ;
  RECT 2679.800 24.170 2680.660 25.170 ;
  RECT 2679.800 36.320 2680.660 37.320 ;
  RECT 2679.800 39.480 2680.660 40.080 ;
  RECT 2679.800 45.560 2680.660 46.160 ;
  RECT 2679.800 57.100 2680.660 61.420 ;
  RECT 2678.380 3.600 2679.520 6.740 ;
  RECT 1370.180 3.600 1378.180 6.740 ;
  RECT 1390.020 3.600 1398.020 6.740 ;
  RECT 1411.100 3.600 1419.100 6.740 ;
  RECT 1430.940 3.600 1438.940 6.740 ;
  RECT 1452.020 3.600 1460.020 6.740 ;
  RECT 1471.860 3.600 1479.860 6.740 ;
  RECT 1492.940 3.600 1500.940 6.740 ;
  RECT 1512.780 3.600 1520.780 6.740 ;
  RECT 1533.860 3.600 1541.860 6.740 ;
  RECT 1553.700 3.600 1561.700 6.740 ;
  RECT 1574.780 3.600 1582.780 6.740 ;
  RECT 1594.620 3.600 1602.620 6.740 ;
  RECT 1615.700 3.600 1623.700 6.740 ;
  RECT 1635.540 3.600 1643.540 6.740 ;
  RECT 1656.620 3.600 1664.620 6.740 ;
  RECT 1676.460 3.600 1684.460 6.740 ;
  RECT 1697.540 3.600 1705.540 6.740 ;
  RECT 1717.380 3.600 1725.380 6.740 ;
  RECT 1738.460 3.600 1746.460 6.740 ;
  RECT 1758.300 3.600 1766.300 6.740 ;
  RECT 1779.380 3.600 1787.380 6.740 ;
  RECT 1799.220 3.600 1807.220 6.740 ;
  RECT 1820.300 3.600 1828.300 6.740 ;
  RECT 1840.140 3.600 1848.140 6.740 ;
  RECT 1861.220 3.600 1869.220 6.740 ;
  RECT 1881.060 3.600 1889.060 6.740 ;
  RECT 1902.140 3.600 1910.140 6.740 ;
  RECT 1921.980 3.600 1929.980 6.740 ;
  RECT 1943.060 3.600 1951.060 6.740 ;
  RECT 1962.900 3.600 1970.900 6.740 ;
  RECT 1983.980 3.600 1991.980 6.740 ;
  RECT 2003.820 3.600 2011.820 6.740 ;
  RECT 2024.900 3.600 2032.900 6.740 ;
  RECT 2044.740 3.600 2052.740 6.740 ;
  RECT 2065.820 3.600 2073.820 6.740 ;
  RECT 2085.660 3.600 2093.660 6.740 ;
  RECT 2106.740 3.600 2114.740 6.740 ;
  RECT 2126.580 3.600 2134.580 6.740 ;
  RECT 2147.660 3.600 2155.660 6.740 ;
  RECT 2167.500 3.600 2175.500 6.740 ;
  RECT 2188.580 3.600 2196.580 6.740 ;
  RECT 2208.420 3.600 2216.420 6.740 ;
  RECT 2229.500 3.600 2237.500 6.740 ;
  RECT 2249.340 3.600 2257.340 6.740 ;
  RECT 2270.420 3.600 2278.420 6.740 ;
  RECT 2290.260 3.600 2298.260 6.740 ;
  RECT 2311.340 3.600 2319.340 6.740 ;
  RECT 2331.180 3.600 2339.180 6.740 ;
  RECT 2352.260 3.600 2360.260 6.740 ;
  RECT 2372.100 3.600 2380.100 6.740 ;
  RECT 2393.180 3.600 2401.180 6.740 ;
  RECT 2413.020 3.600 2421.020 6.740 ;
  RECT 2434.100 3.600 2442.100 6.740 ;
  RECT 2453.940 3.600 2461.940 6.740 ;
  RECT 2475.020 3.600 2483.020 6.740 ;
  RECT 2494.860 3.600 2502.860 6.740 ;
  RECT 2515.940 3.600 2523.940 6.740 ;
  RECT 2535.780 3.600 2543.780 6.740 ;
  RECT 2556.860 3.600 2564.860 6.740 ;
  RECT 2576.700 3.600 2584.700 6.740 ;
  RECT 2597.780 3.600 2605.780 6.740 ;
  RECT 2617.620 3.600 2625.620 6.740 ;
  RECT 2638.700 3.600 2646.700 6.740 ;
  RECT 2658.540 3.600 2666.540 6.740 ;
  RECT 1335.440 3.600 1338.890 6.740 ;
  RECT 1344.290 3.600 1350.210 6.740 ;
  RECT 1327.160 3.600 1328.920 6.740 ;
  RECT 1321.820 3.600 1323.580 6.740 ;
  RECT 1317.820 3.600 1319.580 6.740 ;
  RECT 4.280 57.100 5.140 61.420 ;
  RECT 4.280 45.560 5.140 46.160 ;
  RECT 4.280 39.480 5.140 40.080 ;
  RECT 4.280 36.320 5.140 37.320 ;
  RECT 4.280 24.170 5.140 25.170 ;
  RECT 4.280 21.230 5.140 22.070 ;
  RECT 4.280 18.730 5.140 19.730 ;
  RECT 4.280 14.200 5.140 15.200 ;
  RECT 4.280 9.570 5.140 11.170 ;
  RECT 2.000 34.520 5.420 36.020 ;
  RECT 2.000 37.620 5.420 38.620 ;
  RECT 2.000 42.480 5.420 43.080 ;
  RECT 2.000 27.870 5.420 28.870 ;
  RECT 2.000 12.230 5.420 13.230 ;
  RECT 2.000 16.130 5.420 17.130 ;
  RECT 2.000 22.270 5.420 23.270 ;
  RECT 2.000 62.260 5.420 63.930 ;
  RECT 5.420 3.600 6.560 6.740 ;
  RECT 8.360 3.600 16.360 6.740 ;
  RECT 28.200 3.600 36.200 6.740 ;
  RECT 49.280 3.600 57.280 6.740 ;
  RECT 69.120 3.600 77.120 6.740 ;
  RECT 90.200 3.600 98.200 6.740 ;
  RECT 110.040 3.600 118.040 6.740 ;
  RECT 131.120 3.600 139.120 6.740 ;
  RECT 150.960 3.600 158.960 6.740 ;
  RECT 172.040 3.600 180.040 6.740 ;
  RECT 191.880 3.600 199.880 6.740 ;
  RECT 212.960 3.600 220.960 6.740 ;
  RECT 232.800 3.600 240.800 6.740 ;
  RECT 253.880 3.600 261.880 6.740 ;
  RECT 273.720 3.600 281.720 6.740 ;
  RECT 294.800 3.600 302.800 6.740 ;
  RECT 314.640 3.600 322.640 6.740 ;
  RECT 335.720 3.600 343.720 6.740 ;
  RECT 355.560 3.600 363.560 6.740 ;
  RECT 376.640 3.600 384.640 6.740 ;
  RECT 396.480 3.600 404.480 6.740 ;
  RECT 417.560 3.600 425.560 6.740 ;
  RECT 437.400 3.600 445.400 6.740 ;
  RECT 458.480 3.600 466.480 6.740 ;
  RECT 478.320 3.600 486.320 6.740 ;
  RECT 499.400 3.600 507.400 6.740 ;
  RECT 519.240 3.600 527.240 6.740 ;
  RECT 540.320 3.600 548.320 6.740 ;
  RECT 560.160 3.600 568.160 6.740 ;
  RECT 581.240 3.600 589.240 6.740 ;
  RECT 601.080 3.600 609.080 6.740 ;
  RECT 622.160 3.600 630.160 6.740 ;
  RECT 642.000 3.600 650.000 6.740 ;
  RECT 663.080 3.600 671.080 6.740 ;
  RECT 682.920 3.600 690.920 6.740 ;
  RECT 704.000 3.600 712.000 6.740 ;
  RECT 723.840 3.600 731.840 6.740 ;
  RECT 744.920 3.600 752.920 6.740 ;
  RECT 764.760 3.600 772.760 6.740 ;
  RECT 785.840 3.600 793.840 6.740 ;
  RECT 805.680 3.600 813.680 6.740 ;
  RECT 826.760 3.600 834.760 6.740 ;
  RECT 846.600 3.600 854.600 6.740 ;
  RECT 867.680 3.600 875.680 6.740 ;
  RECT 887.520 3.600 895.520 6.740 ;
  RECT 908.600 3.600 916.600 6.740 ;
  RECT 928.440 3.600 936.440 6.740 ;
  RECT 949.520 3.600 957.520 6.740 ;
  RECT 969.360 3.600 977.360 6.740 ;
  RECT 990.440 3.600 998.440 6.740 ;
  RECT 1010.280 3.600 1018.280 6.740 ;
  RECT 1031.360 3.600 1039.360 6.740 ;
  RECT 1051.200 3.600 1059.200 6.740 ;
  RECT 1072.280 3.600 1080.280 6.740 ;
  RECT 1092.120 3.600 1100.120 6.740 ;
  RECT 1113.200 3.600 1121.200 6.740 ;
  RECT 1133.040 3.600 1141.040 6.740 ;
  RECT 1154.120 3.600 1162.120 6.740 ;
  RECT 1173.960 3.600 1181.960 6.740 ;
  RECT 1195.040 3.600 1203.040 6.740 ;
  RECT 1214.880 3.600 1222.880 6.740 ;
  RECT 1235.960 3.600 1243.960 6.740 ;
  RECT 1255.800 3.600 1263.800 6.740 ;
  RECT 1276.880 3.600 1284.880 6.740 ;
  RECT 1296.720 3.600 1304.720 6.740 ;
  RECT 2679.800 191.940 2680.660 192.320 ;
  RECT 2679.800 184.020 2680.660 184.300 ;
  RECT 2679.520 184.800 2682.940 186.000 ;
  RECT 2679.520 182.320 2682.940 183.520 ;
  RECT 2679.800 180.340 2680.660 180.620 ;
  RECT 2679.520 181.120 2682.940 182.320 ;
  RECT 2679.520 178.640 2682.940 179.840 ;
  RECT 2679.800 176.660 2680.660 176.940 ;
  RECT 2679.520 177.440 2682.940 178.640 ;
  RECT 2679.520 174.960 2682.940 176.160 ;
  RECT 2679.800 172.980 2680.660 173.260 ;
  RECT 2679.520 173.760 2682.940 174.960 ;
  RECT 2679.520 171.280 2682.940 172.480 ;
  RECT 2679.800 169.300 2680.660 169.580 ;
  RECT 2679.520 170.080 2682.940 171.280 ;
  RECT 2679.520 167.600 2682.940 168.800 ;
  RECT 2679.800 165.620 2680.660 165.900 ;
  RECT 2679.520 166.400 2682.940 167.600 ;
  RECT 2679.520 163.920 2682.940 165.120 ;
  RECT 2679.800 161.940 2680.660 162.220 ;
  RECT 2679.520 162.720 2682.940 163.920 ;
  RECT 2679.520 160.240 2682.940 161.440 ;
  RECT 2679.800 158.260 2680.660 158.540 ;
  RECT 2679.520 159.040 2682.940 160.240 ;
  RECT 2679.520 156.560 2682.940 157.760 ;
  RECT 2679.800 154.580 2680.660 154.860 ;
  RECT 2679.520 155.360 2682.940 156.560 ;
  RECT 2679.520 152.880 2682.940 154.080 ;
  RECT 2679.800 150.900 2680.660 151.180 ;
  RECT 2679.520 151.680 2682.940 152.880 ;
  RECT 2679.520 149.200 2682.940 150.400 ;
  RECT 2679.800 147.220 2680.660 147.500 ;
  RECT 2679.520 148.000 2682.940 149.200 ;
  RECT 2679.520 145.520 2682.940 146.720 ;
  RECT 2679.800 143.540 2680.660 143.820 ;
  RECT 2679.520 144.320 2682.940 145.520 ;
  RECT 2679.520 141.840 2682.940 143.040 ;
  RECT 2679.800 139.860 2680.660 140.140 ;
  RECT 2679.520 140.640 2682.940 141.840 ;
  RECT 2679.520 138.160 2682.940 139.360 ;
  RECT 2679.800 136.180 2680.660 136.460 ;
  RECT 2679.520 136.960 2682.940 138.160 ;
  RECT 2679.520 134.480 2682.940 135.680 ;
  RECT 2679.800 132.500 2680.660 132.780 ;
  RECT 2679.520 133.280 2682.940 134.480 ;
  RECT 2679.520 130.800 2682.940 132.000 ;
  RECT 2679.800 128.820 2680.660 129.100 ;
  RECT 2679.520 129.600 2682.940 130.800 ;
  RECT 2679.520 127.120 2682.940 128.320 ;
  RECT 2679.800 125.140 2680.660 125.420 ;
  RECT 2679.520 125.920 2682.940 127.120 ;
  RECT 2679.520 123.440 2682.940 124.640 ;
  RECT 2679.800 121.460 2680.660 121.740 ;
  RECT 2679.520 122.240 2682.940 123.440 ;
  RECT 2679.520 119.760 2682.940 120.960 ;
  RECT 2679.800 117.780 2680.660 118.060 ;
  RECT 2679.520 118.560 2682.940 119.760 ;
  RECT 2679.520 116.080 2682.940 117.280 ;
  RECT 2679.800 114.100 2680.660 114.380 ;
  RECT 2679.520 114.880 2682.940 116.080 ;
  RECT 2679.520 112.400 2682.940 113.600 ;
  RECT 2679.800 110.420 2680.660 110.700 ;
  RECT 2679.520 111.200 2682.940 112.400 ;
  RECT 2679.520 108.720 2682.940 109.920 ;
  RECT 2679.800 106.740 2680.660 107.020 ;
  RECT 2679.520 107.520 2682.940 108.720 ;
  RECT 2679.520 105.040 2682.940 106.240 ;
  RECT 2679.800 103.060 2680.660 103.340 ;
  RECT 2679.520 103.840 2682.940 105.040 ;
  RECT 2679.520 101.360 2682.940 102.560 ;
  RECT 2679.800 99.380 2680.660 99.660 ;
  RECT 2679.520 100.160 2682.940 101.360 ;
  RECT 2679.520 97.680 2682.940 98.880 ;
  RECT 2679.800 95.700 2680.660 95.980 ;
  RECT 2679.520 96.480 2682.940 97.680 ;
  RECT 2679.520 94.000 2682.940 95.200 ;
  RECT 2679.800 92.020 2680.660 92.300 ;
  RECT 2679.520 92.800 2682.940 94.000 ;
  RECT 2679.520 90.320 2682.940 91.520 ;
  RECT 2679.800 88.340 2680.660 88.620 ;
  RECT 2679.520 89.120 2682.940 90.320 ;
  RECT 2679.520 86.640 2682.940 87.840 ;
  RECT 2679.800 84.660 2680.660 84.940 ;
  RECT 2679.520 85.440 2682.940 86.640 ;
  RECT 2679.520 82.960 2682.940 84.160 ;
  RECT 2679.800 80.980 2680.660 81.260 ;
  RECT 2679.520 81.760 2682.940 82.960 ;
  RECT 2679.520 79.280 2682.940 80.480 ;
  RECT 2679.800 77.300 2680.660 77.580 ;
  RECT 2679.520 78.080 2682.940 79.280 ;
  RECT 2679.520 75.600 2682.940 76.800 ;
  RECT 2679.800 73.620 2680.660 73.900 ;
  RECT 2679.520 74.400 2682.940 75.600 ;
  RECT 2679.520 71.920 2682.940 73.120 ;
  RECT 2679.800 69.940 2680.660 70.220 ;
  RECT 2679.520 70.720 2682.940 71.920 ;
  RECT 2679.520 68.240 2682.940 69.440 ;
  RECT 2679.800 65.600 2680.660 65.980 ;
  RECT 1368.250 192.510 1368.500 195.930 ;
  RECT 1368.820 192.790 1369.070 193.650 ;
  RECT 1409.170 192.510 1409.420 195.930 ;
  RECT 1409.740 192.790 1409.990 193.650 ;
  RECT 1450.090 192.510 1450.340 195.930 ;
  RECT 1450.660 192.790 1450.910 193.650 ;
  RECT 1491.010 192.510 1491.260 195.930 ;
  RECT 1491.580 192.790 1491.830 193.650 ;
  RECT 1531.930 192.510 1532.180 195.930 ;
  RECT 1532.500 192.790 1532.750 193.650 ;
  RECT 1572.850 192.510 1573.100 195.930 ;
  RECT 1573.420 192.790 1573.670 193.650 ;
  RECT 1613.770 192.510 1614.020 195.930 ;
  RECT 1614.340 192.790 1614.590 193.650 ;
  RECT 1654.690 192.510 1654.940 195.930 ;
  RECT 1655.260 192.790 1655.510 193.650 ;
  RECT 1695.610 192.510 1695.860 195.930 ;
  RECT 1696.180 192.790 1696.430 193.650 ;
  RECT 1736.530 192.510 1736.780 195.930 ;
  RECT 1737.100 192.790 1737.350 193.650 ;
  RECT 1777.450 192.510 1777.700 195.930 ;
  RECT 1778.020 192.790 1778.270 193.650 ;
  RECT 1818.370 192.510 1818.620 195.930 ;
  RECT 1818.940 192.790 1819.190 193.650 ;
  RECT 1859.290 192.510 1859.540 195.930 ;
  RECT 1859.860 192.790 1860.110 193.650 ;
  RECT 1900.210 192.510 1900.460 195.930 ;
  RECT 1900.780 192.790 1901.030 193.650 ;
  RECT 1941.130 192.510 1941.380 195.930 ;
  RECT 1941.700 192.790 1941.950 193.650 ;
  RECT 1982.050 192.510 1982.300 195.930 ;
  RECT 1982.620 192.790 1982.870 193.650 ;
  RECT 2022.970 192.510 2023.220 195.930 ;
  RECT 2023.540 192.790 2023.790 193.650 ;
  RECT 2063.890 192.510 2064.140 195.930 ;
  RECT 2064.460 192.790 2064.710 193.650 ;
  RECT 2104.810 192.510 2105.060 195.930 ;
  RECT 2105.380 192.790 2105.630 193.650 ;
  RECT 2145.730 192.510 2145.980 195.930 ;
  RECT 2146.300 192.790 2146.550 193.650 ;
  RECT 2186.650 192.510 2186.900 195.930 ;
  RECT 2187.220 192.790 2187.470 193.650 ;
  RECT 2227.570 192.510 2227.820 195.930 ;
  RECT 2228.140 192.790 2228.390 193.650 ;
  RECT 2268.490 192.510 2268.740 195.930 ;
  RECT 2269.060 192.790 2269.310 193.650 ;
  RECT 2309.410 192.510 2309.660 195.930 ;
  RECT 2309.980 192.790 2310.230 193.650 ;
  RECT 2350.330 192.510 2350.580 195.930 ;
  RECT 2350.900 192.790 2351.150 193.650 ;
  RECT 2391.250 192.510 2391.500 195.930 ;
  RECT 2391.820 192.790 2392.070 193.650 ;
  RECT 2432.170 192.510 2432.420 195.930 ;
  RECT 2432.740 192.790 2432.990 193.650 ;
  RECT 2473.090 192.510 2473.340 195.930 ;
  RECT 2473.660 192.790 2473.910 193.650 ;
  RECT 2514.010 192.510 2514.260 195.930 ;
  RECT 2514.580 192.790 2514.830 193.650 ;
  RECT 2554.930 192.510 2555.180 195.930 ;
  RECT 2555.500 192.790 2555.750 193.650 ;
  RECT 2595.850 192.510 2596.100 195.930 ;
  RECT 2596.420 192.790 2596.670 193.650 ;
  RECT 2636.770 192.510 2637.020 195.930 ;
  RECT 2637.340 192.790 2637.590 193.650 ;
  RECT 1364.760 192.510 1365.660 195.930 ;
  RECT 1335.440 192.510 1338.630 195.930 ;
  RECT 1345.440 192.510 1349.760 195.930 ;
  RECT 1351.810 192.790 1354.320 193.650 ;
  RECT 1339.390 192.790 1341.780 193.650 ;
  RECT 1331.880 192.790 1334.940 193.650 ;
  RECT 1356.060 192.790 1358.910 193.650 ;
  RECT 1360.360 192.790 1363.610 193.650 ;
  RECT 1327.160 192.510 1328.920 195.930 ;
  RECT 1329.160 192.790 1330.920 193.650 ;
  RECT 1317.900 192.510 1319.580 195.930 ;
  RECT 1321.820 192.510 1323.580 195.930 ;
  RECT 1319.820 192.790 1321.580 193.650 ;
  RECT 1323.820 192.790 1325.580 193.650 ;
  RECT 1316.800 192.510 1317.700 195.930 ;
  RECT 4.280 65.600 5.140 65.980 ;
  RECT 2.000 68.240 5.420 69.440 ;
  RECT 2.000 70.720 5.420 71.920 ;
  RECT 4.280 69.940 5.140 70.220 ;
  RECT 2.000 71.920 5.420 73.120 ;
  RECT 2.000 74.400 5.420 75.600 ;
  RECT 4.280 73.620 5.140 73.900 ;
  RECT 2.000 75.600 5.420 76.800 ;
  RECT 2.000 78.080 5.420 79.280 ;
  RECT 4.280 77.300 5.140 77.580 ;
  RECT 2.000 79.280 5.420 80.480 ;
  RECT 2.000 81.760 5.420 82.960 ;
  RECT 4.280 80.980 5.140 81.260 ;
  RECT 2.000 82.960 5.420 84.160 ;
  RECT 2.000 85.440 5.420 86.640 ;
  RECT 4.280 84.660 5.140 84.940 ;
  RECT 2.000 86.640 5.420 87.840 ;
  RECT 2.000 89.120 5.420 90.320 ;
  RECT 4.280 88.340 5.140 88.620 ;
  RECT 2.000 90.320 5.420 91.520 ;
  RECT 2.000 92.800 5.420 94.000 ;
  RECT 4.280 92.020 5.140 92.300 ;
  RECT 2.000 94.000 5.420 95.200 ;
  RECT 2.000 96.480 5.420 97.680 ;
  RECT 4.280 95.700 5.140 95.980 ;
  RECT 2.000 97.680 5.420 98.880 ;
  RECT 2.000 100.160 5.420 101.360 ;
  RECT 4.280 99.380 5.140 99.660 ;
  RECT 2.000 101.360 5.420 102.560 ;
  RECT 2.000 103.840 5.420 105.040 ;
  RECT 4.280 103.060 5.140 103.340 ;
  RECT 2.000 105.040 5.420 106.240 ;
  RECT 2.000 107.520 5.420 108.720 ;
  RECT 4.280 106.740 5.140 107.020 ;
  RECT 2.000 108.720 5.420 109.920 ;
  RECT 2.000 111.200 5.420 112.400 ;
  RECT 4.280 110.420 5.140 110.700 ;
  RECT 2.000 112.400 5.420 113.600 ;
  RECT 2.000 114.880 5.420 116.080 ;
  RECT 4.280 114.100 5.140 114.380 ;
  RECT 2.000 116.080 5.420 117.280 ;
  RECT 2.000 118.560 5.420 119.760 ;
  RECT 4.280 117.780 5.140 118.060 ;
  RECT 2.000 119.760 5.420 120.960 ;
  RECT 2.000 122.240 5.420 123.440 ;
  RECT 4.280 121.460 5.140 121.740 ;
  RECT 2.000 123.440 5.420 124.640 ;
  RECT 2.000 125.920 5.420 127.120 ;
  RECT 4.280 125.140 5.140 125.420 ;
  RECT 2.000 127.120 5.420 128.320 ;
  RECT 2.000 129.600 5.420 130.800 ;
  RECT 4.280 128.820 5.140 129.100 ;
  RECT 2.000 130.800 5.420 132.000 ;
  RECT 2.000 133.280 5.420 134.480 ;
  RECT 4.280 132.500 5.140 132.780 ;
  RECT 2.000 134.480 5.420 135.680 ;
  RECT 2.000 136.960 5.420 138.160 ;
  RECT 4.280 136.180 5.140 136.460 ;
  RECT 2.000 138.160 5.420 139.360 ;
  RECT 2.000 140.640 5.420 141.840 ;
  RECT 4.280 139.860 5.140 140.140 ;
  RECT 2.000 141.840 5.420 143.040 ;
  RECT 2.000 144.320 5.420 145.520 ;
  RECT 4.280 143.540 5.140 143.820 ;
  RECT 2.000 145.520 5.420 146.720 ;
  RECT 2.000 148.000 5.420 149.200 ;
  RECT 4.280 147.220 5.140 147.500 ;
  RECT 2.000 149.200 5.420 150.400 ;
  RECT 2.000 151.680 5.420 152.880 ;
  RECT 4.280 150.900 5.140 151.180 ;
  RECT 2.000 152.880 5.420 154.080 ;
  RECT 2.000 155.360 5.420 156.560 ;
  RECT 4.280 154.580 5.140 154.860 ;
  RECT 2.000 156.560 5.420 157.760 ;
  RECT 2.000 159.040 5.420 160.240 ;
  RECT 4.280 158.260 5.140 158.540 ;
  RECT 2.000 160.240 5.420 161.440 ;
  RECT 2.000 162.720 5.420 163.920 ;
  RECT 4.280 161.940 5.140 162.220 ;
  RECT 2.000 163.920 5.420 165.120 ;
  RECT 2.000 166.400 5.420 167.600 ;
  RECT 4.280 165.620 5.140 165.900 ;
  RECT 2.000 167.600 5.420 168.800 ;
  RECT 2.000 170.080 5.420 171.280 ;
  RECT 4.280 169.300 5.140 169.580 ;
  RECT 2.000 171.280 5.420 172.480 ;
  RECT 2.000 173.760 5.420 174.960 ;
  RECT 4.280 172.980 5.140 173.260 ;
  RECT 2.000 174.960 5.420 176.160 ;
  RECT 2.000 177.440 5.420 178.640 ;
  RECT 4.280 176.660 5.140 176.940 ;
  RECT 2.000 178.640 5.420 179.840 ;
  RECT 2.000 181.120 5.420 182.320 ;
  RECT 4.280 180.340 5.140 180.620 ;
  RECT 2.000 182.320 5.420 183.520 ;
  RECT 2.000 184.800 5.420 186.000 ;
  RECT 4.280 184.020 5.140 184.300 ;
  RECT 4.280 191.940 5.140 192.320 ;
  RECT 47.920 192.510 48.170 195.930 ;
  RECT 47.350 192.790 47.600 193.650 ;
  RECT 88.840 192.510 89.090 195.930 ;
  RECT 88.270 192.790 88.520 193.650 ;
  RECT 129.760 192.510 130.010 195.930 ;
  RECT 129.190 192.790 129.440 193.650 ;
  RECT 170.680 192.510 170.930 195.930 ;
  RECT 170.110 192.790 170.360 193.650 ;
  RECT 211.600 192.510 211.850 195.930 ;
  RECT 211.030 192.790 211.280 193.650 ;
  RECT 252.520 192.510 252.770 195.930 ;
  RECT 251.950 192.790 252.200 193.650 ;
  RECT 293.440 192.510 293.690 195.930 ;
  RECT 292.870 192.790 293.120 193.650 ;
  RECT 334.360 192.510 334.610 195.930 ;
  RECT 333.790 192.790 334.040 193.650 ;
  RECT 375.280 192.510 375.530 195.930 ;
  RECT 374.710 192.790 374.960 193.650 ;
  RECT 416.200 192.510 416.450 195.930 ;
  RECT 415.630 192.790 415.880 193.650 ;
  RECT 457.120 192.510 457.370 195.930 ;
  RECT 456.550 192.790 456.800 193.650 ;
  RECT 498.040 192.510 498.290 195.930 ;
  RECT 497.470 192.790 497.720 193.650 ;
  RECT 538.960 192.510 539.210 195.930 ;
  RECT 538.390 192.790 538.640 193.650 ;
  RECT 579.880 192.510 580.130 195.930 ;
  RECT 579.310 192.790 579.560 193.650 ;
  RECT 620.800 192.510 621.050 195.930 ;
  RECT 620.230 192.790 620.480 193.650 ;
  RECT 661.720 192.510 661.970 195.930 ;
  RECT 661.150 192.790 661.400 193.650 ;
  RECT 702.640 192.510 702.890 195.930 ;
  RECT 702.070 192.790 702.320 193.650 ;
  RECT 743.560 192.510 743.810 195.930 ;
  RECT 742.990 192.790 743.240 193.650 ;
  RECT 784.480 192.510 784.730 195.930 ;
  RECT 783.910 192.790 784.160 193.650 ;
  RECT 825.400 192.510 825.650 195.930 ;
  RECT 824.830 192.790 825.080 193.650 ;
  RECT 866.320 192.510 866.570 195.930 ;
  RECT 865.750 192.790 866.000 193.650 ;
  RECT 907.240 192.510 907.490 195.930 ;
  RECT 906.670 192.790 906.920 193.650 ;
  RECT 948.160 192.510 948.410 195.930 ;
  RECT 947.590 192.790 947.840 193.650 ;
  RECT 989.080 192.510 989.330 195.930 ;
  RECT 988.510 192.790 988.760 193.650 ;
  RECT 1030.000 192.510 1030.250 195.930 ;
  RECT 1029.430 192.790 1029.680 193.650 ;
  RECT 1070.920 192.510 1071.170 195.930 ;
  RECT 1070.350 192.790 1070.600 193.650 ;
  RECT 1111.840 192.510 1112.090 195.930 ;
  RECT 1111.270 192.790 1111.520 193.650 ;
  RECT 1152.760 192.510 1153.010 195.930 ;
  RECT 1152.190 192.790 1152.440 193.650 ;
  RECT 1193.680 192.510 1193.930 195.930 ;
  RECT 1193.110 192.790 1193.360 193.650 ;
  RECT 1234.600 192.510 1234.850 195.930 ;
  RECT 1234.030 192.790 1234.280 193.650 ;
  RECT 1275.520 192.510 1275.770 195.930 ;
  RECT 1274.950 192.790 1275.200 193.650 ;
  RECT 0.000 195.930 2684.940 197.930 ;
  RECT 0.000 1.600 2684.940 3.600 ;
  RECT 2682.940 1.600 2684.940 197.930 ;
  RECT 0.000 1.600 2.000 197.930 ;
  LAYER ME2 ;
  RECT 5.420 7.020 2679.520 192.510 ;
  RECT 2683.080 3.460 2684.940 196.070 ;
  RECT 0.000 3.460 1.860 196.070 ;
  RECT 1.860 196.070 2683.080 197.930 ;
  RECT 2674.600 1.600 2683.080 3.460 ;
  RECT 2660.200 1.600 2672.280 3.460 ;
  RECT 2655.000 1.600 2657.650 3.460 ;
  RECT 2640.200 1.600 2652.440 3.460 ;
  RECT 2633.800 1.600 2637.810 3.460 ;
  RECT 2619.400 1.600 2631.360 3.460 ;
  RECT 2614.200 1.600 2616.730 3.460 ;
  RECT 2599.400 1.600 2611.520 3.460 ;
  RECT 2593.000 1.600 2596.890 3.460 ;
  RECT 2578.200 1.600 2590.440 3.460 ;
  RECT 2573.000 1.600 2575.810 3.460 ;
  RECT 2558.600 1.600 2570.600 3.460 ;
  RECT 2552.200 1.600 2555.970 3.460 ;
  RECT 2537.400 1.600 2549.520 3.460 ;
  RECT 2532.200 1.600 2534.890 3.460 ;
  RECT 2517.400 1.600 2529.680 3.460 ;
  RECT 2511.000 1.600 2515.050 3.460 ;
  RECT 2496.600 1.600 2508.600 3.460 ;
  RECT 2491.400 1.600 2493.970 3.460 ;
  RECT 2476.600 1.600 2488.760 3.460 ;
  RECT 2470.200 1.600 2474.130 3.460 ;
  RECT 2455.400 1.600 2467.680 3.460 ;
  RECT 2450.200 1.600 2453.050 3.460 ;
  RECT 2435.800 1.600 2447.840 3.460 ;
  RECT 2429.400 1.600 2433.210 3.460 ;
  RECT 2414.600 1.600 2426.760 3.460 ;
  RECT 2409.400 1.600 2412.130 3.460 ;
  RECT 2394.600 1.600 2406.920 3.460 ;
  RECT 2388.200 1.600 2392.290 3.460 ;
  RECT 2373.800 1.600 2385.840 3.460 ;
  RECT 2368.600 1.600 2371.210 3.460 ;
  RECT 2355.400 1.600 2366.000 3.460 ;
  RECT 2347.400 1.600 2351.370 3.460 ;
  RECT 2332.600 1.600 2344.920 3.460 ;
  RECT 2327.400 1.600 2330.290 3.460 ;
  RECT 2313.000 1.600 2325.080 3.460 ;
  RECT 2306.600 1.600 2310.450 3.460 ;
  RECT 2291.800 1.600 2304.000 3.460 ;
  RECT 2286.600 1.600 2289.370 3.460 ;
  RECT 2272.200 1.600 2284.160 3.460 ;
  RECT 2265.400 1.600 2269.530 3.460 ;
  RECT 2251.000 1.600 2263.080 3.460 ;
  RECT 2245.800 1.600 2248.450 3.460 ;
  RECT 2231.000 1.600 2243.240 3.460 ;
  RECT 2224.600 1.600 2228.610 3.460 ;
  RECT 2210.200 1.600 2222.160 3.460 ;
  RECT 2205.000 1.600 2207.530 3.460 ;
  RECT 2190.200 1.600 2202.320 3.460 ;
  RECT 2183.800 1.600 2187.690 3.460 ;
  RECT 2169.000 1.600 2181.240 3.460 ;
  RECT 2163.800 1.600 2166.610 3.460 ;
  RECT 2149.400 1.600 2161.400 3.460 ;
  RECT 2143.000 1.600 2146.770 3.460 ;
  RECT 2128.200 1.600 2140.320 3.460 ;
  RECT 2123.000 1.600 2125.690 3.460 ;
  RECT 2108.200 1.600 2120.480 3.460 ;
  RECT 2101.800 1.600 2105.850 3.460 ;
  RECT 2087.400 1.600 2099.400 3.460 ;
  RECT 2082.200 1.600 2084.770 3.460 ;
  RECT 2067.400 1.600 2079.560 3.460 ;
  RECT 2061.000 1.600 2064.930 3.460 ;
  RECT 2046.200 1.600 2058.480 3.460 ;
  RECT 2041.000 1.600 2043.850 3.460 ;
  RECT 2028.200 1.600 2038.640 3.460 ;
  RECT 2020.200 1.600 2024.010 3.460 ;
  RECT 2005.400 1.600 2017.560 3.460 ;
  RECT 2000.200 1.600 2002.930 3.460 ;
  RECT 1985.400 1.600 1997.720 3.460 ;
  RECT 1979.000 1.600 1983.090 3.460 ;
  RECT 1964.600 1.600 1976.640 3.460 ;
  RECT 1959.400 1.600 1962.010 3.460 ;
  RECT 1944.600 1.600 1956.800 3.460 ;
  RECT 1938.200 1.600 1942.170 3.460 ;
  RECT 1923.400 1.600 1935.720 3.460 ;
  RECT 1918.200 1.600 1921.090 3.460 ;
  RECT 1903.800 1.600 1915.880 3.460 ;
  RECT 1897.400 1.600 1901.250 3.460 ;
  RECT 1882.600 1.600 1894.800 3.460 ;
  RECT 1877.400 1.600 1880.170 3.460 ;
  RECT 1863.000 1.600 1874.960 3.460 ;
  RECT 1856.200 1.600 1860.330 3.460 ;
  RECT 1841.800 1.600 1853.880 3.460 ;
  RECT 1836.600 1.600 1839.250 3.460 ;
  RECT 1821.800 1.600 1834.040 3.460 ;
  RECT 1815.400 1.600 1819.410 3.460 ;
  RECT 1801.000 1.600 1812.960 3.460 ;
  RECT 1795.800 1.600 1798.330 3.460 ;
  RECT 1781.000 1.600 1793.120 3.460 ;
  RECT 1774.600 1.600 1778.490 3.460 ;
  RECT 1759.800 1.600 1772.040 3.460 ;
  RECT 1754.600 1.600 1757.410 3.460 ;
  RECT 1740.200 1.600 1752.200 3.460 ;
  RECT 1733.800 1.600 1737.570 3.460 ;
  RECT 1719.000 1.600 1731.120 3.460 ;
  RECT 1713.800 1.600 1716.490 3.460 ;
  RECT 1701.000 1.600 1711.280 3.460 ;
  RECT 1692.600 1.600 1696.650 3.460 ;
  RECT 1678.200 1.600 1690.200 3.460 ;
  RECT 1673.000 1.600 1675.570 3.460 ;
  RECT 1658.200 1.600 1670.360 3.460 ;
  RECT 1651.800 1.600 1655.730 3.460 ;
  RECT 1637.000 1.600 1649.280 3.460 ;
  RECT 1631.800 1.600 1634.650 3.460 ;
  RECT 1617.400 1.600 1629.440 3.460 ;
  RECT 1611.000 1.600 1614.810 3.460 ;
  RECT 1596.200 1.600 1608.360 3.460 ;
  RECT 1591.000 1.600 1593.730 3.460 ;
  RECT 1576.200 1.600 1588.520 3.460 ;
  RECT 1569.800 1.600 1573.890 3.460 ;
  RECT 1555.400 1.600 1567.440 3.460 ;
  RECT 1550.200 1.600 1552.810 3.460 ;
  RECT 1535.400 1.600 1547.600 3.460 ;
  RECT 1529.000 1.600 1532.970 3.460 ;
  RECT 1514.200 1.600 1526.520 3.460 ;
  RECT 1509.000 1.600 1511.890 3.460 ;
  RECT 1494.600 1.600 1506.680 3.460 ;
  RECT 1488.200 1.600 1492.050 3.460 ;
  RECT 1473.400 1.600 1485.600 3.460 ;
  RECT 1468.200 1.600 1470.970 3.460 ;
  RECT 1453.800 1.600 1465.760 3.460 ;
  RECT 1447.000 1.600 1451.130 3.460 ;
  RECT 1432.600 1.600 1444.680 3.460 ;
  RECT 1427.400 1.600 1430.050 3.460 ;
  RECT 1412.600 1.600 1424.840 3.460 ;
  RECT 1406.200 1.600 1410.210 3.460 ;
  RECT 1391.800 1.600 1403.760 3.460 ;
  RECT 1386.600 1.600 1389.130 3.460 ;
  RECT 1373.400 1.600 1383.920 3.460 ;
  RECT 1351.000 1.600 1369.290 3.460 ;
  RECT 1339.000 1.600 1342.450 3.460 ;
  RECT 1331.800 1.600 1336.480 3.460 ;
  RECT 1313.000 1.600 1317.360 3.460 ;
  RECT 1298.200 1.600 1310.460 3.460 ;
  RECT 1293.000 1.600 1295.830 3.460 ;
  RECT 1278.600 1.600 1290.620 3.460 ;
  RECT 1272.200 1.600 1275.990 3.460 ;
  RECT 1257.400 1.600 1269.540 3.460 ;
  RECT 1252.200 1.600 1254.910 3.460 ;
  RECT 1237.400 1.600 1249.700 3.460 ;
  RECT 1231.000 1.600 1235.070 3.460 ;
  RECT 1216.600 1.600 1228.620 3.460 ;
  RECT 1211.400 1.600 1213.990 3.460 ;
  RECT 1196.600 1.600 1208.780 3.460 ;
  RECT 1190.200 1.600 1194.150 3.460 ;
  RECT 1175.400 1.600 1187.700 3.460 ;
  RECT 1170.200 1.600 1173.070 3.460 ;
  RECT 1155.800 1.600 1167.860 3.460 ;
  RECT 1149.400 1.600 1153.230 3.460 ;
  RECT 1134.600 1.600 1146.780 3.460 ;
  RECT 1129.400 1.600 1132.150 3.460 ;
  RECT 1115.000 1.600 1126.940 3.460 ;
  RECT 1108.200 1.600 1112.310 3.460 ;
  RECT 1093.800 1.600 1105.860 3.460 ;
  RECT 1088.600 1.600 1091.230 3.460 ;
  RECT 1073.800 1.600 1086.020 3.460 ;
  RECT 1067.400 1.600 1071.390 3.460 ;
  RECT 1053.000 1.600 1064.940 3.460 ;
  RECT 1047.400 1.600 1050.310 3.460 ;
  RECT 1033.000 1.600 1045.100 3.460 ;
  RECT 1026.600 1.600 1030.470 3.460 ;
  RECT 1011.800 1.600 1024.020 3.460 ;
  RECT 1006.600 1.600 1009.390 3.460 ;
  RECT 993.800 1.600 1004.180 3.460 ;
  RECT 985.400 1.600 989.550 3.460 ;
  RECT 971.000 1.600 983.100 3.460 ;
  RECT 965.800 1.600 968.470 3.460 ;
  RECT 951.000 1.600 963.260 3.460 ;
  RECT 944.600 1.600 948.630 3.460 ;
  RECT 930.200 1.600 942.180 3.460 ;
  RECT 925.000 1.600 927.550 3.460 ;
  RECT 910.200 1.600 922.340 3.460 ;
  RECT 903.800 1.600 907.710 3.460 ;
  RECT 889.000 1.600 901.260 3.460 ;
  RECT 883.800 1.600 886.630 3.460 ;
  RECT 869.400 1.600 881.420 3.460 ;
  RECT 863.000 1.600 866.790 3.460 ;
  RECT 848.200 1.600 860.340 3.460 ;
  RECT 843.000 1.600 845.710 3.460 ;
  RECT 828.200 1.600 840.500 3.460 ;
  RECT 821.800 1.600 825.870 3.460 ;
  RECT 807.400 1.600 819.420 3.460 ;
  RECT 802.200 1.600 804.790 3.460 ;
  RECT 787.400 1.600 799.580 3.460 ;
  RECT 781.000 1.600 784.950 3.460 ;
  RECT 766.200 1.600 778.500 3.460 ;
  RECT 761.000 1.600 763.870 3.460 ;
  RECT 746.600 1.600 758.660 3.460 ;
  RECT 740.200 1.600 744.030 3.460 ;
  RECT 725.400 1.600 737.580 3.460 ;
  RECT 720.200 1.600 722.950 3.460 ;
  RECT 705.800 1.600 717.740 3.460 ;
  RECT 699.000 1.600 703.110 3.460 ;
  RECT 684.600 1.600 696.660 3.460 ;
  RECT 679.400 1.600 682.030 3.460 ;
  RECT 666.600 1.600 676.820 3.460 ;
  RECT 658.200 1.600 662.190 3.460 ;
  RECT 643.800 1.600 655.740 3.460 ;
  RECT 638.200 1.600 641.110 3.460 ;
  RECT 623.800 1.600 635.900 3.460 ;
  RECT 617.400 1.600 621.270 3.460 ;
  RECT 602.600 1.600 614.820 3.460 ;
  RECT 597.400 1.600 600.190 3.460 ;
  RECT 583.000 1.600 594.980 3.460 ;
  RECT 576.200 1.600 580.350 3.460 ;
  RECT 561.800 1.600 573.900 3.460 ;
  RECT 556.600 1.600 559.270 3.460 ;
  RECT 541.800 1.600 554.060 3.460 ;
  RECT 535.400 1.600 539.430 3.460 ;
  RECT 521.000 1.600 532.980 3.460 ;
  RECT 515.800 1.600 518.350 3.460 ;
  RECT 501.000 1.600 513.140 3.460 ;
  RECT 494.600 1.600 498.510 3.460 ;
  RECT 479.800 1.600 492.060 3.460 ;
  RECT 474.600 1.600 477.430 3.460 ;
  RECT 460.200 1.600 472.220 3.460 ;
  RECT 453.800 1.600 457.590 3.460 ;
  RECT 439.000 1.600 451.140 3.460 ;
  RECT 433.800 1.600 436.510 3.460 ;
  RECT 419.000 1.600 431.300 3.460 ;
  RECT 412.600 1.600 416.670 3.460 ;
  RECT 398.200 1.600 410.220 3.460 ;
  RECT 393.000 1.600 395.590 3.460 ;
  RECT 378.200 1.600 390.380 3.460 ;
  RECT 371.800 1.600 375.750 3.460 ;
  RECT 357.000 1.600 369.300 3.460 ;
  RECT 351.800 1.600 354.670 3.460 ;
  RECT 339.000 1.600 349.460 3.460 ;
  RECT 331.000 1.600 334.830 3.460 ;
  RECT 316.200 1.600 328.380 3.460 ;
  RECT 311.000 1.600 313.750 3.460 ;
  RECT 296.600 1.600 308.540 3.460 ;
  RECT 289.800 1.600 293.910 3.460 ;
  RECT 275.400 1.600 287.460 3.460 ;
  RECT 270.200 1.600 272.830 3.460 ;
  RECT 255.400 1.600 267.620 3.460 ;
  RECT 249.000 1.600 252.990 3.460 ;
  RECT 234.600 1.600 246.540 3.460 ;
  RECT 229.000 1.600 231.910 3.460 ;
  RECT 214.600 1.600 226.700 3.460 ;
  RECT 208.200 1.600 212.070 3.460 ;
  RECT 193.400 1.600 205.620 3.460 ;
  RECT 188.200 1.600 190.990 3.460 ;
  RECT 173.800 1.600 185.780 3.460 ;
  RECT 167.000 1.600 171.150 3.460 ;
  RECT 152.600 1.600 164.700 3.460 ;
  RECT 147.400 1.600 150.070 3.460 ;
  RECT 132.600 1.600 144.860 3.460 ;
  RECT 126.200 1.600 130.230 3.460 ;
  RECT 111.800 1.600 123.780 3.460 ;
  RECT 106.600 1.600 109.150 3.460 ;
  RECT 91.800 1.600 103.940 3.460 ;
  RECT 85.400 1.600 89.310 3.460 ;
  RECT 70.600 1.600 82.860 3.460 ;
  RECT 65.400 1.600 68.230 3.460 ;
  RECT 51.000 1.600 63.020 3.460 ;
  RECT 44.600 1.600 48.390 3.460 ;
  RECT 29.800 1.600 41.940 3.460 ;
  RECT 24.600 1.600 27.310 3.460 ;
  RECT 11.800 1.600 22.100 3.460 ;
  RECT 1.860 1.600 7.470 3.460 ;
  RECT 2680.940 5.600 2682.800 193.930 ;
  RECT 2.140 5.600 4.000 193.930 ;
  RECT 4.000 193.930 2680.940 195.790 ;
  RECT 2674.600 3.740 2680.940 5.600 ;
  RECT 2660.200 3.740 2672.280 5.600 ;
  RECT 2655.000 3.740 2657.650 5.600 ;
  RECT 2640.200 3.740 2652.440 5.600 ;
  RECT 2633.800 3.740 2637.810 5.600 ;
  RECT 2619.400 3.740 2631.360 5.600 ;
  RECT 2614.200 3.740 2616.730 5.600 ;
  RECT 2599.400 3.740 2611.520 5.600 ;
  RECT 2593.000 3.740 2596.890 5.600 ;
  RECT 2578.200 3.740 2590.440 5.600 ;
  RECT 2573.000 3.740 2575.810 5.600 ;
  RECT 2558.600 3.740 2570.600 5.600 ;
  RECT 2552.200 3.740 2555.970 5.600 ;
  RECT 2537.400 3.740 2549.520 5.600 ;
  RECT 2532.200 3.740 2534.890 5.600 ;
  RECT 2517.400 3.740 2529.680 5.600 ;
  RECT 2511.000 3.740 2515.050 5.600 ;
  RECT 2496.600 3.740 2508.600 5.600 ;
  RECT 2491.400 3.740 2493.970 5.600 ;
  RECT 2476.600 3.740 2488.760 5.600 ;
  RECT 2470.200 3.740 2474.130 5.600 ;
  RECT 2455.400 3.740 2467.680 5.600 ;
  RECT 2450.200 3.740 2453.050 5.600 ;
  RECT 2435.800 3.740 2447.840 5.600 ;
  RECT 2429.400 3.740 2433.210 5.600 ;
  RECT 2414.600 3.740 2426.760 5.600 ;
  RECT 2409.400 3.740 2412.130 5.600 ;
  RECT 2394.600 3.740 2406.920 5.600 ;
  RECT 2388.200 3.740 2392.290 5.600 ;
  RECT 2373.800 3.740 2385.840 5.600 ;
  RECT 2368.600 3.740 2371.210 5.600 ;
  RECT 2355.400 3.740 2366.000 5.600 ;
  RECT 2347.400 3.740 2351.370 5.600 ;
  RECT 2332.600 3.740 2344.920 5.600 ;
  RECT 2327.400 3.740 2330.290 5.600 ;
  RECT 2313.000 3.740 2325.080 5.600 ;
  RECT 2306.600 3.740 2310.450 5.600 ;
  RECT 2291.800 3.740 2304.000 5.600 ;
  RECT 2286.600 3.740 2289.370 5.600 ;
  RECT 2272.200 3.740 2284.160 5.600 ;
  RECT 2265.400 3.740 2269.530 5.600 ;
  RECT 2251.000 3.740 2263.080 5.600 ;
  RECT 2245.800 3.740 2248.450 5.600 ;
  RECT 2231.000 3.740 2243.240 5.600 ;
  RECT 2224.600 3.740 2228.610 5.600 ;
  RECT 2210.200 3.740 2222.160 5.600 ;
  RECT 2205.000 3.740 2207.530 5.600 ;
  RECT 2190.200 3.740 2202.320 5.600 ;
  RECT 2183.800 3.740 2187.690 5.600 ;
  RECT 2169.000 3.740 2181.240 5.600 ;
  RECT 2163.800 3.740 2166.610 5.600 ;
  RECT 2149.400 3.740 2161.400 5.600 ;
  RECT 2143.000 3.740 2146.770 5.600 ;
  RECT 2128.200 3.740 2140.320 5.600 ;
  RECT 2123.000 3.740 2125.690 5.600 ;
  RECT 2108.200 3.740 2120.480 5.600 ;
  RECT 2101.800 3.740 2105.850 5.600 ;
  RECT 2087.400 3.740 2099.400 5.600 ;
  RECT 2082.200 3.740 2084.770 5.600 ;
  RECT 2067.400 3.740 2079.560 5.600 ;
  RECT 2061.000 3.740 2064.930 5.600 ;
  RECT 2046.200 3.740 2058.480 5.600 ;
  RECT 2041.000 3.740 2043.850 5.600 ;
  RECT 2028.200 3.740 2038.640 5.600 ;
  RECT 2020.200 3.740 2024.010 5.600 ;
  RECT 2005.400 3.740 2017.560 5.600 ;
  RECT 2000.200 3.740 2002.930 5.600 ;
  RECT 1985.400 3.740 1997.720 5.600 ;
  RECT 1979.000 3.740 1983.090 5.600 ;
  RECT 1964.600 3.740 1976.640 5.600 ;
  RECT 1959.400 3.740 1962.010 5.600 ;
  RECT 1944.600 3.740 1956.800 5.600 ;
  RECT 1938.200 3.740 1942.170 5.600 ;
  RECT 1923.400 3.740 1935.720 5.600 ;
  RECT 1918.200 3.740 1921.090 5.600 ;
  RECT 1903.800 3.740 1915.880 5.600 ;
  RECT 1897.400 3.740 1901.250 5.600 ;
  RECT 1882.600 3.740 1894.800 5.600 ;
  RECT 1877.400 3.740 1880.170 5.600 ;
  RECT 1863.000 3.740 1874.960 5.600 ;
  RECT 1856.200 3.740 1860.330 5.600 ;
  RECT 1841.800 3.740 1853.880 5.600 ;
  RECT 1836.600 3.740 1839.250 5.600 ;
  RECT 1821.800 3.740 1834.040 5.600 ;
  RECT 1815.400 3.740 1819.410 5.600 ;
  RECT 1801.000 3.740 1812.960 5.600 ;
  RECT 1795.800 3.740 1798.330 5.600 ;
  RECT 1781.000 3.740 1793.120 5.600 ;
  RECT 1774.600 3.740 1778.490 5.600 ;
  RECT 1759.800 3.740 1772.040 5.600 ;
  RECT 1754.600 3.740 1757.410 5.600 ;
  RECT 1740.200 3.740 1752.200 5.600 ;
  RECT 1733.800 3.740 1737.570 5.600 ;
  RECT 1719.000 3.740 1731.120 5.600 ;
  RECT 1713.800 3.740 1716.490 5.600 ;
  RECT 1701.000 3.740 1711.280 5.600 ;
  RECT 1692.600 3.740 1696.650 5.600 ;
  RECT 1678.200 3.740 1690.200 5.600 ;
  RECT 1673.000 3.740 1675.570 5.600 ;
  RECT 1658.200 3.740 1670.360 5.600 ;
  RECT 1651.800 3.740 1655.730 5.600 ;
  RECT 1637.000 3.740 1649.280 5.600 ;
  RECT 1631.800 3.740 1634.650 5.600 ;
  RECT 1617.400 3.740 1629.440 5.600 ;
  RECT 1611.000 3.740 1614.810 5.600 ;
  RECT 1596.200 3.740 1608.360 5.600 ;
  RECT 1591.000 3.740 1593.730 5.600 ;
  RECT 1576.200 3.740 1588.520 5.600 ;
  RECT 1569.800 3.740 1573.890 5.600 ;
  RECT 1555.400 3.740 1567.440 5.600 ;
  RECT 1550.200 3.740 1552.810 5.600 ;
  RECT 1535.400 3.740 1547.600 5.600 ;
  RECT 1529.000 3.740 1532.970 5.600 ;
  RECT 1514.200 3.740 1526.520 5.600 ;
  RECT 1509.000 3.740 1511.890 5.600 ;
  RECT 1494.600 3.740 1506.680 5.600 ;
  RECT 1488.200 3.740 1492.050 5.600 ;
  RECT 1473.400 3.740 1485.600 5.600 ;
  RECT 1468.200 3.740 1470.970 5.600 ;
  RECT 1453.800 3.740 1465.760 5.600 ;
  RECT 1447.000 3.740 1451.130 5.600 ;
  RECT 1432.600 3.740 1444.680 5.600 ;
  RECT 1427.400 3.740 1430.050 5.600 ;
  RECT 1412.600 3.740 1424.840 5.600 ;
  RECT 1406.200 3.740 1410.210 5.600 ;
  RECT 1391.800 3.740 1403.760 5.600 ;
  RECT 1386.600 3.740 1389.130 5.600 ;
  RECT 1373.400 3.740 1383.920 5.600 ;
  RECT 1351.000 3.740 1369.290 5.600 ;
  RECT 1339.000 3.740 1342.450 5.600 ;
  RECT 1331.800 3.740 1336.480 5.600 ;
  RECT 1313.000 3.740 1317.360 5.600 ;
  RECT 1298.200 3.740 1310.460 5.600 ;
  RECT 1293.000 3.740 1295.830 5.600 ;
  RECT 1278.600 3.740 1290.620 5.600 ;
  RECT 1272.200 3.740 1275.990 5.600 ;
  RECT 1257.400 3.740 1269.540 5.600 ;
  RECT 1252.200 3.740 1254.910 5.600 ;
  RECT 1237.400 3.740 1249.700 5.600 ;
  RECT 1231.000 3.740 1235.070 5.600 ;
  RECT 1216.600 3.740 1228.620 5.600 ;
  RECT 1211.400 3.740 1213.990 5.600 ;
  RECT 1196.600 3.740 1208.780 5.600 ;
  RECT 1190.200 3.740 1194.150 5.600 ;
  RECT 1175.400 3.740 1187.700 5.600 ;
  RECT 1170.200 3.740 1173.070 5.600 ;
  RECT 1155.800 3.740 1167.860 5.600 ;
  RECT 1149.400 3.740 1153.230 5.600 ;
  RECT 1134.600 3.740 1146.780 5.600 ;
  RECT 1129.400 3.740 1132.150 5.600 ;
  RECT 1115.000 3.740 1126.940 5.600 ;
  RECT 1108.200 3.740 1112.310 5.600 ;
  RECT 1093.800 3.740 1105.860 5.600 ;
  RECT 1088.600 3.740 1091.230 5.600 ;
  RECT 1073.800 3.740 1086.020 5.600 ;
  RECT 1067.400 3.740 1071.390 5.600 ;
  RECT 1053.000 3.740 1064.940 5.600 ;
  RECT 1047.400 3.740 1050.310 5.600 ;
  RECT 1033.000 3.740 1045.100 5.600 ;
  RECT 1026.600 3.740 1030.470 5.600 ;
  RECT 1011.800 3.740 1024.020 5.600 ;
  RECT 1006.600 3.740 1009.390 5.600 ;
  RECT 993.800 3.740 1004.180 5.600 ;
  RECT 985.400 3.740 989.550 5.600 ;
  RECT 971.000 3.740 983.100 5.600 ;
  RECT 965.800 3.740 968.470 5.600 ;
  RECT 951.000 3.740 963.260 5.600 ;
  RECT 944.600 3.740 948.630 5.600 ;
  RECT 930.200 3.740 942.180 5.600 ;
  RECT 925.000 3.740 927.550 5.600 ;
  RECT 910.200 3.740 922.340 5.600 ;
  RECT 903.800 3.740 907.710 5.600 ;
  RECT 889.000 3.740 901.260 5.600 ;
  RECT 883.800 3.740 886.630 5.600 ;
  RECT 869.400 3.740 881.420 5.600 ;
  RECT 863.000 3.740 866.790 5.600 ;
  RECT 848.200 3.740 860.340 5.600 ;
  RECT 843.000 3.740 845.710 5.600 ;
  RECT 828.200 3.740 840.500 5.600 ;
  RECT 821.800 3.740 825.870 5.600 ;
  RECT 807.400 3.740 819.420 5.600 ;
  RECT 802.200 3.740 804.790 5.600 ;
  RECT 787.400 3.740 799.580 5.600 ;
  RECT 781.000 3.740 784.950 5.600 ;
  RECT 766.200 3.740 778.500 5.600 ;
  RECT 761.000 3.740 763.870 5.600 ;
  RECT 746.600 3.740 758.660 5.600 ;
  RECT 740.200 3.740 744.030 5.600 ;
  RECT 725.400 3.740 737.580 5.600 ;
  RECT 720.200 3.740 722.950 5.600 ;
  RECT 705.800 3.740 717.740 5.600 ;
  RECT 699.000 3.740 703.110 5.600 ;
  RECT 684.600 3.740 696.660 5.600 ;
  RECT 679.400 3.740 682.030 5.600 ;
  RECT 666.600 3.740 676.820 5.600 ;
  RECT 658.200 3.740 662.190 5.600 ;
  RECT 643.800 3.740 655.740 5.600 ;
  RECT 638.200 3.740 641.110 5.600 ;
  RECT 623.800 3.740 635.900 5.600 ;
  RECT 617.400 3.740 621.270 5.600 ;
  RECT 602.600 3.740 614.820 5.600 ;
  RECT 597.400 3.740 600.190 5.600 ;
  RECT 583.000 3.740 594.980 5.600 ;
  RECT 576.200 3.740 580.350 5.600 ;
  RECT 561.800 3.740 573.900 5.600 ;
  RECT 556.600 3.740 559.270 5.600 ;
  RECT 541.800 3.740 554.060 5.600 ;
  RECT 535.400 3.740 539.430 5.600 ;
  RECT 521.000 3.740 532.980 5.600 ;
  RECT 515.800 3.740 518.350 5.600 ;
  RECT 501.000 3.740 513.140 5.600 ;
  RECT 494.600 3.740 498.510 5.600 ;
  RECT 479.800 3.740 492.060 5.600 ;
  RECT 474.600 3.740 477.430 5.600 ;
  RECT 460.200 3.740 472.220 5.600 ;
  RECT 453.800 3.740 457.590 5.600 ;
  RECT 439.000 3.740 451.140 5.600 ;
  RECT 433.800 3.740 436.510 5.600 ;
  RECT 419.000 3.740 431.300 5.600 ;
  RECT 412.600 3.740 416.670 5.600 ;
  RECT 398.200 3.740 410.220 5.600 ;
  RECT 393.000 3.740 395.590 5.600 ;
  RECT 378.200 3.740 390.380 5.600 ;
  RECT 371.800 3.740 375.750 5.600 ;
  RECT 357.000 3.740 369.300 5.600 ;
  RECT 351.800 3.740 354.670 5.600 ;
  RECT 339.000 3.740 349.460 5.600 ;
  RECT 331.000 3.740 334.830 5.600 ;
  RECT 316.200 3.740 328.380 5.600 ;
  RECT 311.000 3.740 313.750 5.600 ;
  RECT 296.600 3.740 308.540 5.600 ;
  RECT 289.800 3.740 293.910 5.600 ;
  RECT 275.400 3.740 287.460 5.600 ;
  RECT 270.200 3.740 272.830 5.600 ;
  RECT 255.400 3.740 267.620 5.600 ;
  RECT 249.000 3.740 252.990 5.600 ;
  RECT 234.600 3.740 246.540 5.600 ;
  RECT 229.000 3.740 231.910 5.600 ;
  RECT 214.600 3.740 226.700 5.600 ;
  RECT 208.200 3.740 212.070 5.600 ;
  RECT 193.400 3.740 205.620 5.600 ;
  RECT 188.200 3.740 190.990 5.600 ;
  RECT 173.800 3.740 185.780 5.600 ;
  RECT 167.000 3.740 171.150 5.600 ;
  RECT 152.600 3.740 164.700 5.600 ;
  RECT 147.400 3.740 150.070 5.600 ;
  RECT 132.600 3.740 144.860 5.600 ;
  RECT 126.200 3.740 130.230 5.600 ;
  RECT 111.800 3.740 123.780 5.600 ;
  RECT 106.600 3.740 109.150 5.600 ;
  RECT 91.800 3.740 103.940 5.600 ;
  RECT 85.400 3.740 89.310 5.600 ;
  RECT 70.600 3.740 82.860 5.600 ;
  RECT 65.400 3.740 68.230 5.600 ;
  RECT 51.000 3.740 63.020 5.600 ;
  RECT 44.600 3.740 48.390 5.600 ;
  RECT 29.800 3.740 41.940 5.600 ;
  RECT 24.600 3.740 27.310 5.600 ;
  RECT 11.800 3.740 22.100 5.600 ;
  RECT 4.000 3.740 7.470 5.600 ;
  RECT 2.140 193.930 4.000 195.790 ;
  RECT 0.000 196.070 1.860 197.930 ;
  RECT 2680.940 3.740 2682.800 5.600 ;
  RECT 2683.080 1.600 2684.940 3.460 ;
  RECT 2680.940 193.930 2682.800 195.790 ;
  RECT 2683.080 196.070 2684.940 197.930 ;
  RECT 2.140 3.740 4.000 5.600 ;
  RECT 0.000 1.600 1.860 3.460 ;
  RECT 2672.800 0.000 2673.600 1.000 ;
  RECT 2673.100 1.000 2673.300 5.200 ;
  RECT 2673.100 5.200 2673.480 5.400 ;
  RECT 2673.280 5.400 2673.480 7.020 ;
  RECT 2658.400 0.000 2659.200 1.000 ;
  RECT 2658.700 1.000 2658.900 5.200 ;
  RECT 2658.650 5.200 2658.900 5.400 ;
  RECT 2658.650 5.400 2658.850 7.020 ;
  RECT 2653.200 0.000 2654.000 1.000 ;
  RECT 2653.500 1.000 2653.700 5.200 ;
  RECT 2653.440 5.200 2653.700 5.400 ;
  RECT 2653.440 5.400 2653.640 7.020 ;
  RECT 2638.400 0.000 2639.200 1.000 ;
  RECT 2638.700 1.000 2638.900 5.200 ;
  RECT 2638.700 5.200 2639.010 5.400 ;
  RECT 2638.810 5.400 2639.010 7.020 ;
  RECT 2632.000 0.000 2632.800 1.000 ;
  RECT 2632.300 1.000 2632.500 5.200 ;
  RECT 2632.300 5.200 2632.560 5.400 ;
  RECT 2632.360 5.400 2632.560 7.020 ;
  RECT 2617.600 0.000 2618.400 1.000 ;
  RECT 2617.900 1.000 2618.100 5.200 ;
  RECT 2617.730 5.200 2618.100 5.400 ;
  RECT 2617.730 5.400 2617.930 7.020 ;
  RECT 2612.400 0.000 2613.200 1.000 ;
  RECT 2612.700 1.000 2612.900 5.200 ;
  RECT 2612.520 5.200 2612.900 5.400 ;
  RECT 2612.520 5.400 2612.720 7.020 ;
  RECT 2597.600 0.000 2598.400 1.000 ;
  RECT 2597.900 1.000 2598.100 5.200 ;
  RECT 2597.890 5.200 2598.100 5.400 ;
  RECT 2597.890 5.400 2598.090 7.020 ;
  RECT 2591.200 0.000 2592.000 1.000 ;
  RECT 2591.500 1.000 2591.700 5.200 ;
  RECT 2591.440 5.200 2591.700 5.400 ;
  RECT 2591.440 5.400 2591.640 7.020 ;
  RECT 2576.400 0.000 2577.200 1.000 ;
  RECT 2576.700 1.000 2576.900 5.200 ;
  RECT 2576.700 5.200 2577.010 5.400 ;
  RECT 2576.810 5.400 2577.010 7.020 ;
  RECT 2571.200 0.000 2572.000 1.000 ;
  RECT 2571.500 1.000 2571.700 5.200 ;
  RECT 2571.500 5.200 2571.800 5.400 ;
  RECT 2571.600 5.400 2571.800 7.020 ;
  RECT 2556.800 0.000 2557.600 1.000 ;
  RECT 2557.100 1.000 2557.300 5.200 ;
  RECT 2556.970 5.200 2557.300 5.400 ;
  RECT 2556.970 5.400 2557.170 7.020 ;
  RECT 2550.400 0.000 2551.200 1.000 ;
  RECT 2550.700 1.000 2550.900 5.200 ;
  RECT 2550.520 5.200 2550.900 5.400 ;
  RECT 2550.520 5.400 2550.720 7.020 ;
  RECT 2535.600 0.000 2536.400 1.000 ;
  RECT 2535.900 1.000 2536.100 5.200 ;
  RECT 2535.890 5.200 2536.100 5.400 ;
  RECT 2535.890 5.400 2536.090 7.020 ;
  RECT 2530.400 0.000 2531.200 1.000 ;
  RECT 2530.700 1.000 2530.900 5.200 ;
  RECT 2530.680 5.200 2530.900 5.400 ;
  RECT 2530.680 5.400 2530.880 7.020 ;
  RECT 2515.600 0.000 2516.400 1.000 ;
  RECT 2515.900 1.000 2516.100 5.200 ;
  RECT 2515.900 5.200 2516.250 5.400 ;
  RECT 2516.050 5.400 2516.250 7.020 ;
  RECT 2509.200 0.000 2510.000 1.000 ;
  RECT 2509.500 1.000 2509.700 5.200 ;
  RECT 2509.500 5.200 2509.800 5.400 ;
  RECT 2509.600 5.400 2509.800 7.020 ;
  RECT 2494.800 0.000 2495.600 1.000 ;
  RECT 2495.100 1.000 2495.300 5.200 ;
  RECT 2494.970 5.200 2495.300 5.400 ;
  RECT 2494.970 5.400 2495.170 7.020 ;
  RECT 2489.600 0.000 2490.400 1.000 ;
  RECT 2489.900 1.000 2490.100 5.200 ;
  RECT 2489.760 5.200 2490.100 5.400 ;
  RECT 2489.760 5.400 2489.960 7.020 ;
  RECT 2474.800 0.000 2475.600 1.000 ;
  RECT 2475.100 1.000 2475.300 5.200 ;
  RECT 2475.100 5.200 2475.330 5.400 ;
  RECT 2475.130 5.400 2475.330 7.020 ;
  RECT 2468.400 0.000 2469.200 1.000 ;
  RECT 2468.700 1.000 2468.900 5.200 ;
  RECT 2468.680 5.200 2468.900 5.400 ;
  RECT 2468.680 5.400 2468.880 7.020 ;
  RECT 2453.600 0.000 2454.400 1.000 ;
  RECT 2453.900 1.000 2454.100 5.200 ;
  RECT 2453.900 5.200 2454.250 5.400 ;
  RECT 2454.050 5.400 2454.250 7.020 ;
  RECT 2448.400 0.000 2449.200 1.000 ;
  RECT 2448.700 1.000 2448.900 5.200 ;
  RECT 2448.700 5.200 2449.040 5.400 ;
  RECT 2448.840 5.400 2449.040 7.020 ;
  RECT 2434.000 0.000 2434.800 1.000 ;
  RECT 2434.300 1.000 2434.500 5.200 ;
  RECT 2434.210 5.200 2434.500 5.400 ;
  RECT 2434.210 5.400 2434.410 7.020 ;
  RECT 2427.600 0.000 2428.400 1.000 ;
  RECT 2427.900 1.000 2428.100 5.200 ;
  RECT 2427.760 5.200 2428.100 5.400 ;
  RECT 2427.760 5.400 2427.960 7.020 ;
  RECT 2412.800 0.000 2413.600 1.000 ;
  RECT 2413.100 1.000 2413.300 5.200 ;
  RECT 2413.100 5.200 2413.330 5.400 ;
  RECT 2413.130 5.400 2413.330 7.020 ;
  RECT 2407.600 0.000 2408.400 1.000 ;
  RECT 2407.900 1.000 2408.100 5.200 ;
  RECT 2407.900 5.200 2408.120 5.400 ;
  RECT 2407.920 5.400 2408.120 7.020 ;
  RECT 2392.800 0.000 2393.600 1.000 ;
  RECT 2393.100 1.000 2393.300 5.200 ;
  RECT 2393.100 5.200 2393.490 5.400 ;
  RECT 2393.290 5.400 2393.490 7.020 ;
  RECT 2386.400 0.000 2387.200 1.000 ;
  RECT 2386.700 1.000 2386.900 5.200 ;
  RECT 2386.700 5.200 2387.040 5.400 ;
  RECT 2386.840 5.400 2387.040 7.020 ;
  RECT 2372.000 0.000 2372.800 1.000 ;
  RECT 2372.300 1.000 2372.500 5.200 ;
  RECT 2372.210 5.200 2372.500 5.400 ;
  RECT 2372.210 5.400 2372.410 7.020 ;
  RECT 2366.800 0.000 2367.600 1.000 ;
  RECT 2367.100 1.000 2367.300 5.200 ;
  RECT 2367.000 5.200 2367.300 5.400 ;
  RECT 2367.000 5.400 2367.200 7.020 ;
  RECT 2353.600 0.000 2354.400 1.000 ;
  RECT 2353.900 1.000 2354.100 5.200 ;
  RECT 2353.900 5.200 2354.290 5.400 ;
  RECT 2354.090 5.400 2354.290 7.020 ;
  RECT 2352.000 0.000 2352.800 1.000 ;
  RECT 2352.300 1.000 2352.500 5.200 ;
  RECT 2352.300 5.200 2352.570 5.400 ;
  RECT 2352.370 5.400 2352.570 7.020 ;
  RECT 2345.600 0.000 2346.400 1.000 ;
  RECT 2345.900 1.000 2346.100 5.200 ;
  RECT 2345.900 5.200 2346.120 5.400 ;
  RECT 2345.920 5.400 2346.120 7.020 ;
  RECT 2330.800 0.000 2331.600 1.000 ;
  RECT 2331.100 1.000 2331.300 5.200 ;
  RECT 2331.100 5.200 2331.490 5.400 ;
  RECT 2331.290 5.400 2331.490 7.020 ;
  RECT 2325.600 0.000 2326.400 1.000 ;
  RECT 2325.900 1.000 2326.100 5.200 ;
  RECT 2325.900 5.200 2326.280 5.400 ;
  RECT 2326.080 5.400 2326.280 7.020 ;
  RECT 2311.200 0.000 2312.000 1.000 ;
  RECT 2311.500 1.000 2311.700 5.200 ;
  RECT 2311.450 5.200 2311.700 5.400 ;
  RECT 2311.450 5.400 2311.650 7.020 ;
  RECT 2304.800 0.000 2305.600 1.000 ;
  RECT 2305.100 1.000 2305.300 5.200 ;
  RECT 2305.000 5.200 2305.300 5.400 ;
  RECT 2305.000 5.400 2305.200 7.020 ;
  RECT 2290.000 0.000 2290.800 1.000 ;
  RECT 2290.300 1.000 2290.500 5.200 ;
  RECT 2290.300 5.200 2290.570 5.400 ;
  RECT 2290.370 5.400 2290.570 7.020 ;
  RECT 2284.800 0.000 2285.600 1.000 ;
  RECT 2285.100 1.000 2285.300 5.200 ;
  RECT 2285.100 5.200 2285.360 5.400 ;
  RECT 2285.160 5.400 2285.360 7.020 ;
  RECT 2270.400 0.000 2271.200 1.000 ;
  RECT 2270.700 1.000 2270.900 5.200 ;
  RECT 2270.530 5.200 2270.900 5.400 ;
  RECT 2270.530 5.400 2270.730 7.020 ;
  RECT 2263.600 0.000 2264.400 1.000 ;
  RECT 2263.900 1.000 2264.100 5.200 ;
  RECT 2263.900 5.200 2264.280 5.400 ;
  RECT 2264.080 5.400 2264.280 7.020 ;
  RECT 2249.200 0.000 2250.000 1.000 ;
  RECT 2249.500 1.000 2249.700 5.200 ;
  RECT 2249.450 5.200 2249.700 5.400 ;
  RECT 2249.450 5.400 2249.650 7.020 ;
  RECT 2244.000 0.000 2244.800 1.000 ;
  RECT 2244.300 1.000 2244.500 5.200 ;
  RECT 2244.240 5.200 2244.500 5.400 ;
  RECT 2244.240 5.400 2244.440 7.020 ;
  RECT 2229.200 0.000 2230.000 1.000 ;
  RECT 2229.500 1.000 2229.700 5.200 ;
  RECT 2229.500 5.200 2229.810 5.400 ;
  RECT 2229.610 5.400 2229.810 7.020 ;
  RECT 2222.800 0.000 2223.600 1.000 ;
  RECT 2223.100 1.000 2223.300 5.200 ;
  RECT 2223.100 5.200 2223.360 5.400 ;
  RECT 2223.160 5.400 2223.360 7.020 ;
  RECT 2208.400 0.000 2209.200 1.000 ;
  RECT 2208.700 1.000 2208.900 5.200 ;
  RECT 2208.530 5.200 2208.900 5.400 ;
  RECT 2208.530 5.400 2208.730 7.020 ;
  RECT 2203.200 0.000 2204.000 1.000 ;
  RECT 2203.500 1.000 2203.700 5.200 ;
  RECT 2203.320 5.200 2203.700 5.400 ;
  RECT 2203.320 5.400 2203.520 7.020 ;
  RECT 2188.400 0.000 2189.200 1.000 ;
  RECT 2188.700 1.000 2188.900 5.200 ;
  RECT 2188.690 5.200 2188.900 5.400 ;
  RECT 2188.690 5.400 2188.890 7.020 ;
  RECT 2182.000 0.000 2182.800 1.000 ;
  RECT 2182.300 1.000 2182.500 5.200 ;
  RECT 2182.240 5.200 2182.500 5.400 ;
  RECT 2182.240 5.400 2182.440 7.020 ;
  RECT 2167.200 0.000 2168.000 1.000 ;
  RECT 2167.500 1.000 2167.700 5.200 ;
  RECT 2167.500 5.200 2167.810 5.400 ;
  RECT 2167.610 5.400 2167.810 7.020 ;
  RECT 2162.000 0.000 2162.800 1.000 ;
  RECT 2162.300 1.000 2162.500 5.200 ;
  RECT 2162.300 5.200 2162.600 5.400 ;
  RECT 2162.400 5.400 2162.600 7.020 ;
  RECT 2147.600 0.000 2148.400 1.000 ;
  RECT 2147.900 1.000 2148.100 5.200 ;
  RECT 2147.770 5.200 2148.100 5.400 ;
  RECT 2147.770 5.400 2147.970 7.020 ;
  RECT 2141.200 0.000 2142.000 1.000 ;
  RECT 2141.500 1.000 2141.700 5.200 ;
  RECT 2141.320 5.200 2141.700 5.400 ;
  RECT 2141.320 5.400 2141.520 7.020 ;
  RECT 2126.400 0.000 2127.200 1.000 ;
  RECT 2126.700 1.000 2126.900 5.200 ;
  RECT 2126.690 5.200 2126.900 5.400 ;
  RECT 2126.690 5.400 2126.890 7.020 ;
  RECT 2121.200 0.000 2122.000 1.000 ;
  RECT 2121.500 1.000 2121.700 5.200 ;
  RECT 2121.480 5.200 2121.700 5.400 ;
  RECT 2121.480 5.400 2121.680 7.020 ;
  RECT 2106.400 0.000 2107.200 1.000 ;
  RECT 2106.700 1.000 2106.900 5.200 ;
  RECT 2106.700 5.200 2107.050 5.400 ;
  RECT 2106.850 5.400 2107.050 7.020 ;
  RECT 2100.000 0.000 2100.800 1.000 ;
  RECT 2100.300 1.000 2100.500 5.200 ;
  RECT 2100.300 5.200 2100.600 5.400 ;
  RECT 2100.400 5.400 2100.600 7.020 ;
  RECT 2085.600 0.000 2086.400 1.000 ;
  RECT 2085.900 1.000 2086.100 5.200 ;
  RECT 2085.770 5.200 2086.100 5.400 ;
  RECT 2085.770 5.400 2085.970 7.020 ;
  RECT 2080.400 0.000 2081.200 1.000 ;
  RECT 2080.700 1.000 2080.900 5.200 ;
  RECT 2080.560 5.200 2080.900 5.400 ;
  RECT 2080.560 5.400 2080.760 7.020 ;
  RECT 2065.600 0.000 2066.400 1.000 ;
  RECT 2065.900 1.000 2066.100 5.200 ;
  RECT 2065.900 5.200 2066.130 5.400 ;
  RECT 2065.930 5.400 2066.130 7.020 ;
  RECT 2059.200 0.000 2060.000 1.000 ;
  RECT 2059.500 1.000 2059.700 5.200 ;
  RECT 2059.480 5.200 2059.700 5.400 ;
  RECT 2059.480 5.400 2059.680 7.020 ;
  RECT 2044.400 0.000 2045.200 1.000 ;
  RECT 2044.700 1.000 2044.900 5.200 ;
  RECT 2044.700 5.200 2045.050 5.400 ;
  RECT 2044.850 5.400 2045.050 7.020 ;
  RECT 2039.200 0.000 2040.000 1.000 ;
  RECT 2039.500 1.000 2039.700 5.200 ;
  RECT 2039.500 5.200 2039.840 5.400 ;
  RECT 2039.640 5.400 2039.840 7.020 ;
  RECT 2026.400 0.000 2027.200 1.000 ;
  RECT 2026.700 1.000 2026.900 5.200 ;
  RECT 2026.700 5.200 2026.930 5.400 ;
  RECT 2026.730 5.400 2026.930 7.020 ;
  RECT 2024.800 0.000 2025.600 1.000 ;
  RECT 2025.100 1.000 2025.300 5.200 ;
  RECT 2025.010 5.200 2025.300 5.400 ;
  RECT 2025.010 5.400 2025.210 7.020 ;
  RECT 2018.400 0.000 2019.200 1.000 ;
  RECT 2018.700 1.000 2018.900 5.200 ;
  RECT 2018.560 5.200 2018.900 5.400 ;
  RECT 2018.560 5.400 2018.760 7.020 ;
  RECT 2003.600 0.000 2004.400 1.000 ;
  RECT 2003.900 1.000 2004.100 5.200 ;
  RECT 2003.900 5.200 2004.130 5.400 ;
  RECT 2003.930 5.400 2004.130 7.020 ;
  RECT 1998.400 0.000 1999.200 1.000 ;
  RECT 1998.700 1.000 1998.900 5.200 ;
  RECT 1998.700 5.200 1998.920 5.400 ;
  RECT 1998.720 5.400 1998.920 7.020 ;
  RECT 1983.600 0.000 1984.400 1.000 ;
  RECT 1983.900 1.000 1984.100 5.200 ;
  RECT 1983.900 5.200 1984.290 5.400 ;
  RECT 1984.090 5.400 1984.290 7.020 ;
  RECT 1977.200 0.000 1978.000 1.000 ;
  RECT 1977.500 1.000 1977.700 5.200 ;
  RECT 1977.500 5.200 1977.840 5.400 ;
  RECT 1977.640 5.400 1977.840 7.020 ;
  RECT 1962.800 0.000 1963.600 1.000 ;
  RECT 1963.100 1.000 1963.300 5.200 ;
  RECT 1963.010 5.200 1963.300 5.400 ;
  RECT 1963.010 5.400 1963.210 7.020 ;
  RECT 1957.600 0.000 1958.400 1.000 ;
  RECT 1957.900 1.000 1958.100 5.200 ;
  RECT 1957.800 5.200 1958.100 5.400 ;
  RECT 1957.800 5.400 1958.000 7.020 ;
  RECT 1942.800 0.000 1943.600 1.000 ;
  RECT 1943.100 1.000 1943.300 5.200 ;
  RECT 1943.100 5.200 1943.370 5.400 ;
  RECT 1943.170 5.400 1943.370 7.020 ;
  RECT 1936.400 0.000 1937.200 1.000 ;
  RECT 1936.700 1.000 1936.900 5.200 ;
  RECT 1936.700 5.200 1936.920 5.400 ;
  RECT 1936.720 5.400 1936.920 7.020 ;
  RECT 1921.600 0.000 1922.400 1.000 ;
  RECT 1921.900 1.000 1922.100 5.200 ;
  RECT 1921.900 5.200 1922.290 5.400 ;
  RECT 1922.090 5.400 1922.290 7.020 ;
  RECT 1916.400 0.000 1917.200 1.000 ;
  RECT 1916.700 1.000 1916.900 5.200 ;
  RECT 1916.700 5.200 1917.080 5.400 ;
  RECT 1916.880 5.400 1917.080 7.020 ;
  RECT 1902.000 0.000 1902.800 1.000 ;
  RECT 1902.300 1.000 1902.500 5.200 ;
  RECT 1902.250 5.200 1902.500 5.400 ;
  RECT 1902.250 5.400 1902.450 7.020 ;
  RECT 1895.600 0.000 1896.400 1.000 ;
  RECT 1895.900 1.000 1896.100 5.200 ;
  RECT 1895.800 5.200 1896.100 5.400 ;
  RECT 1895.800 5.400 1896.000 7.020 ;
  RECT 1880.800 0.000 1881.600 1.000 ;
  RECT 1881.100 1.000 1881.300 5.200 ;
  RECT 1881.100 5.200 1881.370 5.400 ;
  RECT 1881.170 5.400 1881.370 7.020 ;
  RECT 1875.600 0.000 1876.400 1.000 ;
  RECT 1875.900 1.000 1876.100 5.200 ;
  RECT 1875.900 5.200 1876.160 5.400 ;
  RECT 1875.960 5.400 1876.160 7.020 ;
  RECT 1861.200 0.000 1862.000 1.000 ;
  RECT 1861.500 1.000 1861.700 5.200 ;
  RECT 1861.330 5.200 1861.700 5.400 ;
  RECT 1861.330 5.400 1861.530 7.020 ;
  RECT 1854.400 0.000 1855.200 1.000 ;
  RECT 1854.700 1.000 1854.900 5.200 ;
  RECT 1854.700 5.200 1855.080 5.400 ;
  RECT 1854.880 5.400 1855.080 7.020 ;
  RECT 1840.000 0.000 1840.800 1.000 ;
  RECT 1840.300 1.000 1840.500 5.200 ;
  RECT 1840.250 5.200 1840.500 5.400 ;
  RECT 1840.250 5.400 1840.450 7.020 ;
  RECT 1834.800 0.000 1835.600 1.000 ;
  RECT 1835.100 1.000 1835.300 5.200 ;
  RECT 1835.040 5.200 1835.300 5.400 ;
  RECT 1835.040 5.400 1835.240 7.020 ;
  RECT 1820.000 0.000 1820.800 1.000 ;
  RECT 1820.300 1.000 1820.500 5.200 ;
  RECT 1820.300 5.200 1820.610 5.400 ;
  RECT 1820.410 5.400 1820.610 7.020 ;
  RECT 1813.600 0.000 1814.400 1.000 ;
  RECT 1813.900 1.000 1814.100 5.200 ;
  RECT 1813.900 5.200 1814.160 5.400 ;
  RECT 1813.960 5.400 1814.160 7.020 ;
  RECT 1799.200 0.000 1800.000 1.000 ;
  RECT 1799.500 1.000 1799.700 5.200 ;
  RECT 1799.330 5.200 1799.700 5.400 ;
  RECT 1799.330 5.400 1799.530 7.020 ;
  RECT 1794.000 0.000 1794.800 1.000 ;
  RECT 1794.300 1.000 1794.500 5.200 ;
  RECT 1794.120 5.200 1794.500 5.400 ;
  RECT 1794.120 5.400 1794.320 7.020 ;
  RECT 1779.200 0.000 1780.000 1.000 ;
  RECT 1779.500 1.000 1779.700 5.200 ;
  RECT 1779.490 5.200 1779.700 5.400 ;
  RECT 1779.490 5.400 1779.690 7.020 ;
  RECT 1772.800 0.000 1773.600 1.000 ;
  RECT 1773.100 1.000 1773.300 5.200 ;
  RECT 1773.040 5.200 1773.300 5.400 ;
  RECT 1773.040 5.400 1773.240 7.020 ;
  RECT 1758.000 0.000 1758.800 1.000 ;
  RECT 1758.300 1.000 1758.500 5.200 ;
  RECT 1758.300 5.200 1758.610 5.400 ;
  RECT 1758.410 5.400 1758.610 7.020 ;
  RECT 1752.800 0.000 1753.600 1.000 ;
  RECT 1753.100 1.000 1753.300 5.200 ;
  RECT 1753.100 5.200 1753.400 5.400 ;
  RECT 1753.200 5.400 1753.400 7.020 ;
  RECT 1738.400 0.000 1739.200 1.000 ;
  RECT 1738.700 1.000 1738.900 5.200 ;
  RECT 1738.570 5.200 1738.900 5.400 ;
  RECT 1738.570 5.400 1738.770 7.020 ;
  RECT 1732.000 0.000 1732.800 1.000 ;
  RECT 1732.300 1.000 1732.500 5.200 ;
  RECT 1732.120 5.200 1732.500 5.400 ;
  RECT 1732.120 5.400 1732.320 7.020 ;
  RECT 1717.200 0.000 1718.000 1.000 ;
  RECT 1717.500 1.000 1717.700 5.200 ;
  RECT 1717.490 5.200 1717.700 5.400 ;
  RECT 1717.490 5.400 1717.690 7.020 ;
  RECT 1712.000 0.000 1712.800 1.000 ;
  RECT 1712.300 1.000 1712.500 5.200 ;
  RECT 1712.280 5.200 1712.500 5.400 ;
  RECT 1712.280 5.400 1712.480 7.020 ;
  RECT 1699.200 0.000 1700.000 1.000 ;
  RECT 1699.500 1.000 1699.700 5.200 ;
  RECT 1699.370 5.200 1699.700 5.400 ;
  RECT 1699.370 5.400 1699.570 7.020 ;
  RECT 1697.200 0.000 1698.000 1.000 ;
  RECT 1697.500 1.000 1697.700 5.200 ;
  RECT 1697.500 5.200 1697.850 5.400 ;
  RECT 1697.650 5.400 1697.850 7.020 ;
  RECT 1690.800 0.000 1691.600 1.000 ;
  RECT 1691.100 1.000 1691.300 5.200 ;
  RECT 1691.100 5.200 1691.400 5.400 ;
  RECT 1691.200 5.400 1691.400 7.020 ;
  RECT 1676.400 0.000 1677.200 1.000 ;
  RECT 1676.700 1.000 1676.900 5.200 ;
  RECT 1676.570 5.200 1676.900 5.400 ;
  RECT 1676.570 5.400 1676.770 7.020 ;
  RECT 1671.200 0.000 1672.000 1.000 ;
  RECT 1671.500 1.000 1671.700 5.200 ;
  RECT 1671.360 5.200 1671.700 5.400 ;
  RECT 1671.360 5.400 1671.560 7.020 ;
  RECT 1656.400 0.000 1657.200 1.000 ;
  RECT 1656.700 1.000 1656.900 5.200 ;
  RECT 1656.700 5.200 1656.930 5.400 ;
  RECT 1656.730 5.400 1656.930 7.020 ;
  RECT 1650.000 0.000 1650.800 1.000 ;
  RECT 1650.300 1.000 1650.500 5.200 ;
  RECT 1650.280 5.200 1650.500 5.400 ;
  RECT 1650.280 5.400 1650.480 7.020 ;
  RECT 1635.200 0.000 1636.000 1.000 ;
  RECT 1635.500 1.000 1635.700 5.200 ;
  RECT 1635.500 5.200 1635.850 5.400 ;
  RECT 1635.650 5.400 1635.850 7.020 ;
  RECT 1630.000 0.000 1630.800 1.000 ;
  RECT 1630.300 1.000 1630.500 5.200 ;
  RECT 1630.300 5.200 1630.640 5.400 ;
  RECT 1630.440 5.400 1630.640 7.020 ;
  RECT 1615.600 0.000 1616.400 1.000 ;
  RECT 1615.900 1.000 1616.100 5.200 ;
  RECT 1615.810 5.200 1616.100 5.400 ;
  RECT 1615.810 5.400 1616.010 7.020 ;
  RECT 1609.200 0.000 1610.000 1.000 ;
  RECT 1609.500 1.000 1609.700 5.200 ;
  RECT 1609.360 5.200 1609.700 5.400 ;
  RECT 1609.360 5.400 1609.560 7.020 ;
  RECT 1594.400 0.000 1595.200 1.000 ;
  RECT 1594.700 1.000 1594.900 5.200 ;
  RECT 1594.700 5.200 1594.930 5.400 ;
  RECT 1594.730 5.400 1594.930 7.020 ;
  RECT 1589.200 0.000 1590.000 1.000 ;
  RECT 1589.500 1.000 1589.700 5.200 ;
  RECT 1589.500 5.200 1589.720 5.400 ;
  RECT 1589.520 5.400 1589.720 7.020 ;
  RECT 1574.400 0.000 1575.200 1.000 ;
  RECT 1574.700 1.000 1574.900 5.200 ;
  RECT 1574.700 5.200 1575.090 5.400 ;
  RECT 1574.890 5.400 1575.090 7.020 ;
  RECT 1568.000 0.000 1568.800 1.000 ;
  RECT 1568.300 1.000 1568.500 5.200 ;
  RECT 1568.300 5.200 1568.640 5.400 ;
  RECT 1568.440 5.400 1568.640 7.020 ;
  RECT 1553.600 0.000 1554.400 1.000 ;
  RECT 1553.900 1.000 1554.100 5.200 ;
  RECT 1553.810 5.200 1554.100 5.400 ;
  RECT 1553.810 5.400 1554.010 7.020 ;
  RECT 1548.400 0.000 1549.200 1.000 ;
  RECT 1548.700 1.000 1548.900 5.200 ;
  RECT 1548.600 5.200 1548.900 5.400 ;
  RECT 1548.600 5.400 1548.800 7.020 ;
  RECT 1533.600 0.000 1534.400 1.000 ;
  RECT 1533.900 1.000 1534.100 5.200 ;
  RECT 1533.900 5.200 1534.170 5.400 ;
  RECT 1533.970 5.400 1534.170 7.020 ;
  RECT 1527.200 0.000 1528.000 1.000 ;
  RECT 1527.500 1.000 1527.700 5.200 ;
  RECT 1527.500 5.200 1527.720 5.400 ;
  RECT 1527.520 5.400 1527.720 7.020 ;
  RECT 1512.400 0.000 1513.200 1.000 ;
  RECT 1512.700 1.000 1512.900 5.200 ;
  RECT 1512.700 5.200 1513.090 5.400 ;
  RECT 1512.890 5.400 1513.090 7.020 ;
  RECT 1507.200 0.000 1508.000 1.000 ;
  RECT 1507.500 1.000 1507.700 5.200 ;
  RECT 1507.500 5.200 1507.880 5.400 ;
  RECT 1507.680 5.400 1507.880 7.020 ;
  RECT 1492.800 0.000 1493.600 1.000 ;
  RECT 1493.100 1.000 1493.300 5.200 ;
  RECT 1493.050 5.200 1493.300 5.400 ;
  RECT 1493.050 5.400 1493.250 7.020 ;
  RECT 1486.400 0.000 1487.200 1.000 ;
  RECT 1486.700 1.000 1486.900 5.200 ;
  RECT 1486.600 5.200 1486.900 5.400 ;
  RECT 1486.600 5.400 1486.800 7.020 ;
  RECT 1471.600 0.000 1472.400 1.000 ;
  RECT 1471.900 1.000 1472.100 5.200 ;
  RECT 1471.900 5.200 1472.170 5.400 ;
  RECT 1471.970 5.400 1472.170 7.020 ;
  RECT 1466.400 0.000 1467.200 1.000 ;
  RECT 1466.700 1.000 1466.900 5.200 ;
  RECT 1466.700 5.200 1466.960 5.400 ;
  RECT 1466.760 5.400 1466.960 7.020 ;
  RECT 1452.000 0.000 1452.800 1.000 ;
  RECT 1452.300 1.000 1452.500 5.200 ;
  RECT 1452.130 5.200 1452.500 5.400 ;
  RECT 1452.130 5.400 1452.330 7.020 ;
  RECT 1445.200 0.000 1446.000 1.000 ;
  RECT 1445.500 1.000 1445.700 5.200 ;
  RECT 1445.500 5.200 1445.880 5.400 ;
  RECT 1445.680 5.400 1445.880 7.020 ;
  RECT 1430.800 0.000 1431.600 1.000 ;
  RECT 1431.100 1.000 1431.300 5.200 ;
  RECT 1431.050 5.200 1431.300 5.400 ;
  RECT 1431.050 5.400 1431.250 7.020 ;
  RECT 1425.600 0.000 1426.400 1.000 ;
  RECT 1425.900 1.000 1426.100 5.200 ;
  RECT 1425.840 5.200 1426.100 5.400 ;
  RECT 1425.840 5.400 1426.040 7.020 ;
  RECT 1410.800 0.000 1411.600 1.000 ;
  RECT 1411.100 1.000 1411.300 5.200 ;
  RECT 1411.100 5.200 1411.410 5.400 ;
  RECT 1411.210 5.400 1411.410 7.020 ;
  RECT 1404.400 0.000 1405.200 1.000 ;
  RECT 1404.700 1.000 1404.900 5.200 ;
  RECT 1404.700 5.200 1404.960 5.400 ;
  RECT 1404.760 5.400 1404.960 7.020 ;
  RECT 1390.000 0.000 1390.800 1.000 ;
  RECT 1390.300 1.000 1390.500 5.200 ;
  RECT 1390.130 5.200 1390.500 5.400 ;
  RECT 1390.130 5.400 1390.330 7.020 ;
  RECT 1384.800 0.000 1385.600 1.000 ;
  RECT 1385.100 1.000 1385.300 5.200 ;
  RECT 1384.920 5.200 1385.300 5.400 ;
  RECT 1384.920 5.400 1385.120 7.020 ;
  RECT 1371.600 0.000 1372.400 1.000 ;
  RECT 1371.900 1.000 1372.100 5.200 ;
  RECT 1371.900 5.200 1372.210 5.400 ;
  RECT 1372.010 5.400 1372.210 7.020 ;
  RECT 1370.000 0.000 1370.800 1.000 ;
  RECT 1370.300 1.000 1370.500 5.200 ;
  RECT 1370.290 5.200 1370.500 5.400 ;
  RECT 1370.290 5.400 1370.490 7.020 ;
  RECT 1349.200 0.000 1350.000 1.000 ;
  RECT 1349.500 1.000 1349.700 5.200 ;
  RECT 1349.500 5.200 1349.720 5.400 ;
  RECT 1349.520 5.400 1349.720 7.020 ;
  RECT 1348.000 0.000 1348.800 1.000 ;
  RECT 1348.300 1.000 1348.500 5.200 ;
  RECT 1348.300 5.200 1348.570 5.400 ;
  RECT 1348.370 5.400 1348.570 7.020 ;
  RECT 1346.800 0.000 1347.600 1.000 ;
  RECT 1347.100 1.000 1347.300 5.200 ;
  RECT 1347.100 5.200 1347.400 5.400 ;
  RECT 1347.200 5.400 1347.400 7.020 ;
  RECT 1345.600 0.000 1346.400 1.000 ;
  RECT 1345.900 1.000 1346.100 5.200 ;
  RECT 1345.900 5.200 1346.150 5.400 ;
  RECT 1345.950 5.400 1346.150 7.020 ;
  RECT 1344.400 0.000 1345.200 1.000 ;
  RECT 1344.700 1.000 1344.900 5.200 ;
  RECT 1344.700 5.200 1344.900 5.400 ;
  RECT 1344.700 5.400 1344.900 7.020 ;
  RECT 1343.200 0.000 1344.000 1.000 ;
  RECT 1343.500 1.000 1343.700 5.200 ;
  RECT 1343.450 5.200 1343.700 5.400 ;
  RECT 1343.450 5.400 1343.650 7.020 ;
  RECT 1337.200 0.000 1338.000 1.000 ;
  RECT 1337.500 1.000 1337.700 5.200 ;
  RECT 1337.480 5.200 1337.700 5.400 ;
  RECT 1337.480 5.400 1337.680 7.020 ;
  RECT 1330.000 0.000 1330.800 1.000 ;
  RECT 1330.300 1.000 1330.500 5.200 ;
  RECT 1330.180 5.200 1330.500 5.400 ;
  RECT 1330.180 5.400 1330.380 7.020 ;
  RECT 1327.200 0.000 1328.000 1.000 ;
  RECT 1327.500 1.000 1327.700 5.200 ;
  RECT 1327.500 5.200 1327.900 5.400 ;
  RECT 1327.700 5.400 1327.900 7.020 ;
  RECT 1324.400 0.000 1325.200 1.000 ;
  RECT 1324.700 1.000 1324.900 5.200 ;
  RECT 1324.700 5.200 1325.040 5.400 ;
  RECT 1324.840 5.400 1325.040 7.020 ;
  RECT 1322.000 0.000 1322.800 1.000 ;
  RECT 1322.300 1.000 1322.500 5.200 ;
  RECT 1322.300 5.200 1322.560 5.400 ;
  RECT 1322.360 5.400 1322.560 7.020 ;
  RECT 1320.400 0.000 1321.200 1.000 ;
  RECT 1320.700 1.000 1320.900 5.200 ;
  RECT 1320.700 5.200 1321.040 5.400 ;
  RECT 1320.840 5.400 1321.040 7.020 ;
  RECT 1318.000 0.000 1318.800 1.000 ;
  RECT 1318.300 1.000 1318.500 5.200 ;
  RECT 1318.300 5.200 1318.560 5.400 ;
  RECT 1318.360 5.400 1318.560 7.020 ;
  RECT 1311.200 0.000 1312.000 1.000 ;
  RECT 1311.500 1.000 1311.700 5.200 ;
  RECT 1311.460 5.200 1311.700 5.400 ;
  RECT 1311.460 5.400 1311.660 7.020 ;
  RECT 1296.400 0.000 1297.200 1.000 ;
  RECT 1296.700 1.000 1296.900 5.200 ;
  RECT 1296.700 5.200 1297.030 5.400 ;
  RECT 1296.830 5.400 1297.030 7.020 ;
  RECT 1291.200 0.000 1292.000 1.000 ;
  RECT 1291.500 1.000 1291.700 5.200 ;
  RECT 1291.500 5.200 1291.820 5.400 ;
  RECT 1291.620 5.400 1291.820 7.020 ;
  RECT 1276.800 0.000 1277.600 1.000 ;
  RECT 1277.100 1.000 1277.300 5.200 ;
  RECT 1276.990 5.200 1277.300 5.400 ;
  RECT 1276.990 5.400 1277.190 7.020 ;
  RECT 1270.400 0.000 1271.200 1.000 ;
  RECT 1270.700 1.000 1270.900 5.200 ;
  RECT 1270.540 5.200 1270.900 5.400 ;
  RECT 1270.540 5.400 1270.740 7.020 ;
  RECT 1255.600 0.000 1256.400 1.000 ;
  RECT 1255.900 1.000 1256.100 5.200 ;
  RECT 1255.900 5.200 1256.110 5.400 ;
  RECT 1255.910 5.400 1256.110 7.020 ;
  RECT 1250.400 0.000 1251.200 1.000 ;
  RECT 1250.700 1.000 1250.900 5.200 ;
  RECT 1250.700 5.200 1250.900 5.400 ;
  RECT 1250.700 5.400 1250.900 7.020 ;
  RECT 1235.600 0.000 1236.400 1.000 ;
  RECT 1235.900 1.000 1236.100 5.200 ;
  RECT 1235.900 5.200 1236.270 5.400 ;
  RECT 1236.070 5.400 1236.270 7.020 ;
  RECT 1229.200 0.000 1230.000 1.000 ;
  RECT 1229.500 1.000 1229.700 5.200 ;
  RECT 1229.500 5.200 1229.820 5.400 ;
  RECT 1229.620 5.400 1229.820 7.020 ;
  RECT 1214.800 0.000 1215.600 1.000 ;
  RECT 1215.100 1.000 1215.300 5.200 ;
  RECT 1214.990 5.200 1215.300 5.400 ;
  RECT 1214.990 5.400 1215.190 7.020 ;
  RECT 1209.600 0.000 1210.400 1.000 ;
  RECT 1209.900 1.000 1210.100 5.200 ;
  RECT 1209.780 5.200 1210.100 5.400 ;
  RECT 1209.780 5.400 1209.980 7.020 ;
  RECT 1194.800 0.000 1195.600 1.000 ;
  RECT 1195.100 1.000 1195.300 5.200 ;
  RECT 1195.100 5.200 1195.350 5.400 ;
  RECT 1195.150 5.400 1195.350 7.020 ;
  RECT 1188.400 0.000 1189.200 1.000 ;
  RECT 1188.700 1.000 1188.900 5.200 ;
  RECT 1188.700 5.200 1188.900 5.400 ;
  RECT 1188.700 5.400 1188.900 7.020 ;
  RECT 1173.600 0.000 1174.400 1.000 ;
  RECT 1173.900 1.000 1174.100 5.200 ;
  RECT 1173.900 5.200 1174.270 5.400 ;
  RECT 1174.070 5.400 1174.270 7.020 ;
  RECT 1168.400 0.000 1169.200 1.000 ;
  RECT 1168.700 1.000 1168.900 5.200 ;
  RECT 1168.700 5.200 1169.060 5.400 ;
  RECT 1168.860 5.400 1169.060 7.020 ;
  RECT 1154.000 0.000 1154.800 1.000 ;
  RECT 1154.300 1.000 1154.500 5.200 ;
  RECT 1154.230 5.200 1154.500 5.400 ;
  RECT 1154.230 5.400 1154.430 7.020 ;
  RECT 1147.600 0.000 1148.400 1.000 ;
  RECT 1147.900 1.000 1148.100 5.200 ;
  RECT 1147.780 5.200 1148.100 5.400 ;
  RECT 1147.780 5.400 1147.980 7.020 ;
  RECT 1132.800 0.000 1133.600 1.000 ;
  RECT 1133.100 1.000 1133.300 5.200 ;
  RECT 1133.100 5.200 1133.350 5.400 ;
  RECT 1133.150 5.400 1133.350 7.020 ;
  RECT 1127.600 0.000 1128.400 1.000 ;
  RECT 1127.900 1.000 1128.100 5.200 ;
  RECT 1127.900 5.200 1128.140 5.400 ;
  RECT 1127.940 5.400 1128.140 7.020 ;
  RECT 1113.200 0.000 1114.000 1.000 ;
  RECT 1113.500 1.000 1113.700 5.200 ;
  RECT 1113.310 5.200 1113.700 5.400 ;
  RECT 1113.310 5.400 1113.510 7.020 ;
  RECT 1106.400 0.000 1107.200 1.000 ;
  RECT 1106.700 1.000 1106.900 5.200 ;
  RECT 1106.700 5.200 1107.060 5.400 ;
  RECT 1106.860 5.400 1107.060 7.020 ;
  RECT 1092.000 0.000 1092.800 1.000 ;
  RECT 1092.300 1.000 1092.500 5.200 ;
  RECT 1092.230 5.200 1092.500 5.400 ;
  RECT 1092.230 5.400 1092.430 7.020 ;
  RECT 1086.800 0.000 1087.600 1.000 ;
  RECT 1087.100 1.000 1087.300 5.200 ;
  RECT 1087.020 5.200 1087.300 5.400 ;
  RECT 1087.020 5.400 1087.220 7.020 ;
  RECT 1072.000 0.000 1072.800 1.000 ;
  RECT 1072.300 1.000 1072.500 5.200 ;
  RECT 1072.300 5.200 1072.590 5.400 ;
  RECT 1072.390 5.400 1072.590 7.020 ;
  RECT 1065.600 0.000 1066.400 1.000 ;
  RECT 1065.900 1.000 1066.100 5.200 ;
  RECT 1065.900 5.200 1066.140 5.400 ;
  RECT 1065.940 5.400 1066.140 7.020 ;
  RECT 1051.200 0.000 1052.000 1.000 ;
  RECT 1051.500 1.000 1051.700 5.200 ;
  RECT 1051.310 5.200 1051.700 5.400 ;
  RECT 1051.310 5.400 1051.510 7.020 ;
  RECT 1045.600 0.000 1046.400 1.000 ;
  RECT 1045.900 1.000 1046.100 5.200 ;
  RECT 1045.900 5.200 1046.300 5.400 ;
  RECT 1046.100 5.400 1046.300 7.020 ;
  RECT 1031.200 0.000 1032.000 1.000 ;
  RECT 1031.500 1.000 1031.700 5.200 ;
  RECT 1031.470 5.200 1031.700 5.400 ;
  RECT 1031.470 5.400 1031.670 7.020 ;
  RECT 1024.800 0.000 1025.600 1.000 ;
  RECT 1025.100 1.000 1025.300 5.200 ;
  RECT 1025.020 5.200 1025.300 5.400 ;
  RECT 1025.020 5.400 1025.220 7.020 ;
  RECT 1010.000 0.000 1010.800 1.000 ;
  RECT 1010.300 1.000 1010.500 5.200 ;
  RECT 1010.300 5.200 1010.590 5.400 ;
  RECT 1010.390 5.400 1010.590 7.020 ;
  RECT 1004.800 0.000 1005.600 1.000 ;
  RECT 1005.100 1.000 1005.300 5.200 ;
  RECT 1005.100 5.200 1005.380 5.400 ;
  RECT 1005.180 5.400 1005.380 7.020 ;
  RECT 992.000 0.000 992.800 1.000 ;
  RECT 992.300 1.000 992.500 5.200 ;
  RECT 992.270 5.200 992.500 5.400 ;
  RECT 992.270 5.400 992.470 7.020 ;
  RECT 990.400 0.000 991.200 1.000 ;
  RECT 990.700 1.000 990.900 5.200 ;
  RECT 990.550 5.200 990.900 5.400 ;
  RECT 990.550 5.400 990.750 7.020 ;
  RECT 983.600 0.000 984.400 1.000 ;
  RECT 983.900 1.000 984.100 5.200 ;
  RECT 983.900 5.200 984.300 5.400 ;
  RECT 984.100 5.400 984.300 7.020 ;
  RECT 969.200 0.000 970.000 1.000 ;
  RECT 969.500 1.000 969.700 5.200 ;
  RECT 969.470 5.200 969.700 5.400 ;
  RECT 969.470 5.400 969.670 7.020 ;
  RECT 964.000 0.000 964.800 1.000 ;
  RECT 964.300 1.000 964.500 5.200 ;
  RECT 964.260 5.200 964.500 5.400 ;
  RECT 964.260 5.400 964.460 7.020 ;
  RECT 949.200 0.000 950.000 1.000 ;
  RECT 949.500 1.000 949.700 5.200 ;
  RECT 949.500 5.200 949.830 5.400 ;
  RECT 949.630 5.400 949.830 7.020 ;
  RECT 942.800 0.000 943.600 1.000 ;
  RECT 943.100 1.000 943.300 5.200 ;
  RECT 943.100 5.200 943.380 5.400 ;
  RECT 943.180 5.400 943.380 7.020 ;
  RECT 928.400 0.000 929.200 1.000 ;
  RECT 928.700 1.000 928.900 5.200 ;
  RECT 928.550 5.200 928.900 5.400 ;
  RECT 928.550 5.400 928.750 7.020 ;
  RECT 923.200 0.000 924.000 1.000 ;
  RECT 923.500 1.000 923.700 5.200 ;
  RECT 923.340 5.200 923.700 5.400 ;
  RECT 923.340 5.400 923.540 7.020 ;
  RECT 908.400 0.000 909.200 1.000 ;
  RECT 908.700 1.000 908.900 5.200 ;
  RECT 908.700 5.200 908.910 5.400 ;
  RECT 908.710 5.400 908.910 7.020 ;
  RECT 902.000 0.000 902.800 1.000 ;
  RECT 902.300 1.000 902.500 5.200 ;
  RECT 902.260 5.200 902.500 5.400 ;
  RECT 902.260 5.400 902.460 7.020 ;
  RECT 887.200 0.000 888.000 1.000 ;
  RECT 887.500 1.000 887.700 5.200 ;
  RECT 887.500 5.200 887.830 5.400 ;
  RECT 887.630 5.400 887.830 7.020 ;
  RECT 882.000 0.000 882.800 1.000 ;
  RECT 882.300 1.000 882.500 5.200 ;
  RECT 882.300 5.200 882.620 5.400 ;
  RECT 882.420 5.400 882.620 7.020 ;
  RECT 867.600 0.000 868.400 1.000 ;
  RECT 867.900 1.000 868.100 5.200 ;
  RECT 867.790 5.200 868.100 5.400 ;
  RECT 867.790 5.400 867.990 7.020 ;
  RECT 861.200 0.000 862.000 1.000 ;
  RECT 861.500 1.000 861.700 5.200 ;
  RECT 861.340 5.200 861.700 5.400 ;
  RECT 861.340 5.400 861.540 7.020 ;
  RECT 846.400 0.000 847.200 1.000 ;
  RECT 846.700 1.000 846.900 5.200 ;
  RECT 846.700 5.200 846.910 5.400 ;
  RECT 846.710 5.400 846.910 7.020 ;
  RECT 841.200 0.000 842.000 1.000 ;
  RECT 841.500 1.000 841.700 5.200 ;
  RECT 841.500 5.200 841.700 5.400 ;
  RECT 841.500 5.400 841.700 7.020 ;
  RECT 826.400 0.000 827.200 1.000 ;
  RECT 826.700 1.000 826.900 5.200 ;
  RECT 826.700 5.200 827.070 5.400 ;
  RECT 826.870 5.400 827.070 7.020 ;
  RECT 820.000 0.000 820.800 1.000 ;
  RECT 820.300 1.000 820.500 5.200 ;
  RECT 820.300 5.200 820.620 5.400 ;
  RECT 820.420 5.400 820.620 7.020 ;
  RECT 805.600 0.000 806.400 1.000 ;
  RECT 805.900 1.000 806.100 5.200 ;
  RECT 805.790 5.200 806.100 5.400 ;
  RECT 805.790 5.400 805.990 7.020 ;
  RECT 800.400 0.000 801.200 1.000 ;
  RECT 800.700 1.000 800.900 5.200 ;
  RECT 800.580 5.200 800.900 5.400 ;
  RECT 800.580 5.400 800.780 7.020 ;
  RECT 785.600 0.000 786.400 1.000 ;
  RECT 785.900 1.000 786.100 5.200 ;
  RECT 785.900 5.200 786.150 5.400 ;
  RECT 785.950 5.400 786.150 7.020 ;
  RECT 779.200 0.000 780.000 1.000 ;
  RECT 779.500 1.000 779.700 5.200 ;
  RECT 779.500 5.200 779.700 5.400 ;
  RECT 779.500 5.400 779.700 7.020 ;
  RECT 764.400 0.000 765.200 1.000 ;
  RECT 764.700 1.000 764.900 5.200 ;
  RECT 764.700 5.200 765.070 5.400 ;
  RECT 764.870 5.400 765.070 7.020 ;
  RECT 759.200 0.000 760.000 1.000 ;
  RECT 759.500 1.000 759.700 5.200 ;
  RECT 759.500 5.200 759.860 5.400 ;
  RECT 759.660 5.400 759.860 7.020 ;
  RECT 744.800 0.000 745.600 1.000 ;
  RECT 745.100 1.000 745.300 5.200 ;
  RECT 745.030 5.200 745.300 5.400 ;
  RECT 745.030 5.400 745.230 7.020 ;
  RECT 738.400 0.000 739.200 1.000 ;
  RECT 738.700 1.000 738.900 5.200 ;
  RECT 738.580 5.200 738.900 5.400 ;
  RECT 738.580 5.400 738.780 7.020 ;
  RECT 723.600 0.000 724.400 1.000 ;
  RECT 723.900 1.000 724.100 5.200 ;
  RECT 723.900 5.200 724.150 5.400 ;
  RECT 723.950 5.400 724.150 7.020 ;
  RECT 718.400 0.000 719.200 1.000 ;
  RECT 718.700 1.000 718.900 5.200 ;
  RECT 718.700 5.200 718.940 5.400 ;
  RECT 718.740 5.400 718.940 7.020 ;
  RECT 704.000 0.000 704.800 1.000 ;
  RECT 704.300 1.000 704.500 5.200 ;
  RECT 704.110 5.200 704.500 5.400 ;
  RECT 704.110 5.400 704.310 7.020 ;
  RECT 697.200 0.000 698.000 1.000 ;
  RECT 697.500 1.000 697.700 5.200 ;
  RECT 697.500 5.200 697.860 5.400 ;
  RECT 697.660 5.400 697.860 7.020 ;
  RECT 682.800 0.000 683.600 1.000 ;
  RECT 683.100 1.000 683.300 5.200 ;
  RECT 683.030 5.200 683.300 5.400 ;
  RECT 683.030 5.400 683.230 7.020 ;
  RECT 677.600 0.000 678.400 1.000 ;
  RECT 677.900 1.000 678.100 5.200 ;
  RECT 677.820 5.200 678.100 5.400 ;
  RECT 677.820 5.400 678.020 7.020 ;
  RECT 664.800 0.000 665.600 1.000 ;
  RECT 665.100 1.000 665.300 5.200 ;
  RECT 664.910 5.200 665.300 5.400 ;
  RECT 664.910 5.400 665.110 7.020 ;
  RECT 662.800 0.000 663.600 1.000 ;
  RECT 663.100 1.000 663.300 5.200 ;
  RECT 663.100 5.200 663.390 5.400 ;
  RECT 663.190 5.400 663.390 7.020 ;
  RECT 656.400 0.000 657.200 1.000 ;
  RECT 656.700 1.000 656.900 5.200 ;
  RECT 656.700 5.200 656.940 5.400 ;
  RECT 656.740 5.400 656.940 7.020 ;
  RECT 642.000 0.000 642.800 1.000 ;
  RECT 642.300 1.000 642.500 5.200 ;
  RECT 642.110 5.200 642.500 5.400 ;
  RECT 642.110 5.400 642.310 7.020 ;
  RECT 636.400 0.000 637.200 1.000 ;
  RECT 636.700 1.000 636.900 5.200 ;
  RECT 636.700 5.200 637.100 5.400 ;
  RECT 636.900 5.400 637.100 7.020 ;
  RECT 622.000 0.000 622.800 1.000 ;
  RECT 622.300 1.000 622.500 5.200 ;
  RECT 622.270 5.200 622.500 5.400 ;
  RECT 622.270 5.400 622.470 7.020 ;
  RECT 615.600 0.000 616.400 1.000 ;
  RECT 615.900 1.000 616.100 5.200 ;
  RECT 615.820 5.200 616.100 5.400 ;
  RECT 615.820 5.400 616.020 7.020 ;
  RECT 600.800 0.000 601.600 1.000 ;
  RECT 601.100 1.000 601.300 5.200 ;
  RECT 601.100 5.200 601.390 5.400 ;
  RECT 601.190 5.400 601.390 7.020 ;
  RECT 595.600 0.000 596.400 1.000 ;
  RECT 595.900 1.000 596.100 5.200 ;
  RECT 595.900 5.200 596.180 5.400 ;
  RECT 595.980 5.400 596.180 7.020 ;
  RECT 581.200 0.000 582.000 1.000 ;
  RECT 581.500 1.000 581.700 5.200 ;
  RECT 581.350 5.200 581.700 5.400 ;
  RECT 581.350 5.400 581.550 7.020 ;
  RECT 574.400 0.000 575.200 1.000 ;
  RECT 574.700 1.000 574.900 5.200 ;
  RECT 574.700 5.200 575.100 5.400 ;
  RECT 574.900 5.400 575.100 7.020 ;
  RECT 560.000 0.000 560.800 1.000 ;
  RECT 560.300 1.000 560.500 5.200 ;
  RECT 560.270 5.200 560.500 5.400 ;
  RECT 560.270 5.400 560.470 7.020 ;
  RECT 554.800 0.000 555.600 1.000 ;
  RECT 555.100 1.000 555.300 5.200 ;
  RECT 555.060 5.200 555.300 5.400 ;
  RECT 555.060 5.400 555.260 7.020 ;
  RECT 540.000 0.000 540.800 1.000 ;
  RECT 540.300 1.000 540.500 5.200 ;
  RECT 540.300 5.200 540.630 5.400 ;
  RECT 540.430 5.400 540.630 7.020 ;
  RECT 533.600 0.000 534.400 1.000 ;
  RECT 533.900 1.000 534.100 5.200 ;
  RECT 533.900 5.200 534.180 5.400 ;
  RECT 533.980 5.400 534.180 7.020 ;
  RECT 519.200 0.000 520.000 1.000 ;
  RECT 519.500 1.000 519.700 5.200 ;
  RECT 519.350 5.200 519.700 5.400 ;
  RECT 519.350 5.400 519.550 7.020 ;
  RECT 514.000 0.000 514.800 1.000 ;
  RECT 514.300 1.000 514.500 5.200 ;
  RECT 514.140 5.200 514.500 5.400 ;
  RECT 514.140 5.400 514.340 7.020 ;
  RECT 499.200 0.000 500.000 1.000 ;
  RECT 499.500 1.000 499.700 5.200 ;
  RECT 499.500 5.200 499.710 5.400 ;
  RECT 499.510 5.400 499.710 7.020 ;
  RECT 492.800 0.000 493.600 1.000 ;
  RECT 493.100 1.000 493.300 5.200 ;
  RECT 493.060 5.200 493.300 5.400 ;
  RECT 493.060 5.400 493.260 7.020 ;
  RECT 478.000 0.000 478.800 1.000 ;
  RECT 478.300 1.000 478.500 5.200 ;
  RECT 478.300 5.200 478.630 5.400 ;
  RECT 478.430 5.400 478.630 7.020 ;
  RECT 472.800 0.000 473.600 1.000 ;
  RECT 473.100 1.000 473.300 5.200 ;
  RECT 473.100 5.200 473.420 5.400 ;
  RECT 473.220 5.400 473.420 7.020 ;
  RECT 458.400 0.000 459.200 1.000 ;
  RECT 458.700 1.000 458.900 5.200 ;
  RECT 458.590 5.200 458.900 5.400 ;
  RECT 458.590 5.400 458.790 7.020 ;
  RECT 452.000 0.000 452.800 1.000 ;
  RECT 452.300 1.000 452.500 5.200 ;
  RECT 452.140 5.200 452.500 5.400 ;
  RECT 452.140 5.400 452.340 7.020 ;
  RECT 437.200 0.000 438.000 1.000 ;
  RECT 437.500 1.000 437.700 5.200 ;
  RECT 437.500 5.200 437.710 5.400 ;
  RECT 437.510 5.400 437.710 7.020 ;
  RECT 432.000 0.000 432.800 1.000 ;
  RECT 432.300 1.000 432.500 5.200 ;
  RECT 432.300 5.200 432.500 5.400 ;
  RECT 432.300 5.400 432.500 7.020 ;
  RECT 417.200 0.000 418.000 1.000 ;
  RECT 417.500 1.000 417.700 5.200 ;
  RECT 417.500 5.200 417.870 5.400 ;
  RECT 417.670 5.400 417.870 7.020 ;
  RECT 410.800 0.000 411.600 1.000 ;
  RECT 411.100 1.000 411.300 5.200 ;
  RECT 411.100 5.200 411.420 5.400 ;
  RECT 411.220 5.400 411.420 7.020 ;
  RECT 396.400 0.000 397.200 1.000 ;
  RECT 396.700 1.000 396.900 5.200 ;
  RECT 396.590 5.200 396.900 5.400 ;
  RECT 396.590 5.400 396.790 7.020 ;
  RECT 391.200 0.000 392.000 1.000 ;
  RECT 391.500 1.000 391.700 5.200 ;
  RECT 391.380 5.200 391.700 5.400 ;
  RECT 391.380 5.400 391.580 7.020 ;
  RECT 376.400 0.000 377.200 1.000 ;
  RECT 376.700 1.000 376.900 5.200 ;
  RECT 376.700 5.200 376.950 5.400 ;
  RECT 376.750 5.400 376.950 7.020 ;
  RECT 370.000 0.000 370.800 1.000 ;
  RECT 370.300 1.000 370.500 5.200 ;
  RECT 370.300 5.200 370.500 5.400 ;
  RECT 370.300 5.400 370.500 7.020 ;
  RECT 355.200 0.000 356.000 1.000 ;
  RECT 355.500 1.000 355.700 5.200 ;
  RECT 355.500 5.200 355.870 5.400 ;
  RECT 355.670 5.400 355.870 7.020 ;
  RECT 350.000 0.000 350.800 1.000 ;
  RECT 350.300 1.000 350.500 5.200 ;
  RECT 350.300 5.200 350.660 5.400 ;
  RECT 350.460 5.400 350.660 7.020 ;
  RECT 337.200 0.000 338.000 1.000 ;
  RECT 337.500 1.000 337.700 5.200 ;
  RECT 337.500 5.200 337.750 5.400 ;
  RECT 337.550 5.400 337.750 7.020 ;
  RECT 335.600 0.000 336.400 1.000 ;
  RECT 335.900 1.000 336.100 5.200 ;
  RECT 335.830 5.200 336.100 5.400 ;
  RECT 335.830 5.400 336.030 7.020 ;
  RECT 329.200 0.000 330.000 1.000 ;
  RECT 329.500 1.000 329.700 5.200 ;
  RECT 329.380 5.200 329.700 5.400 ;
  RECT 329.380 5.400 329.580 7.020 ;
  RECT 314.400 0.000 315.200 1.000 ;
  RECT 314.700 1.000 314.900 5.200 ;
  RECT 314.700 5.200 314.950 5.400 ;
  RECT 314.750 5.400 314.950 7.020 ;
  RECT 309.200 0.000 310.000 1.000 ;
  RECT 309.500 1.000 309.700 5.200 ;
  RECT 309.500 5.200 309.740 5.400 ;
  RECT 309.540 5.400 309.740 7.020 ;
  RECT 294.800 0.000 295.600 1.000 ;
  RECT 295.100 1.000 295.300 5.200 ;
  RECT 294.910 5.200 295.300 5.400 ;
  RECT 294.910 5.400 295.110 7.020 ;
  RECT 288.000 0.000 288.800 1.000 ;
  RECT 288.300 1.000 288.500 5.200 ;
  RECT 288.300 5.200 288.660 5.400 ;
  RECT 288.460 5.400 288.660 7.020 ;
  RECT 273.600 0.000 274.400 1.000 ;
  RECT 273.900 1.000 274.100 5.200 ;
  RECT 273.830 5.200 274.100 5.400 ;
  RECT 273.830 5.400 274.030 7.020 ;
  RECT 268.400 0.000 269.200 1.000 ;
  RECT 268.700 1.000 268.900 5.200 ;
  RECT 268.620 5.200 268.900 5.400 ;
  RECT 268.620 5.400 268.820 7.020 ;
  RECT 253.600 0.000 254.400 1.000 ;
  RECT 253.900 1.000 254.100 5.200 ;
  RECT 253.900 5.200 254.190 5.400 ;
  RECT 253.990 5.400 254.190 7.020 ;
  RECT 247.200 0.000 248.000 1.000 ;
  RECT 247.500 1.000 247.700 5.200 ;
  RECT 247.500 5.200 247.740 5.400 ;
  RECT 247.540 5.400 247.740 7.020 ;
  RECT 232.800 0.000 233.600 1.000 ;
  RECT 233.100 1.000 233.300 5.200 ;
  RECT 232.910 5.200 233.300 5.400 ;
  RECT 232.910 5.400 233.110 7.020 ;
  RECT 227.200 0.000 228.000 1.000 ;
  RECT 227.500 1.000 227.700 5.200 ;
  RECT 227.500 5.200 227.900 5.400 ;
  RECT 227.700 5.400 227.900 7.020 ;
  RECT 212.800 0.000 213.600 1.000 ;
  RECT 213.100 1.000 213.300 5.200 ;
  RECT 213.070 5.200 213.300 5.400 ;
  RECT 213.070 5.400 213.270 7.020 ;
  RECT 206.400 0.000 207.200 1.000 ;
  RECT 206.700 1.000 206.900 5.200 ;
  RECT 206.620 5.200 206.900 5.400 ;
  RECT 206.620 5.400 206.820 7.020 ;
  RECT 191.600 0.000 192.400 1.000 ;
  RECT 191.900 1.000 192.100 5.200 ;
  RECT 191.900 5.200 192.190 5.400 ;
  RECT 191.990 5.400 192.190 7.020 ;
  RECT 186.400 0.000 187.200 1.000 ;
  RECT 186.700 1.000 186.900 5.200 ;
  RECT 186.700 5.200 186.980 5.400 ;
  RECT 186.780 5.400 186.980 7.020 ;
  RECT 172.000 0.000 172.800 1.000 ;
  RECT 172.300 1.000 172.500 5.200 ;
  RECT 172.150 5.200 172.500 5.400 ;
  RECT 172.150 5.400 172.350 7.020 ;
  RECT 165.200 0.000 166.000 1.000 ;
  RECT 165.500 1.000 165.700 5.200 ;
  RECT 165.500 5.200 165.900 5.400 ;
  RECT 165.700 5.400 165.900 7.020 ;
  RECT 150.800 0.000 151.600 1.000 ;
  RECT 151.100 1.000 151.300 5.200 ;
  RECT 151.070 5.200 151.300 5.400 ;
  RECT 151.070 5.400 151.270 7.020 ;
  RECT 145.600 0.000 146.400 1.000 ;
  RECT 145.900 1.000 146.100 5.200 ;
  RECT 145.860 5.200 146.100 5.400 ;
  RECT 145.860 5.400 146.060 7.020 ;
  RECT 130.800 0.000 131.600 1.000 ;
  RECT 131.100 1.000 131.300 5.200 ;
  RECT 131.100 5.200 131.430 5.400 ;
  RECT 131.230 5.400 131.430 7.020 ;
  RECT 124.400 0.000 125.200 1.000 ;
  RECT 124.700 1.000 124.900 5.200 ;
  RECT 124.700 5.200 124.980 5.400 ;
  RECT 124.780 5.400 124.980 7.020 ;
  RECT 110.000 0.000 110.800 1.000 ;
  RECT 110.300 1.000 110.500 5.200 ;
  RECT 110.150 5.200 110.500 5.400 ;
  RECT 110.150 5.400 110.350 7.020 ;
  RECT 104.800 0.000 105.600 1.000 ;
  RECT 105.100 1.000 105.300 5.200 ;
  RECT 104.940 5.200 105.300 5.400 ;
  RECT 104.940 5.400 105.140 7.020 ;
  RECT 90.000 0.000 90.800 1.000 ;
  RECT 90.300 1.000 90.500 5.200 ;
  RECT 90.300 5.200 90.510 5.400 ;
  RECT 90.310 5.400 90.510 7.020 ;
  RECT 83.600 0.000 84.400 1.000 ;
  RECT 83.900 1.000 84.100 5.200 ;
  RECT 83.860 5.200 84.100 5.400 ;
  RECT 83.860 5.400 84.060 7.020 ;
  RECT 68.800 0.000 69.600 1.000 ;
  RECT 69.100 1.000 69.300 5.200 ;
  RECT 69.100 5.200 69.430 5.400 ;
  RECT 69.230 5.400 69.430 7.020 ;
  RECT 63.600 0.000 64.400 1.000 ;
  RECT 63.900 1.000 64.100 5.200 ;
  RECT 63.900 5.200 64.220 5.400 ;
  RECT 64.020 5.400 64.220 7.020 ;
  RECT 49.200 0.000 50.000 1.000 ;
  RECT 49.500 1.000 49.700 5.200 ;
  RECT 49.390 5.200 49.700 5.400 ;
  RECT 49.390 5.400 49.590 7.020 ;
  RECT 42.800 0.000 43.600 1.000 ;
  RECT 43.100 1.000 43.300 5.200 ;
  RECT 42.940 5.200 43.300 5.400 ;
  RECT 42.940 5.400 43.140 7.020 ;
  RECT 28.000 0.000 28.800 1.000 ;
  RECT 28.300 1.000 28.500 5.200 ;
  RECT 28.300 5.200 28.510 5.400 ;
  RECT 28.310 5.400 28.510 7.020 ;
  RECT 22.800 0.000 23.600 1.000 ;
  RECT 23.100 1.000 23.300 5.200 ;
  RECT 23.100 5.200 23.300 5.400 ;
  RECT 23.100 5.400 23.300 7.020 ;
  RECT 10.000 0.000 10.800 1.000 ;
  RECT 10.300 1.000 10.500 5.200 ;
  RECT 10.190 5.200 10.500 5.400 ;
  RECT 10.190 5.400 10.390 7.020 ;
  RECT 8.000 0.000 8.800 1.000 ;
  RECT 8.300 1.000 8.500 5.200 ;
  RECT 8.300 5.200 8.670 5.400 ;
  RECT 8.470 5.400 8.670 7.020 ;
  RECT 2679.520 9.570 2680.660 11.170 ;
  RECT 2679.520 14.200 2680.660 15.200 ;
  RECT 2679.520 18.730 2680.660 19.730 ;
  RECT 2679.520 21.230 2680.660 22.070 ;
  RECT 2679.520 24.170 2680.660 25.170 ;
  RECT 2679.520 36.320 2680.660 37.320 ;
  RECT 2679.520 39.480 2680.660 40.080 ;
  RECT 2679.520 45.560 2680.660 46.160 ;
  RECT 2679.520 57.100 2680.660 61.420 ;
  RECT 4.280 57.100 5.420 61.420 ;
  RECT 4.280 45.560 5.420 46.160 ;
  RECT 4.280 39.480 5.420 40.080 ;
  RECT 4.280 36.320 5.420 37.320 ;
  RECT 4.280 24.170 5.420 25.170 ;
  RECT 4.280 21.230 5.420 22.070 ;
  RECT 4.280 18.730 5.420 19.730 ;
  RECT 4.280 14.200 5.420 15.200 ;
  RECT 4.280 9.570 5.420 11.170 ;
  RECT 2679.520 191.940 2680.660 192.320 ;
  RECT 2679.520 184.020 2680.660 184.300 ;
  RECT 2679.520 180.340 2680.660 180.620 ;
  RECT 2679.520 176.660 2680.660 176.940 ;
  RECT 2679.520 172.980 2680.660 173.260 ;
  RECT 2679.520 169.300 2680.660 169.580 ;
  RECT 2679.520 165.620 2680.660 165.900 ;
  RECT 2679.520 161.940 2680.660 162.220 ;
  RECT 2679.520 158.260 2680.660 158.540 ;
  RECT 2679.520 154.580 2680.660 154.860 ;
  RECT 2679.520 150.900 2680.660 151.180 ;
  RECT 2679.520 147.220 2680.660 147.500 ;
  RECT 2679.520 143.540 2680.660 143.820 ;
  RECT 2679.520 139.860 2680.660 140.140 ;
  RECT 2679.520 136.180 2680.660 136.460 ;
  RECT 2679.520 132.500 2680.660 132.780 ;
  RECT 2679.520 128.820 2680.660 129.100 ;
  RECT 2679.520 125.140 2680.660 125.420 ;
  RECT 2679.520 121.460 2680.660 121.740 ;
  RECT 2679.520 117.780 2680.660 118.060 ;
  RECT 2679.520 114.100 2680.660 114.380 ;
  RECT 2679.520 110.420 2680.660 110.700 ;
  RECT 2679.520 106.740 2680.660 107.020 ;
  RECT 2679.520 103.060 2680.660 103.340 ;
  RECT 2679.520 99.380 2680.660 99.660 ;
  RECT 2679.520 95.700 2680.660 95.980 ;
  RECT 2679.520 92.020 2680.660 92.300 ;
  RECT 2679.520 88.340 2680.660 88.620 ;
  RECT 2679.520 84.660 2680.660 84.940 ;
  RECT 2679.520 80.980 2680.660 81.260 ;
  RECT 2679.520 77.300 2680.660 77.580 ;
  RECT 2679.520 73.620 2680.660 73.900 ;
  RECT 2679.520 69.940 2680.660 70.220 ;
  RECT 2679.520 65.600 2680.660 65.980 ;
  RECT 1368.820 192.510 1369.070 193.650 ;
  RECT 1409.740 192.510 1409.990 193.650 ;
  RECT 1450.660 192.510 1450.910 193.650 ;
  RECT 1491.580 192.510 1491.830 193.650 ;
  RECT 1532.500 192.510 1532.750 193.650 ;
  RECT 1573.420 192.510 1573.670 193.650 ;
  RECT 1614.340 192.510 1614.590 193.650 ;
  RECT 1655.260 192.510 1655.510 193.650 ;
  RECT 1696.180 192.510 1696.430 193.650 ;
  RECT 1737.100 192.510 1737.350 193.650 ;
  RECT 1778.020 192.510 1778.270 193.650 ;
  RECT 1818.940 192.510 1819.190 193.650 ;
  RECT 1859.860 192.510 1860.110 193.650 ;
  RECT 1900.780 192.510 1901.030 193.650 ;
  RECT 1941.700 192.510 1941.950 193.650 ;
  RECT 1982.620 192.510 1982.870 193.650 ;
  RECT 2023.540 192.510 2023.790 193.650 ;
  RECT 2064.460 192.510 2064.710 193.650 ;
  RECT 2105.380 192.510 2105.630 193.650 ;
  RECT 2146.300 192.510 2146.550 193.650 ;
  RECT 2187.220 192.510 2187.470 193.650 ;
  RECT 2228.140 192.510 2228.390 193.650 ;
  RECT 2269.060 192.510 2269.310 193.650 ;
  RECT 2309.980 192.510 2310.230 193.650 ;
  RECT 2350.900 192.510 2351.150 193.650 ;
  RECT 2391.820 192.510 2392.070 193.650 ;
  RECT 2432.740 192.510 2432.990 193.650 ;
  RECT 2473.660 192.510 2473.910 193.650 ;
  RECT 2514.580 192.510 2514.830 193.650 ;
  RECT 2555.500 192.510 2555.750 193.650 ;
  RECT 2596.420 192.510 2596.670 193.650 ;
  RECT 2637.340 192.510 2637.590 193.650 ;
  RECT 1351.810 192.510 1354.320 193.650 ;
  RECT 1339.390 192.510 1341.780 193.650 ;
  RECT 1331.880 192.510 1334.940 193.650 ;
  RECT 1356.060 192.510 1358.910 193.650 ;
  RECT 1360.360 192.510 1363.610 193.650 ;
  RECT 1329.160 192.510 1330.920 193.650 ;
  RECT 1319.820 192.510 1321.580 193.650 ;
  RECT 1323.820 192.510 1325.580 193.650 ;
  RECT 4.280 65.600 5.420 65.980 ;
  RECT 4.280 69.940 5.420 70.220 ;
  RECT 4.280 73.620 5.420 73.900 ;
  RECT 4.280 77.300 5.420 77.580 ;
  RECT 4.280 80.980 5.420 81.260 ;
  RECT 4.280 84.660 5.420 84.940 ;
  RECT 4.280 88.340 5.420 88.620 ;
  RECT 4.280 92.020 5.420 92.300 ;
  RECT 4.280 95.700 5.420 95.980 ;
  RECT 4.280 99.380 5.420 99.660 ;
  RECT 4.280 103.060 5.420 103.340 ;
  RECT 4.280 106.740 5.420 107.020 ;
  RECT 4.280 110.420 5.420 110.700 ;
  RECT 4.280 114.100 5.420 114.380 ;
  RECT 4.280 117.780 5.420 118.060 ;
  RECT 4.280 121.460 5.420 121.740 ;
  RECT 4.280 125.140 5.420 125.420 ;
  RECT 4.280 128.820 5.420 129.100 ;
  RECT 4.280 132.500 5.420 132.780 ;
  RECT 4.280 136.180 5.420 136.460 ;
  RECT 4.280 139.860 5.420 140.140 ;
  RECT 4.280 143.540 5.420 143.820 ;
  RECT 4.280 147.220 5.420 147.500 ;
  RECT 4.280 150.900 5.420 151.180 ;
  RECT 4.280 154.580 5.420 154.860 ;
  RECT 4.280 158.260 5.420 158.540 ;
  RECT 4.280 161.940 5.420 162.220 ;
  RECT 4.280 165.620 5.420 165.900 ;
  RECT 4.280 169.300 5.420 169.580 ;
  RECT 4.280 172.980 5.420 173.260 ;
  RECT 4.280 176.660 5.420 176.940 ;
  RECT 4.280 180.340 5.420 180.620 ;
  RECT 4.280 184.020 5.420 184.300 ;
  RECT 4.280 191.940 5.420 192.320 ;
  RECT 47.350 192.510 47.600 193.650 ;
  RECT 88.270 192.510 88.520 193.650 ;
  RECT 129.190 192.510 129.440 193.650 ;
  RECT 170.110 192.510 170.360 193.650 ;
  RECT 211.030 192.510 211.280 193.650 ;
  RECT 251.950 192.510 252.200 193.650 ;
  RECT 292.870 192.510 293.120 193.650 ;
  RECT 333.790 192.510 334.040 193.650 ;
  RECT 374.710 192.510 374.960 193.650 ;
  RECT 415.630 192.510 415.880 193.650 ;
  RECT 456.550 192.510 456.800 193.650 ;
  RECT 497.470 192.510 497.720 193.650 ;
  RECT 538.390 192.510 538.640 193.650 ;
  RECT 579.310 192.510 579.560 193.650 ;
  RECT 620.230 192.510 620.480 193.650 ;
  RECT 661.150 192.510 661.400 193.650 ;
  RECT 702.070 192.510 702.320 193.650 ;
  RECT 742.990 192.510 743.240 193.650 ;
  RECT 783.910 192.510 784.160 193.650 ;
  RECT 824.830 192.510 825.080 193.650 ;
  RECT 865.750 192.510 866.000 193.650 ;
  RECT 906.670 192.510 906.920 193.650 ;
  RECT 947.590 192.510 947.840 193.650 ;
  RECT 988.510 192.510 988.760 193.650 ;
  RECT 1029.430 192.510 1029.680 193.650 ;
  RECT 1070.350 192.510 1070.600 193.650 ;
  RECT 1111.270 192.510 1111.520 193.650 ;
  RECT 1152.190 192.510 1152.440 193.650 ;
  RECT 1193.110 192.510 1193.360 193.650 ;
  RECT 1234.030 192.510 1234.280 193.650 ;
  RECT 1274.950 192.510 1275.200 193.650 ;
  LAYER ME1 ;
  RECT 5.420 7.020 2679.520 192.510 ;
  RECT 2683.080 3.460 2684.940 196.070 ;
  RECT 0.000 3.460 1.860 196.070 ;
  RECT 1.860 196.070 2683.080 197.930 ;
  RECT 1.860 1.600 2683.080 3.460 ;
  RECT 2680.940 5.600 2682.800 193.930 ;
  RECT 2.140 5.600 4.000 193.930 ;
  RECT 4.000 193.930 2680.940 195.790 ;
  RECT 4.000 3.740 2680.940 5.600 ;
  RECT 2.140 193.930 4.000 195.790 ;
  RECT 0.000 196.070 1.860 197.930 ;
  RECT 2680.940 3.740 2682.800 5.600 ;
  RECT 2683.080 1.600 2684.940 3.460 ;
  RECT 2680.940 193.930 2682.800 195.790 ;
  RECT 2683.080 196.070 2684.940 197.930 ;
  RECT 2.140 3.740 4.000 5.600 ;
  RECT 0.000 1.600 1.860 3.460 ;
  RECT 2672.800 0.000 2673.600 1.000 ;
  RECT 2658.400 0.000 2659.200 1.000 ;
  RECT 2653.200 0.000 2654.000 1.000 ;
  RECT 2638.400 0.000 2639.200 1.000 ;
  RECT 2632.000 0.000 2632.800 1.000 ;
  RECT 2617.600 0.000 2618.400 1.000 ;
  RECT 2612.400 0.000 2613.200 1.000 ;
  RECT 2597.600 0.000 2598.400 1.000 ;
  RECT 2591.200 0.000 2592.000 1.000 ;
  RECT 2576.400 0.000 2577.200 1.000 ;
  RECT 2571.200 0.000 2572.000 1.000 ;
  RECT 2556.800 0.000 2557.600 1.000 ;
  RECT 2550.400 0.000 2551.200 1.000 ;
  RECT 2535.600 0.000 2536.400 1.000 ;
  RECT 2530.400 0.000 2531.200 1.000 ;
  RECT 2515.600 0.000 2516.400 1.000 ;
  RECT 2509.200 0.000 2510.000 1.000 ;
  RECT 2494.800 0.000 2495.600 1.000 ;
  RECT 2489.600 0.000 2490.400 1.000 ;
  RECT 2474.800 0.000 2475.600 1.000 ;
  RECT 2468.400 0.000 2469.200 1.000 ;
  RECT 2453.600 0.000 2454.400 1.000 ;
  RECT 2448.400 0.000 2449.200 1.000 ;
  RECT 2434.000 0.000 2434.800 1.000 ;
  RECT 2427.600 0.000 2428.400 1.000 ;
  RECT 2412.800 0.000 2413.600 1.000 ;
  RECT 2407.600 0.000 2408.400 1.000 ;
  RECT 2392.800 0.000 2393.600 1.000 ;
  RECT 2386.400 0.000 2387.200 1.000 ;
  RECT 2372.000 0.000 2372.800 1.000 ;
  RECT 2366.800 0.000 2367.600 1.000 ;
  RECT 2353.600 0.000 2354.400 1.000 ;
  RECT 2352.000 0.000 2352.800 1.000 ;
  RECT 2345.600 0.000 2346.400 1.000 ;
  RECT 2330.800 0.000 2331.600 1.000 ;
  RECT 2325.600 0.000 2326.400 1.000 ;
  RECT 2311.200 0.000 2312.000 1.000 ;
  RECT 2304.800 0.000 2305.600 1.000 ;
  RECT 2290.000 0.000 2290.800 1.000 ;
  RECT 2284.800 0.000 2285.600 1.000 ;
  RECT 2270.400 0.000 2271.200 1.000 ;
  RECT 2263.600 0.000 2264.400 1.000 ;
  RECT 2249.200 0.000 2250.000 1.000 ;
  RECT 2244.000 0.000 2244.800 1.000 ;
  RECT 2229.200 0.000 2230.000 1.000 ;
  RECT 2222.800 0.000 2223.600 1.000 ;
  RECT 2208.400 0.000 2209.200 1.000 ;
  RECT 2203.200 0.000 2204.000 1.000 ;
  RECT 2188.400 0.000 2189.200 1.000 ;
  RECT 2182.000 0.000 2182.800 1.000 ;
  RECT 2167.200 0.000 2168.000 1.000 ;
  RECT 2162.000 0.000 2162.800 1.000 ;
  RECT 2147.600 0.000 2148.400 1.000 ;
  RECT 2141.200 0.000 2142.000 1.000 ;
  RECT 2126.400 0.000 2127.200 1.000 ;
  RECT 2121.200 0.000 2122.000 1.000 ;
  RECT 2106.400 0.000 2107.200 1.000 ;
  RECT 2100.000 0.000 2100.800 1.000 ;
  RECT 2085.600 0.000 2086.400 1.000 ;
  RECT 2080.400 0.000 2081.200 1.000 ;
  RECT 2065.600 0.000 2066.400 1.000 ;
  RECT 2059.200 0.000 2060.000 1.000 ;
  RECT 2044.400 0.000 2045.200 1.000 ;
  RECT 2039.200 0.000 2040.000 1.000 ;
  RECT 2026.400 0.000 2027.200 1.000 ;
  RECT 2024.800 0.000 2025.600 1.000 ;
  RECT 2018.400 0.000 2019.200 1.000 ;
  RECT 2003.600 0.000 2004.400 1.000 ;
  RECT 1998.400 0.000 1999.200 1.000 ;
  RECT 1983.600 0.000 1984.400 1.000 ;
  RECT 1977.200 0.000 1978.000 1.000 ;
  RECT 1962.800 0.000 1963.600 1.000 ;
  RECT 1957.600 0.000 1958.400 1.000 ;
  RECT 1942.800 0.000 1943.600 1.000 ;
  RECT 1936.400 0.000 1937.200 1.000 ;
  RECT 1921.600 0.000 1922.400 1.000 ;
  RECT 1916.400 0.000 1917.200 1.000 ;
  RECT 1902.000 0.000 1902.800 1.000 ;
  RECT 1895.600 0.000 1896.400 1.000 ;
  RECT 1880.800 0.000 1881.600 1.000 ;
  RECT 1875.600 0.000 1876.400 1.000 ;
  RECT 1861.200 0.000 1862.000 1.000 ;
  RECT 1854.400 0.000 1855.200 1.000 ;
  RECT 1840.000 0.000 1840.800 1.000 ;
  RECT 1834.800 0.000 1835.600 1.000 ;
  RECT 1820.000 0.000 1820.800 1.000 ;
  RECT 1813.600 0.000 1814.400 1.000 ;
  RECT 1799.200 0.000 1800.000 1.000 ;
  RECT 1794.000 0.000 1794.800 1.000 ;
  RECT 1779.200 0.000 1780.000 1.000 ;
  RECT 1772.800 0.000 1773.600 1.000 ;
  RECT 1758.000 0.000 1758.800 1.000 ;
  RECT 1752.800 0.000 1753.600 1.000 ;
  RECT 1738.400 0.000 1739.200 1.000 ;
  RECT 1732.000 0.000 1732.800 1.000 ;
  RECT 1717.200 0.000 1718.000 1.000 ;
  RECT 1712.000 0.000 1712.800 1.000 ;
  RECT 1699.200 0.000 1700.000 1.000 ;
  RECT 1697.200 0.000 1698.000 1.000 ;
  RECT 1690.800 0.000 1691.600 1.000 ;
  RECT 1676.400 0.000 1677.200 1.000 ;
  RECT 1671.200 0.000 1672.000 1.000 ;
  RECT 1656.400 0.000 1657.200 1.000 ;
  RECT 1650.000 0.000 1650.800 1.000 ;
  RECT 1635.200 0.000 1636.000 1.000 ;
  RECT 1630.000 0.000 1630.800 1.000 ;
  RECT 1615.600 0.000 1616.400 1.000 ;
  RECT 1609.200 0.000 1610.000 1.000 ;
  RECT 1594.400 0.000 1595.200 1.000 ;
  RECT 1589.200 0.000 1590.000 1.000 ;
  RECT 1574.400 0.000 1575.200 1.000 ;
  RECT 1568.000 0.000 1568.800 1.000 ;
  RECT 1553.600 0.000 1554.400 1.000 ;
  RECT 1548.400 0.000 1549.200 1.000 ;
  RECT 1533.600 0.000 1534.400 1.000 ;
  RECT 1527.200 0.000 1528.000 1.000 ;
  RECT 1512.400 0.000 1513.200 1.000 ;
  RECT 1507.200 0.000 1508.000 1.000 ;
  RECT 1492.800 0.000 1493.600 1.000 ;
  RECT 1486.400 0.000 1487.200 1.000 ;
  RECT 1471.600 0.000 1472.400 1.000 ;
  RECT 1466.400 0.000 1467.200 1.000 ;
  RECT 1452.000 0.000 1452.800 1.000 ;
  RECT 1445.200 0.000 1446.000 1.000 ;
  RECT 1430.800 0.000 1431.600 1.000 ;
  RECT 1425.600 0.000 1426.400 1.000 ;
  RECT 1410.800 0.000 1411.600 1.000 ;
  RECT 1404.400 0.000 1405.200 1.000 ;
  RECT 1390.000 0.000 1390.800 1.000 ;
  RECT 1384.800 0.000 1385.600 1.000 ;
  RECT 1371.600 0.000 1372.400 1.000 ;
  RECT 1370.000 0.000 1370.800 1.000 ;
  RECT 1349.200 0.000 1350.000 1.000 ;
  RECT 1348.000 0.000 1348.800 1.000 ;
  RECT 1346.800 0.000 1347.600 1.000 ;
  RECT 1345.600 0.000 1346.400 1.000 ;
  RECT 1344.400 0.000 1345.200 1.000 ;
  RECT 1343.200 0.000 1344.000 1.000 ;
  RECT 1337.200 0.000 1338.000 1.000 ;
  RECT 1330.000 0.000 1330.800 1.000 ;
  RECT 1327.200 0.000 1328.000 1.000 ;
  RECT 1324.400 0.000 1325.200 1.000 ;
  RECT 1322.000 0.000 1322.800 1.000 ;
  RECT 1320.400 0.000 1321.200 1.000 ;
  RECT 1318.000 0.000 1318.800 1.000 ;
  RECT 1311.200 0.000 1312.000 1.000 ;
  RECT 1296.400 0.000 1297.200 1.000 ;
  RECT 1291.200 0.000 1292.000 1.000 ;
  RECT 1276.800 0.000 1277.600 1.000 ;
  RECT 1270.400 0.000 1271.200 1.000 ;
  RECT 1255.600 0.000 1256.400 1.000 ;
  RECT 1250.400 0.000 1251.200 1.000 ;
  RECT 1235.600 0.000 1236.400 1.000 ;
  RECT 1229.200 0.000 1230.000 1.000 ;
  RECT 1214.800 0.000 1215.600 1.000 ;
  RECT 1209.600 0.000 1210.400 1.000 ;
  RECT 1194.800 0.000 1195.600 1.000 ;
  RECT 1188.400 0.000 1189.200 1.000 ;
  RECT 1173.600 0.000 1174.400 1.000 ;
  RECT 1168.400 0.000 1169.200 1.000 ;
  RECT 1154.000 0.000 1154.800 1.000 ;
  RECT 1147.600 0.000 1148.400 1.000 ;
  RECT 1132.800 0.000 1133.600 1.000 ;
  RECT 1127.600 0.000 1128.400 1.000 ;
  RECT 1113.200 0.000 1114.000 1.000 ;
  RECT 1106.400 0.000 1107.200 1.000 ;
  RECT 1092.000 0.000 1092.800 1.000 ;
  RECT 1086.800 0.000 1087.600 1.000 ;
  RECT 1072.000 0.000 1072.800 1.000 ;
  RECT 1065.600 0.000 1066.400 1.000 ;
  RECT 1051.200 0.000 1052.000 1.000 ;
  RECT 1045.600 0.000 1046.400 1.000 ;
  RECT 1031.200 0.000 1032.000 1.000 ;
  RECT 1024.800 0.000 1025.600 1.000 ;
  RECT 1010.000 0.000 1010.800 1.000 ;
  RECT 1004.800 0.000 1005.600 1.000 ;
  RECT 992.000 0.000 992.800 1.000 ;
  RECT 990.400 0.000 991.200 1.000 ;
  RECT 983.600 0.000 984.400 1.000 ;
  RECT 969.200 0.000 970.000 1.000 ;
  RECT 964.000 0.000 964.800 1.000 ;
  RECT 949.200 0.000 950.000 1.000 ;
  RECT 942.800 0.000 943.600 1.000 ;
  RECT 928.400 0.000 929.200 1.000 ;
  RECT 923.200 0.000 924.000 1.000 ;
  RECT 908.400 0.000 909.200 1.000 ;
  RECT 902.000 0.000 902.800 1.000 ;
  RECT 887.200 0.000 888.000 1.000 ;
  RECT 882.000 0.000 882.800 1.000 ;
  RECT 867.600 0.000 868.400 1.000 ;
  RECT 861.200 0.000 862.000 1.000 ;
  RECT 846.400 0.000 847.200 1.000 ;
  RECT 841.200 0.000 842.000 1.000 ;
  RECT 826.400 0.000 827.200 1.000 ;
  RECT 820.000 0.000 820.800 1.000 ;
  RECT 805.600 0.000 806.400 1.000 ;
  RECT 800.400 0.000 801.200 1.000 ;
  RECT 785.600 0.000 786.400 1.000 ;
  RECT 779.200 0.000 780.000 1.000 ;
  RECT 764.400 0.000 765.200 1.000 ;
  RECT 759.200 0.000 760.000 1.000 ;
  RECT 744.800 0.000 745.600 1.000 ;
  RECT 738.400 0.000 739.200 1.000 ;
  RECT 723.600 0.000 724.400 1.000 ;
  RECT 718.400 0.000 719.200 1.000 ;
  RECT 704.000 0.000 704.800 1.000 ;
  RECT 697.200 0.000 698.000 1.000 ;
  RECT 682.800 0.000 683.600 1.000 ;
  RECT 677.600 0.000 678.400 1.000 ;
  RECT 664.800 0.000 665.600 1.000 ;
  RECT 662.800 0.000 663.600 1.000 ;
  RECT 656.400 0.000 657.200 1.000 ;
  RECT 642.000 0.000 642.800 1.000 ;
  RECT 636.400 0.000 637.200 1.000 ;
  RECT 622.000 0.000 622.800 1.000 ;
  RECT 615.600 0.000 616.400 1.000 ;
  RECT 600.800 0.000 601.600 1.000 ;
  RECT 595.600 0.000 596.400 1.000 ;
  RECT 581.200 0.000 582.000 1.000 ;
  RECT 574.400 0.000 575.200 1.000 ;
  RECT 560.000 0.000 560.800 1.000 ;
  RECT 554.800 0.000 555.600 1.000 ;
  RECT 540.000 0.000 540.800 1.000 ;
  RECT 533.600 0.000 534.400 1.000 ;
  RECT 519.200 0.000 520.000 1.000 ;
  RECT 514.000 0.000 514.800 1.000 ;
  RECT 499.200 0.000 500.000 1.000 ;
  RECT 492.800 0.000 493.600 1.000 ;
  RECT 478.000 0.000 478.800 1.000 ;
  RECT 472.800 0.000 473.600 1.000 ;
  RECT 458.400 0.000 459.200 1.000 ;
  RECT 452.000 0.000 452.800 1.000 ;
  RECT 437.200 0.000 438.000 1.000 ;
  RECT 432.000 0.000 432.800 1.000 ;
  RECT 417.200 0.000 418.000 1.000 ;
  RECT 410.800 0.000 411.600 1.000 ;
  RECT 396.400 0.000 397.200 1.000 ;
  RECT 391.200 0.000 392.000 1.000 ;
  RECT 376.400 0.000 377.200 1.000 ;
  RECT 370.000 0.000 370.800 1.000 ;
  RECT 355.200 0.000 356.000 1.000 ;
  RECT 350.000 0.000 350.800 1.000 ;
  RECT 337.200 0.000 338.000 1.000 ;
  RECT 335.600 0.000 336.400 1.000 ;
  RECT 329.200 0.000 330.000 1.000 ;
  RECT 314.400 0.000 315.200 1.000 ;
  RECT 309.200 0.000 310.000 1.000 ;
  RECT 294.800 0.000 295.600 1.000 ;
  RECT 288.000 0.000 288.800 1.000 ;
  RECT 273.600 0.000 274.400 1.000 ;
  RECT 268.400 0.000 269.200 1.000 ;
  RECT 253.600 0.000 254.400 1.000 ;
  RECT 247.200 0.000 248.000 1.000 ;
  RECT 232.800 0.000 233.600 1.000 ;
  RECT 227.200 0.000 228.000 1.000 ;
  RECT 212.800 0.000 213.600 1.000 ;
  RECT 206.400 0.000 207.200 1.000 ;
  RECT 191.600 0.000 192.400 1.000 ;
  RECT 186.400 0.000 187.200 1.000 ;
  RECT 172.000 0.000 172.800 1.000 ;
  RECT 165.200 0.000 166.000 1.000 ;
  RECT 150.800 0.000 151.600 1.000 ;
  RECT 145.600 0.000 146.400 1.000 ;
  RECT 130.800 0.000 131.600 1.000 ;
  RECT 124.400 0.000 125.200 1.000 ;
  RECT 110.000 0.000 110.800 1.000 ;
  RECT 104.800 0.000 105.600 1.000 ;
  RECT 90.000 0.000 90.800 1.000 ;
  RECT 83.600 0.000 84.400 1.000 ;
  RECT 68.800 0.000 69.600 1.000 ;
  RECT 63.600 0.000 64.400 1.000 ;
  RECT 49.200 0.000 50.000 1.000 ;
  RECT 42.800 0.000 43.600 1.000 ;
  RECT 28.000 0.000 28.800 1.000 ;
  RECT 22.800 0.000 23.600 1.000 ;
  RECT 10.000 0.000 10.800 1.000 ;
  RECT 8.000 0.000 8.800 1.000 ;
  LAYER VI2 ;
  RECT 2683.080 3.600 2684.940 195.930 ;
  LAYER VI1 ;
  RECT 2683.080 3.460 2684.940 196.070 ;
  LAYER VI2 ;
  RECT 0.000 3.600 1.860 195.930 ;
  LAYER VI1 ;
  RECT 0.000 3.460 1.860 196.070 ;
  LAYER VI2 ;
  RECT 2.000 196.070 2682.940 197.930 ;
  LAYER VI1 ;
  RECT 1.860 196.070 2683.080 197.930 ;
  LAYER VI2 ;
  RECT 2674.600 1.600 2682.940 3.460 ;
  LAYER VI2 ;
  RECT 2660.200 1.600 2672.280 3.460 ;
  LAYER VI2 ;
  RECT 2655.000 1.600 2657.650 3.460 ;
  LAYER VI2 ;
  RECT 2640.200 1.600 2652.440 3.460 ;
  LAYER VI2 ;
  RECT 2633.800 1.600 2637.810 3.460 ;
  LAYER VI2 ;
  RECT 2619.400 1.600 2631.360 3.460 ;
  LAYER VI2 ;
  RECT 2614.200 1.600 2616.730 3.460 ;
  LAYER VI2 ;
  RECT 2599.400 1.600 2611.520 3.460 ;
  LAYER VI2 ;
  RECT 2593.000 1.600 2596.890 3.460 ;
  LAYER VI2 ;
  RECT 2578.200 1.600 2590.440 3.460 ;
  LAYER VI2 ;
  RECT 2573.000 1.600 2575.810 3.460 ;
  LAYER VI2 ;
  RECT 2558.600 1.600 2570.600 3.460 ;
  LAYER VI2 ;
  RECT 2552.200 1.600 2555.970 3.460 ;
  LAYER VI2 ;
  RECT 2537.400 1.600 2549.520 3.460 ;
  LAYER VI2 ;
  RECT 2532.200 1.600 2534.890 3.460 ;
  LAYER VI2 ;
  RECT 2517.400 1.600 2529.680 3.460 ;
  LAYER VI2 ;
  RECT 2511.000 1.600 2515.050 3.460 ;
  LAYER VI2 ;
  RECT 2496.600 1.600 2508.600 3.460 ;
  LAYER VI2 ;
  RECT 2491.400 1.600 2493.970 3.460 ;
  LAYER VI2 ;
  RECT 2476.600 1.600 2488.760 3.460 ;
  LAYER VI2 ;
  RECT 2470.200 1.600 2474.130 3.460 ;
  LAYER VI2 ;
  RECT 2455.400 1.600 2467.680 3.460 ;
  LAYER VI2 ;
  RECT 2450.200 1.600 2453.050 3.460 ;
  LAYER VI2 ;
  RECT 2435.800 1.600 2447.840 3.460 ;
  LAYER VI2 ;
  RECT 2429.400 1.600 2433.210 3.460 ;
  LAYER VI2 ;
  RECT 2414.600 1.600 2426.760 3.460 ;
  LAYER VI2 ;
  RECT 2409.400 1.600 2412.130 3.460 ;
  LAYER VI2 ;
  RECT 2394.600 1.600 2406.920 3.460 ;
  LAYER VI2 ;
  RECT 2388.200 1.600 2392.290 3.460 ;
  LAYER VI2 ;
  RECT 2373.800 1.600 2385.840 3.460 ;
  LAYER VI2 ;
  RECT 2368.600 1.600 2371.210 3.460 ;
  LAYER VI2 ;
  RECT 2355.400 1.600 2366.000 3.460 ;
  LAYER VI2 ;
  RECT 2347.400 1.600 2351.370 3.460 ;
  LAYER VI2 ;
  RECT 2332.600 1.600 2344.920 3.460 ;
  LAYER VI2 ;
  RECT 2327.400 1.600 2330.290 3.460 ;
  LAYER VI2 ;
  RECT 2313.000 1.600 2325.080 3.460 ;
  LAYER VI2 ;
  RECT 2306.600 1.600 2310.450 3.460 ;
  LAYER VI2 ;
  RECT 2291.800 1.600 2304.000 3.460 ;
  LAYER VI2 ;
  RECT 2286.600 1.600 2289.370 3.460 ;
  LAYER VI2 ;
  RECT 2272.200 1.600 2284.160 3.460 ;
  LAYER VI2 ;
  RECT 2265.400 1.600 2269.530 3.460 ;
  LAYER VI2 ;
  RECT 2251.000 1.600 2263.080 3.460 ;
  LAYER VI2 ;
  RECT 2245.800 1.600 2248.450 3.460 ;
  LAYER VI2 ;
  RECT 2231.000 1.600 2243.240 3.460 ;
  LAYER VI2 ;
  RECT 2224.600 1.600 2228.610 3.460 ;
  LAYER VI2 ;
  RECT 2210.200 1.600 2222.160 3.460 ;
  LAYER VI2 ;
  RECT 2205.000 1.600 2207.530 3.460 ;
  LAYER VI2 ;
  RECT 2190.200 1.600 2202.320 3.460 ;
  LAYER VI2 ;
  RECT 2183.800 1.600 2187.690 3.460 ;
  LAYER VI2 ;
  RECT 2169.000 1.600 2181.240 3.460 ;
  LAYER VI2 ;
  RECT 2163.800 1.600 2166.610 3.460 ;
  LAYER VI2 ;
  RECT 2149.400 1.600 2161.400 3.460 ;
  LAYER VI2 ;
  RECT 2143.000 1.600 2146.770 3.460 ;
  LAYER VI2 ;
  RECT 2128.200 1.600 2140.320 3.460 ;
  LAYER VI2 ;
  RECT 2123.000 1.600 2125.690 3.460 ;
  LAYER VI2 ;
  RECT 2108.200 1.600 2120.480 3.460 ;
  LAYER VI2 ;
  RECT 2101.800 1.600 2105.850 3.460 ;
  LAYER VI2 ;
  RECT 2087.400 1.600 2099.400 3.460 ;
  LAYER VI2 ;
  RECT 2082.200 1.600 2084.770 3.460 ;
  LAYER VI2 ;
  RECT 2067.400 1.600 2079.560 3.460 ;
  LAYER VI2 ;
  RECT 2061.000 1.600 2064.930 3.460 ;
  LAYER VI2 ;
  RECT 2046.200 1.600 2058.480 3.460 ;
  LAYER VI2 ;
  RECT 2041.000 1.600 2043.850 3.460 ;
  LAYER VI2 ;
  RECT 2028.200 1.600 2038.640 3.460 ;
  LAYER VI2 ;
  RECT 2020.200 1.600 2024.010 3.460 ;
  LAYER VI2 ;
  RECT 2005.400 1.600 2017.560 3.460 ;
  LAYER VI2 ;
  RECT 2000.200 1.600 2002.930 3.460 ;
  LAYER VI2 ;
  RECT 1985.400 1.600 1997.720 3.460 ;
  LAYER VI2 ;
  RECT 1979.000 1.600 1983.090 3.460 ;
  LAYER VI2 ;
  RECT 1964.600 1.600 1976.640 3.460 ;
  LAYER VI2 ;
  RECT 1959.400 1.600 1962.010 3.460 ;
  LAYER VI2 ;
  RECT 1944.600 1.600 1956.800 3.460 ;
  LAYER VI2 ;
  RECT 1938.200 1.600 1942.170 3.460 ;
  LAYER VI2 ;
  RECT 1923.400 1.600 1935.720 3.460 ;
  LAYER VI2 ;
  RECT 1918.200 1.600 1921.090 3.460 ;
  LAYER VI2 ;
  RECT 1903.800 1.600 1915.880 3.460 ;
  LAYER VI2 ;
  RECT 1897.400 1.600 1901.250 3.460 ;
  LAYER VI2 ;
  RECT 1882.600 1.600 1894.800 3.460 ;
  LAYER VI2 ;
  RECT 1877.400 1.600 1880.170 3.460 ;
  LAYER VI2 ;
  RECT 1863.000 1.600 1874.960 3.460 ;
  LAYER VI2 ;
  RECT 1856.200 1.600 1860.330 3.460 ;
  LAYER VI2 ;
  RECT 1841.800 1.600 1853.880 3.460 ;
  LAYER VI2 ;
  RECT 1836.600 1.600 1839.250 3.460 ;
  LAYER VI2 ;
  RECT 1821.800 1.600 1834.040 3.460 ;
  LAYER VI2 ;
  RECT 1815.400 1.600 1819.410 3.460 ;
  LAYER VI2 ;
  RECT 1801.000 1.600 1812.960 3.460 ;
  LAYER VI2 ;
  RECT 1795.800 1.600 1798.330 3.460 ;
  LAYER VI2 ;
  RECT 1781.000 1.600 1793.120 3.460 ;
  LAYER VI2 ;
  RECT 1774.600 1.600 1778.490 3.460 ;
  LAYER VI2 ;
  RECT 1759.800 1.600 1772.040 3.460 ;
  LAYER VI2 ;
  RECT 1754.600 1.600 1757.410 3.460 ;
  LAYER VI2 ;
  RECT 1740.200 1.600 1752.200 3.460 ;
  LAYER VI2 ;
  RECT 1733.800 1.600 1737.570 3.460 ;
  LAYER VI2 ;
  RECT 1719.000 1.600 1731.120 3.460 ;
  LAYER VI2 ;
  RECT 1713.800 1.600 1716.490 3.460 ;
  LAYER VI2 ;
  RECT 1701.000 1.600 1711.280 3.460 ;
  LAYER VI2 ;
  RECT 1692.600 1.600 1696.650 3.460 ;
  LAYER VI2 ;
  RECT 1678.200 1.600 1690.200 3.460 ;
  LAYER VI2 ;
  RECT 1673.000 1.600 1675.570 3.460 ;
  LAYER VI2 ;
  RECT 1658.200 1.600 1670.360 3.460 ;
  LAYER VI2 ;
  RECT 1651.800 1.600 1655.730 3.460 ;
  LAYER VI2 ;
  RECT 1637.000 1.600 1649.280 3.460 ;
  LAYER VI2 ;
  RECT 1631.800 1.600 1634.650 3.460 ;
  LAYER VI2 ;
  RECT 1617.400 1.600 1629.440 3.460 ;
  LAYER VI2 ;
  RECT 1611.000 1.600 1614.810 3.460 ;
  LAYER VI2 ;
  RECT 1596.200 1.600 1608.360 3.460 ;
  LAYER VI2 ;
  RECT 1591.000 1.600 1593.730 3.460 ;
  LAYER VI2 ;
  RECT 1576.200 1.600 1588.520 3.460 ;
  LAYER VI2 ;
  RECT 1569.800 1.600 1573.890 3.460 ;
  LAYER VI2 ;
  RECT 1555.400 1.600 1567.440 3.460 ;
  LAYER VI2 ;
  RECT 1550.200 1.600 1552.810 3.460 ;
  LAYER VI2 ;
  RECT 1535.400 1.600 1547.600 3.460 ;
  LAYER VI2 ;
  RECT 1529.000 1.600 1532.970 3.460 ;
  LAYER VI2 ;
  RECT 1514.200 1.600 1526.520 3.460 ;
  LAYER VI2 ;
  RECT 1509.000 1.600 1511.890 3.460 ;
  LAYER VI2 ;
  RECT 1494.600 1.600 1506.680 3.460 ;
  LAYER VI2 ;
  RECT 1488.200 1.600 1492.050 3.460 ;
  LAYER VI2 ;
  RECT 1473.400 1.600 1485.600 3.460 ;
  LAYER VI2 ;
  RECT 1468.200 1.600 1470.970 3.460 ;
  LAYER VI2 ;
  RECT 1453.800 1.600 1465.760 3.460 ;
  LAYER VI2 ;
  RECT 1447.000 1.600 1451.130 3.460 ;
  LAYER VI2 ;
  RECT 1432.600 1.600 1444.680 3.460 ;
  LAYER VI2 ;
  RECT 1427.400 1.600 1430.050 3.460 ;
  LAYER VI2 ;
  RECT 1412.600 1.600 1424.840 3.460 ;
  LAYER VI2 ;
  RECT 1406.200 1.600 1410.210 3.460 ;
  LAYER VI2 ;
  RECT 1391.800 1.600 1403.760 3.460 ;
  LAYER VI2 ;
  RECT 1386.600 1.600 1389.130 3.460 ;
  LAYER VI2 ;
  RECT 1373.400 1.600 1383.920 3.460 ;
  LAYER VI2 ;
  RECT 1351.000 1.600 1369.290 3.460 ;
  LAYER VI2 ;
  RECT 1339.000 1.600 1342.450 3.460 ;
  LAYER VI2 ;
  RECT 1331.800 1.600 1336.480 3.460 ;
  LAYER VI2 ;
  RECT 1313.000 1.600 1317.360 3.460 ;
  LAYER VI2 ;
  RECT 1298.200 1.600 1310.460 3.460 ;
  LAYER VI2 ;
  RECT 1293.000 1.600 1295.830 3.460 ;
  LAYER VI2 ;
  RECT 1278.600 1.600 1290.620 3.460 ;
  LAYER VI2 ;
  RECT 1272.200 1.600 1275.990 3.460 ;
  LAYER VI2 ;
  RECT 1257.400 1.600 1269.540 3.460 ;
  LAYER VI2 ;
  RECT 1252.200 1.600 1254.910 3.460 ;
  LAYER VI2 ;
  RECT 1237.400 1.600 1249.700 3.460 ;
  LAYER VI2 ;
  RECT 1231.000 1.600 1235.070 3.460 ;
  LAYER VI2 ;
  RECT 1216.600 1.600 1228.620 3.460 ;
  LAYER VI2 ;
  RECT 1211.400 1.600 1213.990 3.460 ;
  LAYER VI2 ;
  RECT 1196.600 1.600 1208.780 3.460 ;
  LAYER VI2 ;
  RECT 1190.200 1.600 1194.150 3.460 ;
  LAYER VI2 ;
  RECT 1175.400 1.600 1187.700 3.460 ;
  LAYER VI2 ;
  RECT 1170.200 1.600 1173.070 3.460 ;
  LAYER VI2 ;
  RECT 1155.800 1.600 1167.860 3.460 ;
  LAYER VI2 ;
  RECT 1149.400 1.600 1153.230 3.460 ;
  LAYER VI2 ;
  RECT 1134.600 1.600 1146.780 3.460 ;
  LAYER VI2 ;
  RECT 1129.400 1.600 1132.150 3.460 ;
  LAYER VI2 ;
  RECT 1115.000 1.600 1126.940 3.460 ;
  LAYER VI2 ;
  RECT 1108.200 1.600 1112.310 3.460 ;
  LAYER VI2 ;
  RECT 1093.800 1.600 1105.860 3.460 ;
  LAYER VI2 ;
  RECT 1088.600 1.600 1091.230 3.460 ;
  LAYER VI2 ;
  RECT 1073.800 1.600 1086.020 3.460 ;
  LAYER VI2 ;
  RECT 1067.400 1.600 1071.390 3.460 ;
  LAYER VI2 ;
  RECT 1053.000 1.600 1064.940 3.460 ;
  LAYER VI2 ;
  RECT 1047.400 1.600 1050.310 3.460 ;
  LAYER VI2 ;
  RECT 1033.000 1.600 1045.100 3.460 ;
  LAYER VI2 ;
  RECT 1026.600 1.600 1030.470 3.460 ;
  LAYER VI2 ;
  RECT 1011.800 1.600 1024.020 3.460 ;
  LAYER VI2 ;
  RECT 1006.600 1.600 1009.390 3.460 ;
  LAYER VI2 ;
  RECT 993.800 1.600 1004.180 3.460 ;
  LAYER VI2 ;
  RECT 985.400 1.600 989.550 3.460 ;
  LAYER VI2 ;
  RECT 971.000 1.600 983.100 3.460 ;
  LAYER VI2 ;
  RECT 965.800 1.600 968.470 3.460 ;
  LAYER VI2 ;
  RECT 951.000 1.600 963.260 3.460 ;
  LAYER VI2 ;
  RECT 944.600 1.600 948.630 3.460 ;
  LAYER VI2 ;
  RECT 930.200 1.600 942.180 3.460 ;
  LAYER VI2 ;
  RECT 925.000 1.600 927.550 3.460 ;
  LAYER VI2 ;
  RECT 910.200 1.600 922.340 3.460 ;
  LAYER VI2 ;
  RECT 903.800 1.600 907.710 3.460 ;
  LAYER VI2 ;
  RECT 889.000 1.600 901.260 3.460 ;
  LAYER VI2 ;
  RECT 883.800 1.600 886.630 3.460 ;
  LAYER VI2 ;
  RECT 869.400 1.600 881.420 3.460 ;
  LAYER VI2 ;
  RECT 863.000 1.600 866.790 3.460 ;
  LAYER VI2 ;
  RECT 848.200 1.600 860.340 3.460 ;
  LAYER VI2 ;
  RECT 843.000 1.600 845.710 3.460 ;
  LAYER VI2 ;
  RECT 828.200 1.600 840.500 3.460 ;
  LAYER VI2 ;
  RECT 821.800 1.600 825.870 3.460 ;
  LAYER VI2 ;
  RECT 807.400 1.600 819.420 3.460 ;
  LAYER VI2 ;
  RECT 802.200 1.600 804.790 3.460 ;
  LAYER VI2 ;
  RECT 787.400 1.600 799.580 3.460 ;
  LAYER VI2 ;
  RECT 781.000 1.600 784.950 3.460 ;
  LAYER VI2 ;
  RECT 766.200 1.600 778.500 3.460 ;
  LAYER VI2 ;
  RECT 761.000 1.600 763.870 3.460 ;
  LAYER VI2 ;
  RECT 746.600 1.600 758.660 3.460 ;
  LAYER VI2 ;
  RECT 740.200 1.600 744.030 3.460 ;
  LAYER VI2 ;
  RECT 725.400 1.600 737.580 3.460 ;
  LAYER VI2 ;
  RECT 720.200 1.600 722.950 3.460 ;
  LAYER VI2 ;
  RECT 705.800 1.600 717.740 3.460 ;
  LAYER VI2 ;
  RECT 699.000 1.600 703.110 3.460 ;
  LAYER VI2 ;
  RECT 684.600 1.600 696.660 3.460 ;
  LAYER VI2 ;
  RECT 679.400 1.600 682.030 3.460 ;
  LAYER VI2 ;
  RECT 666.600 1.600 676.820 3.460 ;
  LAYER VI2 ;
  RECT 658.200 1.600 662.190 3.460 ;
  LAYER VI2 ;
  RECT 643.800 1.600 655.740 3.460 ;
  LAYER VI2 ;
  RECT 638.200 1.600 641.110 3.460 ;
  LAYER VI2 ;
  RECT 623.800 1.600 635.900 3.460 ;
  LAYER VI2 ;
  RECT 617.400 1.600 621.270 3.460 ;
  LAYER VI2 ;
  RECT 602.600 1.600 614.820 3.460 ;
  LAYER VI2 ;
  RECT 597.400 1.600 600.190 3.460 ;
  LAYER VI2 ;
  RECT 583.000 1.600 594.980 3.460 ;
  LAYER VI2 ;
  RECT 576.200 1.600 580.350 3.460 ;
  LAYER VI2 ;
  RECT 561.800 1.600 573.900 3.460 ;
  LAYER VI2 ;
  RECT 556.600 1.600 559.270 3.460 ;
  LAYER VI2 ;
  RECT 541.800 1.600 554.060 3.460 ;
  LAYER VI2 ;
  RECT 535.400 1.600 539.430 3.460 ;
  LAYER VI2 ;
  RECT 521.000 1.600 532.980 3.460 ;
  LAYER VI2 ;
  RECT 515.800 1.600 518.350 3.460 ;
  LAYER VI2 ;
  RECT 501.000 1.600 513.140 3.460 ;
  LAYER VI2 ;
  RECT 494.600 1.600 498.510 3.460 ;
  LAYER VI2 ;
  RECT 479.800 1.600 492.060 3.460 ;
  LAYER VI2 ;
  RECT 474.600 1.600 477.430 3.460 ;
  LAYER VI2 ;
  RECT 460.200 1.600 472.220 3.460 ;
  LAYER VI2 ;
  RECT 453.800 1.600 457.590 3.460 ;
  LAYER VI2 ;
  RECT 439.000 1.600 451.140 3.460 ;
  LAYER VI2 ;
  RECT 433.800 1.600 436.510 3.460 ;
  LAYER VI2 ;
  RECT 419.000 1.600 431.300 3.460 ;
  LAYER VI2 ;
  RECT 412.600 1.600 416.670 3.460 ;
  LAYER VI2 ;
  RECT 398.200 1.600 410.220 3.460 ;
  LAYER VI2 ;
  RECT 393.000 1.600 395.590 3.460 ;
  LAYER VI2 ;
  RECT 378.200 1.600 390.380 3.460 ;
  LAYER VI2 ;
  RECT 371.800 1.600 375.750 3.460 ;
  LAYER VI2 ;
  RECT 357.000 1.600 369.300 3.460 ;
  LAYER VI2 ;
  RECT 351.800 1.600 354.670 3.460 ;
  LAYER VI2 ;
  RECT 339.000 1.600 349.460 3.460 ;
  LAYER VI2 ;
  RECT 331.000 1.600 334.830 3.460 ;
  LAYER VI2 ;
  RECT 316.200 1.600 328.380 3.460 ;
  LAYER VI2 ;
  RECT 311.000 1.600 313.750 3.460 ;
  LAYER VI2 ;
  RECT 296.600 1.600 308.540 3.460 ;
  LAYER VI2 ;
  RECT 289.800 1.600 293.910 3.460 ;
  LAYER VI2 ;
  RECT 275.400 1.600 287.460 3.460 ;
  LAYER VI2 ;
  RECT 270.200 1.600 272.830 3.460 ;
  LAYER VI2 ;
  RECT 255.400 1.600 267.620 3.460 ;
  LAYER VI2 ;
  RECT 249.000 1.600 252.990 3.460 ;
  LAYER VI2 ;
  RECT 234.600 1.600 246.540 3.460 ;
  LAYER VI2 ;
  RECT 229.000 1.600 231.910 3.460 ;
  LAYER VI2 ;
  RECT 214.600 1.600 226.700 3.460 ;
  LAYER VI2 ;
  RECT 208.200 1.600 212.070 3.460 ;
  LAYER VI2 ;
  RECT 193.400 1.600 205.620 3.460 ;
  LAYER VI2 ;
  RECT 188.200 1.600 190.990 3.460 ;
  LAYER VI2 ;
  RECT 173.800 1.600 185.780 3.460 ;
  LAYER VI2 ;
  RECT 167.000 1.600 171.150 3.460 ;
  LAYER VI2 ;
  RECT 152.600 1.600 164.700 3.460 ;
  LAYER VI2 ;
  RECT 147.400 1.600 150.070 3.460 ;
  LAYER VI2 ;
  RECT 132.600 1.600 144.860 3.460 ;
  LAYER VI2 ;
  RECT 126.200 1.600 130.230 3.460 ;
  LAYER VI2 ;
  RECT 111.800 1.600 123.780 3.460 ;
  LAYER VI2 ;
  RECT 106.600 1.600 109.150 3.460 ;
  LAYER VI2 ;
  RECT 91.800 1.600 103.940 3.460 ;
  LAYER VI2 ;
  RECT 85.400 1.600 89.310 3.460 ;
  LAYER VI2 ;
  RECT 70.600 1.600 82.860 3.460 ;
  LAYER VI2 ;
  RECT 65.400 1.600 68.230 3.460 ;
  LAYER VI2 ;
  RECT 51.000 1.600 63.020 3.460 ;
  LAYER VI2 ;
  RECT 44.600 1.600 48.390 3.460 ;
  LAYER VI2 ;
  RECT 29.800 1.600 41.940 3.460 ;
  LAYER VI2 ;
  RECT 24.600 1.600 27.310 3.460 ;
  LAYER VI2 ;
  RECT 11.800 1.600 22.100 3.460 ;
  LAYER VI2 ;
  RECT 2.000 1.600 7.470 3.460 ;
  LAYER VI1 ;
  RECT 2674.600 1.600 2683.080 3.460 ;
  LAYER VI1 ;
  RECT 2660.200 1.600 2672.280 3.460 ;
  LAYER VI1 ;
  RECT 2655.000 1.600 2657.650 3.460 ;
  LAYER VI1 ;
  RECT 2640.200 1.600 2652.440 3.460 ;
  LAYER VI1 ;
  RECT 2633.800 1.600 2637.810 3.460 ;
  LAYER VI1 ;
  RECT 2619.400 1.600 2631.360 3.460 ;
  LAYER VI1 ;
  RECT 2614.200 1.600 2616.730 3.460 ;
  LAYER VI1 ;
  RECT 2599.400 1.600 2611.520 3.460 ;
  LAYER VI1 ;
  RECT 2593.000 1.600 2596.890 3.460 ;
  LAYER VI1 ;
  RECT 2578.200 1.600 2590.440 3.460 ;
  LAYER VI1 ;
  RECT 2573.000 1.600 2575.810 3.460 ;
  LAYER VI1 ;
  RECT 2558.600 1.600 2570.600 3.460 ;
  LAYER VI1 ;
  RECT 2552.200 1.600 2555.970 3.460 ;
  LAYER VI1 ;
  RECT 2537.400 1.600 2549.520 3.460 ;
  LAYER VI1 ;
  RECT 2532.200 1.600 2534.890 3.460 ;
  LAYER VI1 ;
  RECT 2517.400 1.600 2529.680 3.460 ;
  LAYER VI1 ;
  RECT 2511.000 1.600 2515.050 3.460 ;
  LAYER VI1 ;
  RECT 2496.600 1.600 2508.600 3.460 ;
  LAYER VI1 ;
  RECT 2491.400 1.600 2493.970 3.460 ;
  LAYER VI1 ;
  RECT 2476.600 1.600 2488.760 3.460 ;
  LAYER VI1 ;
  RECT 2470.200 1.600 2474.130 3.460 ;
  LAYER VI1 ;
  RECT 2455.400 1.600 2467.680 3.460 ;
  LAYER VI1 ;
  RECT 2450.200 1.600 2453.050 3.460 ;
  LAYER VI1 ;
  RECT 2435.800 1.600 2447.840 3.460 ;
  LAYER VI1 ;
  RECT 2429.400 1.600 2433.210 3.460 ;
  LAYER VI1 ;
  RECT 2414.600 1.600 2426.760 3.460 ;
  LAYER VI1 ;
  RECT 2409.400 1.600 2412.130 3.460 ;
  LAYER VI1 ;
  RECT 2394.600 1.600 2406.920 3.460 ;
  LAYER VI1 ;
  RECT 2388.200 1.600 2392.290 3.460 ;
  LAYER VI1 ;
  RECT 2373.800 1.600 2385.840 3.460 ;
  LAYER VI1 ;
  RECT 2368.600 1.600 2371.210 3.460 ;
  LAYER VI1 ;
  RECT 2355.400 1.600 2366.000 3.460 ;
  LAYER VI1 ;
  RECT 2347.400 1.600 2351.370 3.460 ;
  LAYER VI1 ;
  RECT 2332.600 1.600 2344.920 3.460 ;
  LAYER VI1 ;
  RECT 2327.400 1.600 2330.290 3.460 ;
  LAYER VI1 ;
  RECT 2313.000 1.600 2325.080 3.460 ;
  LAYER VI1 ;
  RECT 2306.600 1.600 2310.450 3.460 ;
  LAYER VI1 ;
  RECT 2291.800 1.600 2304.000 3.460 ;
  LAYER VI1 ;
  RECT 2286.600 1.600 2289.370 3.460 ;
  LAYER VI1 ;
  RECT 2272.200 1.600 2284.160 3.460 ;
  LAYER VI1 ;
  RECT 2265.400 1.600 2269.530 3.460 ;
  LAYER VI1 ;
  RECT 2251.000 1.600 2263.080 3.460 ;
  LAYER VI1 ;
  RECT 2245.800 1.600 2248.450 3.460 ;
  LAYER VI1 ;
  RECT 2231.000 1.600 2243.240 3.460 ;
  LAYER VI1 ;
  RECT 2224.600 1.600 2228.610 3.460 ;
  LAYER VI1 ;
  RECT 2210.200 1.600 2222.160 3.460 ;
  LAYER VI1 ;
  RECT 2205.000 1.600 2207.530 3.460 ;
  LAYER VI1 ;
  RECT 2190.200 1.600 2202.320 3.460 ;
  LAYER VI1 ;
  RECT 2183.800 1.600 2187.690 3.460 ;
  LAYER VI1 ;
  RECT 2169.000 1.600 2181.240 3.460 ;
  LAYER VI1 ;
  RECT 2163.800 1.600 2166.610 3.460 ;
  LAYER VI1 ;
  RECT 2149.400 1.600 2161.400 3.460 ;
  LAYER VI1 ;
  RECT 2143.000 1.600 2146.770 3.460 ;
  LAYER VI1 ;
  RECT 2128.200 1.600 2140.320 3.460 ;
  LAYER VI1 ;
  RECT 2123.000 1.600 2125.690 3.460 ;
  LAYER VI1 ;
  RECT 2108.200 1.600 2120.480 3.460 ;
  LAYER VI1 ;
  RECT 2101.800 1.600 2105.850 3.460 ;
  LAYER VI1 ;
  RECT 2087.400 1.600 2099.400 3.460 ;
  LAYER VI1 ;
  RECT 2082.200 1.600 2084.770 3.460 ;
  LAYER VI1 ;
  RECT 2067.400 1.600 2079.560 3.460 ;
  LAYER VI1 ;
  RECT 2061.000 1.600 2064.930 3.460 ;
  LAYER VI1 ;
  RECT 2046.200 1.600 2058.480 3.460 ;
  LAYER VI1 ;
  RECT 2041.000 1.600 2043.850 3.460 ;
  LAYER VI1 ;
  RECT 2028.200 1.600 2038.640 3.460 ;
  LAYER VI1 ;
  RECT 2020.200 1.600 2024.010 3.460 ;
  LAYER VI1 ;
  RECT 2005.400 1.600 2017.560 3.460 ;
  LAYER VI1 ;
  RECT 2000.200 1.600 2002.930 3.460 ;
  LAYER VI1 ;
  RECT 1985.400 1.600 1997.720 3.460 ;
  LAYER VI1 ;
  RECT 1979.000 1.600 1983.090 3.460 ;
  LAYER VI1 ;
  RECT 1964.600 1.600 1976.640 3.460 ;
  LAYER VI1 ;
  RECT 1959.400 1.600 1962.010 3.460 ;
  LAYER VI1 ;
  RECT 1944.600 1.600 1956.800 3.460 ;
  LAYER VI1 ;
  RECT 1938.200 1.600 1942.170 3.460 ;
  LAYER VI1 ;
  RECT 1923.400 1.600 1935.720 3.460 ;
  LAYER VI1 ;
  RECT 1918.200 1.600 1921.090 3.460 ;
  LAYER VI1 ;
  RECT 1903.800 1.600 1915.880 3.460 ;
  LAYER VI1 ;
  RECT 1897.400 1.600 1901.250 3.460 ;
  LAYER VI1 ;
  RECT 1882.600 1.600 1894.800 3.460 ;
  LAYER VI1 ;
  RECT 1877.400 1.600 1880.170 3.460 ;
  LAYER VI1 ;
  RECT 1863.000 1.600 1874.960 3.460 ;
  LAYER VI1 ;
  RECT 1856.200 1.600 1860.330 3.460 ;
  LAYER VI1 ;
  RECT 1841.800 1.600 1853.880 3.460 ;
  LAYER VI1 ;
  RECT 1836.600 1.600 1839.250 3.460 ;
  LAYER VI1 ;
  RECT 1821.800 1.600 1834.040 3.460 ;
  LAYER VI1 ;
  RECT 1815.400 1.600 1819.410 3.460 ;
  LAYER VI1 ;
  RECT 1801.000 1.600 1812.960 3.460 ;
  LAYER VI1 ;
  RECT 1795.800 1.600 1798.330 3.460 ;
  LAYER VI1 ;
  RECT 1781.000 1.600 1793.120 3.460 ;
  LAYER VI1 ;
  RECT 1774.600 1.600 1778.490 3.460 ;
  LAYER VI1 ;
  RECT 1759.800 1.600 1772.040 3.460 ;
  LAYER VI1 ;
  RECT 1754.600 1.600 1757.410 3.460 ;
  LAYER VI1 ;
  RECT 1740.200 1.600 1752.200 3.460 ;
  LAYER VI1 ;
  RECT 1733.800 1.600 1737.570 3.460 ;
  LAYER VI1 ;
  RECT 1719.000 1.600 1731.120 3.460 ;
  LAYER VI1 ;
  RECT 1713.800 1.600 1716.490 3.460 ;
  LAYER VI1 ;
  RECT 1701.000 1.600 1711.280 3.460 ;
  LAYER VI1 ;
  RECT 1692.600 1.600 1696.650 3.460 ;
  LAYER VI1 ;
  RECT 1678.200 1.600 1690.200 3.460 ;
  LAYER VI1 ;
  RECT 1673.000 1.600 1675.570 3.460 ;
  LAYER VI1 ;
  RECT 1658.200 1.600 1670.360 3.460 ;
  LAYER VI1 ;
  RECT 1651.800 1.600 1655.730 3.460 ;
  LAYER VI1 ;
  RECT 1637.000 1.600 1649.280 3.460 ;
  LAYER VI1 ;
  RECT 1631.800 1.600 1634.650 3.460 ;
  LAYER VI1 ;
  RECT 1617.400 1.600 1629.440 3.460 ;
  LAYER VI1 ;
  RECT 1611.000 1.600 1614.810 3.460 ;
  LAYER VI1 ;
  RECT 1596.200 1.600 1608.360 3.460 ;
  LAYER VI1 ;
  RECT 1591.000 1.600 1593.730 3.460 ;
  LAYER VI1 ;
  RECT 1576.200 1.600 1588.520 3.460 ;
  LAYER VI1 ;
  RECT 1569.800 1.600 1573.890 3.460 ;
  LAYER VI1 ;
  RECT 1555.400 1.600 1567.440 3.460 ;
  LAYER VI1 ;
  RECT 1550.200 1.600 1552.810 3.460 ;
  LAYER VI1 ;
  RECT 1535.400 1.600 1547.600 3.460 ;
  LAYER VI1 ;
  RECT 1529.000 1.600 1532.970 3.460 ;
  LAYER VI1 ;
  RECT 1514.200 1.600 1526.520 3.460 ;
  LAYER VI1 ;
  RECT 1509.000 1.600 1511.890 3.460 ;
  LAYER VI1 ;
  RECT 1494.600 1.600 1506.680 3.460 ;
  LAYER VI1 ;
  RECT 1488.200 1.600 1492.050 3.460 ;
  LAYER VI1 ;
  RECT 1473.400 1.600 1485.600 3.460 ;
  LAYER VI1 ;
  RECT 1468.200 1.600 1470.970 3.460 ;
  LAYER VI1 ;
  RECT 1453.800 1.600 1465.760 3.460 ;
  LAYER VI1 ;
  RECT 1447.000 1.600 1451.130 3.460 ;
  LAYER VI1 ;
  RECT 1432.600 1.600 1444.680 3.460 ;
  LAYER VI1 ;
  RECT 1427.400 1.600 1430.050 3.460 ;
  LAYER VI1 ;
  RECT 1412.600 1.600 1424.840 3.460 ;
  LAYER VI1 ;
  RECT 1406.200 1.600 1410.210 3.460 ;
  LAYER VI1 ;
  RECT 1391.800 1.600 1403.760 3.460 ;
  LAYER VI1 ;
  RECT 1386.600 1.600 1389.130 3.460 ;
  LAYER VI1 ;
  RECT 1373.400 1.600 1383.920 3.460 ;
  LAYER VI1 ;
  RECT 1351.000 1.600 1369.290 3.460 ;
  LAYER VI1 ;
  RECT 1339.000 1.600 1342.450 3.460 ;
  LAYER VI1 ;
  RECT 1331.800 1.600 1336.480 3.460 ;
  LAYER VI1 ;
  RECT 1313.000 1.600 1317.360 3.460 ;
  LAYER VI1 ;
  RECT 1298.200 1.600 1310.460 3.460 ;
  LAYER VI1 ;
  RECT 1293.000 1.600 1295.830 3.460 ;
  LAYER VI1 ;
  RECT 1278.600 1.600 1290.620 3.460 ;
  LAYER VI1 ;
  RECT 1272.200 1.600 1275.990 3.460 ;
  LAYER VI1 ;
  RECT 1257.400 1.600 1269.540 3.460 ;
  LAYER VI1 ;
  RECT 1252.200 1.600 1254.910 3.460 ;
  LAYER VI1 ;
  RECT 1237.400 1.600 1249.700 3.460 ;
  LAYER VI1 ;
  RECT 1231.000 1.600 1235.070 3.460 ;
  LAYER VI1 ;
  RECT 1216.600 1.600 1228.620 3.460 ;
  LAYER VI1 ;
  RECT 1211.400 1.600 1213.990 3.460 ;
  LAYER VI1 ;
  RECT 1196.600 1.600 1208.780 3.460 ;
  LAYER VI1 ;
  RECT 1190.200 1.600 1194.150 3.460 ;
  LAYER VI1 ;
  RECT 1175.400 1.600 1187.700 3.460 ;
  LAYER VI1 ;
  RECT 1170.200 1.600 1173.070 3.460 ;
  LAYER VI1 ;
  RECT 1155.800 1.600 1167.860 3.460 ;
  LAYER VI1 ;
  RECT 1149.400 1.600 1153.230 3.460 ;
  LAYER VI1 ;
  RECT 1134.600 1.600 1146.780 3.460 ;
  LAYER VI1 ;
  RECT 1129.400 1.600 1132.150 3.460 ;
  LAYER VI1 ;
  RECT 1115.000 1.600 1126.940 3.460 ;
  LAYER VI1 ;
  RECT 1108.200 1.600 1112.310 3.460 ;
  LAYER VI1 ;
  RECT 1093.800 1.600 1105.860 3.460 ;
  LAYER VI1 ;
  RECT 1088.600 1.600 1091.230 3.460 ;
  LAYER VI1 ;
  RECT 1073.800 1.600 1086.020 3.460 ;
  LAYER VI1 ;
  RECT 1067.400 1.600 1071.390 3.460 ;
  LAYER VI1 ;
  RECT 1053.000 1.600 1064.940 3.460 ;
  LAYER VI1 ;
  RECT 1047.400 1.600 1050.310 3.460 ;
  LAYER VI1 ;
  RECT 1033.000 1.600 1045.100 3.460 ;
  LAYER VI1 ;
  RECT 1026.600 1.600 1030.470 3.460 ;
  LAYER VI1 ;
  RECT 1011.800 1.600 1024.020 3.460 ;
  LAYER VI1 ;
  RECT 1006.600 1.600 1009.390 3.460 ;
  LAYER VI1 ;
  RECT 993.800 1.600 1004.180 3.460 ;
  LAYER VI1 ;
  RECT 985.400 1.600 989.550 3.460 ;
  LAYER VI1 ;
  RECT 971.000 1.600 983.100 3.460 ;
  LAYER VI1 ;
  RECT 965.800 1.600 968.470 3.460 ;
  LAYER VI1 ;
  RECT 951.000 1.600 963.260 3.460 ;
  LAYER VI1 ;
  RECT 944.600 1.600 948.630 3.460 ;
  LAYER VI1 ;
  RECT 930.200 1.600 942.180 3.460 ;
  LAYER VI1 ;
  RECT 925.000 1.600 927.550 3.460 ;
  LAYER VI1 ;
  RECT 910.200 1.600 922.340 3.460 ;
  LAYER VI1 ;
  RECT 903.800 1.600 907.710 3.460 ;
  LAYER VI1 ;
  RECT 889.000 1.600 901.260 3.460 ;
  LAYER VI1 ;
  RECT 883.800 1.600 886.630 3.460 ;
  LAYER VI1 ;
  RECT 869.400 1.600 881.420 3.460 ;
  LAYER VI1 ;
  RECT 863.000 1.600 866.790 3.460 ;
  LAYER VI1 ;
  RECT 848.200 1.600 860.340 3.460 ;
  LAYER VI1 ;
  RECT 843.000 1.600 845.710 3.460 ;
  LAYER VI1 ;
  RECT 828.200 1.600 840.500 3.460 ;
  LAYER VI1 ;
  RECT 821.800 1.600 825.870 3.460 ;
  LAYER VI1 ;
  RECT 807.400 1.600 819.420 3.460 ;
  LAYER VI1 ;
  RECT 802.200 1.600 804.790 3.460 ;
  LAYER VI1 ;
  RECT 787.400 1.600 799.580 3.460 ;
  LAYER VI1 ;
  RECT 781.000 1.600 784.950 3.460 ;
  LAYER VI1 ;
  RECT 766.200 1.600 778.500 3.460 ;
  LAYER VI1 ;
  RECT 761.000 1.600 763.870 3.460 ;
  LAYER VI1 ;
  RECT 746.600 1.600 758.660 3.460 ;
  LAYER VI1 ;
  RECT 740.200 1.600 744.030 3.460 ;
  LAYER VI1 ;
  RECT 725.400 1.600 737.580 3.460 ;
  LAYER VI1 ;
  RECT 720.200 1.600 722.950 3.460 ;
  LAYER VI1 ;
  RECT 705.800 1.600 717.740 3.460 ;
  LAYER VI1 ;
  RECT 699.000 1.600 703.110 3.460 ;
  LAYER VI1 ;
  RECT 684.600 1.600 696.660 3.460 ;
  LAYER VI1 ;
  RECT 679.400 1.600 682.030 3.460 ;
  LAYER VI1 ;
  RECT 666.600 1.600 676.820 3.460 ;
  LAYER VI1 ;
  RECT 658.200 1.600 662.190 3.460 ;
  LAYER VI1 ;
  RECT 643.800 1.600 655.740 3.460 ;
  LAYER VI1 ;
  RECT 638.200 1.600 641.110 3.460 ;
  LAYER VI1 ;
  RECT 623.800 1.600 635.900 3.460 ;
  LAYER VI1 ;
  RECT 617.400 1.600 621.270 3.460 ;
  LAYER VI1 ;
  RECT 602.600 1.600 614.820 3.460 ;
  LAYER VI1 ;
  RECT 597.400 1.600 600.190 3.460 ;
  LAYER VI1 ;
  RECT 583.000 1.600 594.980 3.460 ;
  LAYER VI1 ;
  RECT 576.200 1.600 580.350 3.460 ;
  LAYER VI1 ;
  RECT 561.800 1.600 573.900 3.460 ;
  LAYER VI1 ;
  RECT 556.600 1.600 559.270 3.460 ;
  LAYER VI1 ;
  RECT 541.800 1.600 554.060 3.460 ;
  LAYER VI1 ;
  RECT 535.400 1.600 539.430 3.460 ;
  LAYER VI1 ;
  RECT 521.000 1.600 532.980 3.460 ;
  LAYER VI1 ;
  RECT 515.800 1.600 518.350 3.460 ;
  LAYER VI1 ;
  RECT 501.000 1.600 513.140 3.460 ;
  LAYER VI1 ;
  RECT 494.600 1.600 498.510 3.460 ;
  LAYER VI1 ;
  RECT 479.800 1.600 492.060 3.460 ;
  LAYER VI1 ;
  RECT 474.600 1.600 477.430 3.460 ;
  LAYER VI1 ;
  RECT 460.200 1.600 472.220 3.460 ;
  LAYER VI1 ;
  RECT 453.800 1.600 457.590 3.460 ;
  LAYER VI1 ;
  RECT 439.000 1.600 451.140 3.460 ;
  LAYER VI1 ;
  RECT 433.800 1.600 436.510 3.460 ;
  LAYER VI1 ;
  RECT 419.000 1.600 431.300 3.460 ;
  LAYER VI1 ;
  RECT 412.600 1.600 416.670 3.460 ;
  LAYER VI1 ;
  RECT 398.200 1.600 410.220 3.460 ;
  LAYER VI1 ;
  RECT 393.000 1.600 395.590 3.460 ;
  LAYER VI1 ;
  RECT 378.200 1.600 390.380 3.460 ;
  LAYER VI1 ;
  RECT 371.800 1.600 375.750 3.460 ;
  LAYER VI1 ;
  RECT 357.000 1.600 369.300 3.460 ;
  LAYER VI1 ;
  RECT 351.800 1.600 354.670 3.460 ;
  LAYER VI1 ;
  RECT 339.000 1.600 349.460 3.460 ;
  LAYER VI1 ;
  RECT 331.000 1.600 334.830 3.460 ;
  LAYER VI1 ;
  RECT 316.200 1.600 328.380 3.460 ;
  LAYER VI1 ;
  RECT 311.000 1.600 313.750 3.460 ;
  LAYER VI1 ;
  RECT 296.600 1.600 308.540 3.460 ;
  LAYER VI1 ;
  RECT 289.800 1.600 293.910 3.460 ;
  LAYER VI1 ;
  RECT 275.400 1.600 287.460 3.460 ;
  LAYER VI1 ;
  RECT 270.200 1.600 272.830 3.460 ;
  LAYER VI1 ;
  RECT 255.400 1.600 267.620 3.460 ;
  LAYER VI1 ;
  RECT 249.000 1.600 252.990 3.460 ;
  LAYER VI1 ;
  RECT 234.600 1.600 246.540 3.460 ;
  LAYER VI1 ;
  RECT 229.000 1.600 231.910 3.460 ;
  LAYER VI1 ;
  RECT 214.600 1.600 226.700 3.460 ;
  LAYER VI1 ;
  RECT 208.200 1.600 212.070 3.460 ;
  LAYER VI1 ;
  RECT 193.400 1.600 205.620 3.460 ;
  LAYER VI1 ;
  RECT 188.200 1.600 190.990 3.460 ;
  LAYER VI1 ;
  RECT 173.800 1.600 185.780 3.460 ;
  LAYER VI1 ;
  RECT 167.000 1.600 171.150 3.460 ;
  LAYER VI1 ;
  RECT 152.600 1.600 164.700 3.460 ;
  LAYER VI1 ;
  RECT 147.400 1.600 150.070 3.460 ;
  LAYER VI1 ;
  RECT 132.600 1.600 144.860 3.460 ;
  LAYER VI1 ;
  RECT 126.200 1.600 130.230 3.460 ;
  LAYER VI1 ;
  RECT 111.800 1.600 123.780 3.460 ;
  LAYER VI1 ;
  RECT 106.600 1.600 109.150 3.460 ;
  LAYER VI1 ;
  RECT 91.800 1.600 103.940 3.460 ;
  LAYER VI1 ;
  RECT 85.400 1.600 89.310 3.460 ;
  LAYER VI1 ;
  RECT 70.600 1.600 82.860 3.460 ;
  LAYER VI1 ;
  RECT 65.400 1.600 68.230 3.460 ;
  LAYER VI1 ;
  RECT 51.000 1.600 63.020 3.460 ;
  LAYER VI1 ;
  RECT 44.600 1.600 48.390 3.460 ;
  LAYER VI1 ;
  RECT 29.800 1.600 41.940 3.460 ;
  LAYER VI1 ;
  RECT 24.600 1.600 27.310 3.460 ;
  LAYER VI1 ;
  RECT 11.800 1.600 22.100 3.460 ;
  LAYER VI1 ;
  RECT 1.860 1.600 7.470 3.460 ;
  LAYER VI3 ;
  RECT 2680.940 187.000 2682.660 193.930 ;
  LAYER VI3 ;
  RECT 2680.940 64.930 2682.660 67.240 ;
  LAYER VI3 ;
  RECT 2680.940 44.080 2682.660 61.260 ;
  LAYER VI3 ;
  RECT 2680.940 39.620 2682.660 41.480 ;
  LAYER VI3 ;
  RECT 2680.940 29.870 2682.660 33.520 ;
  LAYER VI3 ;
  RECT 2680.940 24.270 2682.660 26.870 ;
  LAYER VI3 ;
  RECT 2680.940 18.130 2682.660 21.270 ;
  LAYER VI3 ;
  RECT 2680.940 5.600 2682.660 11.230 ;
  LAYER VI2 ;
  RECT 2680.940 187.000 2682.660 193.930 ;
  LAYER VI2 ;
  RECT 2680.940 64.930 2682.660 67.240 ;
  LAYER VI2 ;
  RECT 2680.940 44.080 2682.660 61.260 ;
  LAYER VI2 ;
  RECT 2680.940 39.620 2682.660 41.480 ;
  LAYER VI2 ;
  RECT 2680.940 29.870 2682.660 33.520 ;
  LAYER VI2 ;
  RECT 2680.940 24.270 2682.660 26.870 ;
  LAYER VI2 ;
  RECT 2680.940 18.130 2682.660 21.270 ;
  LAYER VI2 ;
  RECT 2680.940 5.600 2682.660 11.230 ;
  LAYER VI1 ;
  RECT 2680.940 5.600 2682.800 193.930 ;
  LAYER VI3 ;
  RECT 2.280 187.000 4.000 193.930 ;
  LAYER VI3 ;
  RECT 2.280 64.930 4.000 67.240 ;
  LAYER VI3 ;
  RECT 2.280 44.080 4.000 61.260 ;
  LAYER VI3 ;
  RECT 2.280 39.620 4.000 41.480 ;
  LAYER VI3 ;
  RECT 2.280 29.870 4.000 33.520 ;
  LAYER VI3 ;
  RECT 2.280 24.270 4.000 26.870 ;
  LAYER VI3 ;
  RECT 2.280 18.130 4.000 21.270 ;
  LAYER VI3 ;
  RECT 2.280 5.600 4.000 11.230 ;
  LAYER VI2 ;
  RECT 2.280 187.000 4.000 193.930 ;
  LAYER VI2 ;
  RECT 2.280 64.930 4.000 67.240 ;
  LAYER VI2 ;
  RECT 2.280 44.080 4.000 61.260 ;
  LAYER VI2 ;
  RECT 2.280 39.620 4.000 41.480 ;
  LAYER VI2 ;
  RECT 2.280 29.870 4.000 33.520 ;
  LAYER VI2 ;
  RECT 2.280 24.270 4.000 26.870 ;
  LAYER VI2 ;
  RECT 2.280 18.130 4.000 21.270 ;
  LAYER VI2 ;
  RECT 2.280 5.600 4.000 11.230 ;
  LAYER VI1 ;
  RECT 2.140 5.600 4.000 193.930 ;
  LAYER VI3 ;
  RECT 2638.020 193.930 2680.940 195.650 ;
  LAYER VI3 ;
  RECT 2597.100 193.930 2635.770 195.650 ;
  LAYER VI3 ;
  RECT 2556.180 193.930 2594.850 195.650 ;
  LAYER VI3 ;
  RECT 2515.260 193.930 2553.930 195.650 ;
  LAYER VI3 ;
  RECT 2474.340 193.930 2513.010 195.650 ;
  LAYER VI3 ;
  RECT 2433.420 193.930 2472.090 195.650 ;
  LAYER VI3 ;
  RECT 2392.500 193.930 2431.170 195.650 ;
  LAYER VI3 ;
  RECT 2351.580 193.930 2390.250 195.650 ;
  LAYER VI3 ;
  RECT 2310.660 193.930 2349.330 195.650 ;
  LAYER VI3 ;
  RECT 2269.740 193.930 2308.410 195.650 ;
  LAYER VI3 ;
  RECT 2228.820 193.930 2267.490 195.650 ;
  LAYER VI3 ;
  RECT 2187.900 193.930 2226.570 195.650 ;
  LAYER VI3 ;
  RECT 2146.980 193.930 2185.650 195.650 ;
  LAYER VI3 ;
  RECT 2106.060 193.930 2144.730 195.650 ;
  LAYER VI3 ;
  RECT 2065.140 193.930 2103.810 195.650 ;
  LAYER VI3 ;
  RECT 2024.220 193.930 2062.890 195.650 ;
  LAYER VI3 ;
  RECT 1983.300 193.930 2021.970 195.650 ;
  LAYER VI3 ;
  RECT 1942.380 193.930 1981.050 195.650 ;
  LAYER VI3 ;
  RECT 1901.460 193.930 1940.130 195.650 ;
  LAYER VI3 ;
  RECT 1860.540 193.930 1899.210 195.650 ;
  LAYER VI3 ;
  RECT 1819.620 193.930 1858.290 195.650 ;
  LAYER VI3 ;
  RECT 1778.700 193.930 1817.370 195.650 ;
  LAYER VI3 ;
  RECT 1737.780 193.930 1776.450 195.650 ;
  LAYER VI3 ;
  RECT 1696.860 193.930 1735.530 195.650 ;
  LAYER VI3 ;
  RECT 1655.940 193.930 1694.610 195.650 ;
  LAYER VI3 ;
  RECT 1615.020 193.930 1653.690 195.650 ;
  LAYER VI3 ;
  RECT 1574.100 193.930 1612.770 195.650 ;
  LAYER VI3 ;
  RECT 1533.180 193.930 1571.850 195.650 ;
  LAYER VI3 ;
  RECT 1492.260 193.930 1530.930 195.650 ;
  LAYER VI3 ;
  RECT 1451.340 193.930 1490.010 195.650 ;
  LAYER VI3 ;
  RECT 1410.420 193.930 1449.090 195.650 ;
  LAYER VI3 ;
  RECT 1369.500 193.930 1408.170 195.650 ;
  LAYER VI3 ;
  RECT 1350.760 193.930 1363.760 195.650 ;
  LAYER VI3 ;
  RECT 1339.630 193.930 1344.440 195.650 ;
  LAYER VI3 ;
  RECT 1329.920 193.930 1334.440 195.650 ;
  LAYER VI3 ;
  RECT 1324.580 193.930 1326.160 195.650 ;
  LAYER VI3 ;
  RECT 1276.770 193.930 1315.800 195.650 ;
  LAYER VI3 ;
  RECT 1235.850 193.930 1274.520 195.650 ;
  LAYER VI3 ;
  RECT 1194.930 193.930 1233.600 195.650 ;
  LAYER VI3 ;
  RECT 1154.010 193.930 1192.680 195.650 ;
  LAYER VI3 ;
  RECT 1113.090 193.930 1151.760 195.650 ;
  LAYER VI3 ;
  RECT 1072.170 193.930 1110.840 195.650 ;
  LAYER VI3 ;
  RECT 1031.250 193.930 1069.920 195.650 ;
  LAYER VI3 ;
  RECT 990.330 193.930 1029.000 195.650 ;
  LAYER VI3 ;
  RECT 949.410 193.930 988.080 195.650 ;
  LAYER VI3 ;
  RECT 908.490 193.930 947.160 195.650 ;
  LAYER VI3 ;
  RECT 867.570 193.930 906.240 195.650 ;
  LAYER VI3 ;
  RECT 826.650 193.930 865.320 195.650 ;
  LAYER VI3 ;
  RECT 785.730 193.930 824.400 195.650 ;
  LAYER VI3 ;
  RECT 744.810 193.930 783.480 195.650 ;
  LAYER VI3 ;
  RECT 703.890 193.930 742.560 195.650 ;
  LAYER VI3 ;
  RECT 662.970 193.930 701.640 195.650 ;
  LAYER VI3 ;
  RECT 622.050 193.930 660.720 195.650 ;
  LAYER VI3 ;
  RECT 581.130 193.930 619.800 195.650 ;
  LAYER VI3 ;
  RECT 540.210 193.930 578.880 195.650 ;
  LAYER VI3 ;
  RECT 499.290 193.930 537.960 195.650 ;
  LAYER VI3 ;
  RECT 458.370 193.930 497.040 195.650 ;
  LAYER VI3 ;
  RECT 417.450 193.930 456.120 195.650 ;
  LAYER VI3 ;
  RECT 376.530 193.930 415.200 195.650 ;
  LAYER VI3 ;
  RECT 335.610 193.930 374.280 195.650 ;
  LAYER VI3 ;
  RECT 294.690 193.930 333.360 195.650 ;
  LAYER VI3 ;
  RECT 253.770 193.930 292.440 195.650 ;
  LAYER VI3 ;
  RECT 212.850 193.930 251.520 195.650 ;
  LAYER VI3 ;
  RECT 171.930 193.930 210.600 195.650 ;
  LAYER VI3 ;
  RECT 131.010 193.930 169.680 195.650 ;
  LAYER VI3 ;
  RECT 90.090 193.930 128.760 195.650 ;
  LAYER VI3 ;
  RECT 49.170 193.930 87.840 195.650 ;
  LAYER VI3 ;
  RECT 4.000 193.930 46.920 195.650 ;
  LAYER VI2 ;
  RECT 2638.020 193.930 2680.940 195.650 ;
  LAYER VI2 ;
  RECT 2597.100 193.930 2635.770 195.650 ;
  LAYER VI2 ;
  RECT 2556.180 193.930 2594.850 195.650 ;
  LAYER VI2 ;
  RECT 2515.260 193.930 2553.930 195.650 ;
  LAYER VI2 ;
  RECT 2474.340 193.930 2513.010 195.650 ;
  LAYER VI2 ;
  RECT 2433.420 193.930 2472.090 195.650 ;
  LAYER VI2 ;
  RECT 2392.500 193.930 2431.170 195.650 ;
  LAYER VI2 ;
  RECT 2351.580 193.930 2390.250 195.650 ;
  LAYER VI2 ;
  RECT 2310.660 193.930 2349.330 195.650 ;
  LAYER VI2 ;
  RECT 2269.740 193.930 2308.410 195.650 ;
  LAYER VI2 ;
  RECT 2228.820 193.930 2267.490 195.650 ;
  LAYER VI2 ;
  RECT 2187.900 193.930 2226.570 195.650 ;
  LAYER VI2 ;
  RECT 2146.980 193.930 2185.650 195.650 ;
  LAYER VI2 ;
  RECT 2106.060 193.930 2144.730 195.650 ;
  LAYER VI2 ;
  RECT 2065.140 193.930 2103.810 195.650 ;
  LAYER VI2 ;
  RECT 2024.220 193.930 2062.890 195.650 ;
  LAYER VI2 ;
  RECT 1983.300 193.930 2021.970 195.650 ;
  LAYER VI2 ;
  RECT 1942.380 193.930 1981.050 195.650 ;
  LAYER VI2 ;
  RECT 1901.460 193.930 1940.130 195.650 ;
  LAYER VI2 ;
  RECT 1860.540 193.930 1899.210 195.650 ;
  LAYER VI2 ;
  RECT 1819.620 193.930 1858.290 195.650 ;
  LAYER VI2 ;
  RECT 1778.700 193.930 1817.370 195.650 ;
  LAYER VI2 ;
  RECT 1737.780 193.930 1776.450 195.650 ;
  LAYER VI2 ;
  RECT 1696.860 193.930 1735.530 195.650 ;
  LAYER VI2 ;
  RECT 1655.940 193.930 1694.610 195.650 ;
  LAYER VI2 ;
  RECT 1615.020 193.930 1653.690 195.650 ;
  LAYER VI2 ;
  RECT 1574.100 193.930 1612.770 195.650 ;
  LAYER VI2 ;
  RECT 1533.180 193.930 1571.850 195.650 ;
  LAYER VI2 ;
  RECT 1492.260 193.930 1530.930 195.650 ;
  LAYER VI2 ;
  RECT 1451.340 193.930 1490.010 195.650 ;
  LAYER VI2 ;
  RECT 1410.420 193.930 1449.090 195.650 ;
  LAYER VI2 ;
  RECT 1369.500 193.930 1408.170 195.650 ;
  LAYER VI2 ;
  RECT 1350.760 193.930 1363.760 195.650 ;
  LAYER VI2 ;
  RECT 1339.630 193.930 1344.440 195.650 ;
  LAYER VI2 ;
  RECT 1329.920 193.930 1334.440 195.650 ;
  LAYER VI2 ;
  RECT 1324.580 193.930 1326.160 195.650 ;
  LAYER VI2 ;
  RECT 1276.770 193.930 1315.800 195.650 ;
  LAYER VI2 ;
  RECT 1235.850 193.930 1274.520 195.650 ;
  LAYER VI2 ;
  RECT 1194.930 193.930 1233.600 195.650 ;
  LAYER VI2 ;
  RECT 1154.010 193.930 1192.680 195.650 ;
  LAYER VI2 ;
  RECT 1113.090 193.930 1151.760 195.650 ;
  LAYER VI2 ;
  RECT 1072.170 193.930 1110.840 195.650 ;
  LAYER VI2 ;
  RECT 1031.250 193.930 1069.920 195.650 ;
  LAYER VI2 ;
  RECT 990.330 193.930 1029.000 195.650 ;
  LAYER VI2 ;
  RECT 949.410 193.930 988.080 195.650 ;
  LAYER VI2 ;
  RECT 908.490 193.930 947.160 195.650 ;
  LAYER VI2 ;
  RECT 867.570 193.930 906.240 195.650 ;
  LAYER VI2 ;
  RECT 826.650 193.930 865.320 195.650 ;
  LAYER VI2 ;
  RECT 785.730 193.930 824.400 195.650 ;
  LAYER VI2 ;
  RECT 744.810 193.930 783.480 195.650 ;
  LAYER VI2 ;
  RECT 703.890 193.930 742.560 195.650 ;
  LAYER VI2 ;
  RECT 662.970 193.930 701.640 195.650 ;
  LAYER VI2 ;
  RECT 622.050 193.930 660.720 195.650 ;
  LAYER VI2 ;
  RECT 581.130 193.930 619.800 195.650 ;
  LAYER VI2 ;
  RECT 540.210 193.930 578.880 195.650 ;
  LAYER VI2 ;
  RECT 499.290 193.930 537.960 195.650 ;
  LAYER VI2 ;
  RECT 458.370 193.930 497.040 195.650 ;
  LAYER VI2 ;
  RECT 417.450 193.930 456.120 195.650 ;
  LAYER VI2 ;
  RECT 376.530 193.930 415.200 195.650 ;
  LAYER VI2 ;
  RECT 335.610 193.930 374.280 195.650 ;
  LAYER VI2 ;
  RECT 294.690 193.930 333.360 195.650 ;
  LAYER VI2 ;
  RECT 253.770 193.930 292.440 195.650 ;
  LAYER VI2 ;
  RECT 212.850 193.930 251.520 195.650 ;
  LAYER VI2 ;
  RECT 171.930 193.930 210.600 195.650 ;
  LAYER VI2 ;
  RECT 131.010 193.930 169.680 195.650 ;
  LAYER VI2 ;
  RECT 90.090 193.930 128.760 195.650 ;
  LAYER VI2 ;
  RECT 49.170 193.930 87.840 195.650 ;
  LAYER VI2 ;
  RECT 4.000 193.930 46.920 195.650 ;
  LAYER VI1 ;
  RECT 4.000 193.930 2680.940 195.790 ;
  LAYER VI3 ;
  RECT 2667.540 3.880 2677.380 5.600 ;
  LAYER VI3 ;
  RECT 2647.700 3.880 2657.540 5.600 ;
  LAYER VI3 ;
  RECT 2626.620 3.880 2637.700 5.600 ;
  LAYER VI3 ;
  RECT 2606.780 3.880 2616.620 5.600 ;
  LAYER VI3 ;
  RECT 2585.700 3.880 2596.780 5.600 ;
  LAYER VI3 ;
  RECT 2565.860 3.880 2575.700 5.600 ;
  LAYER VI3 ;
  RECT 2544.780 3.880 2555.860 5.600 ;
  LAYER VI3 ;
  RECT 2524.940 3.880 2534.780 5.600 ;
  LAYER VI3 ;
  RECT 2503.860 3.880 2514.940 5.600 ;
  LAYER VI3 ;
  RECT 2484.020 3.880 2493.860 5.600 ;
  LAYER VI3 ;
  RECT 2462.940 3.880 2474.020 5.600 ;
  LAYER VI3 ;
  RECT 2443.100 3.880 2452.940 5.600 ;
  LAYER VI3 ;
  RECT 2422.020 3.880 2433.100 5.600 ;
  LAYER VI3 ;
  RECT 2402.180 3.880 2412.020 5.600 ;
  LAYER VI3 ;
  RECT 2381.100 3.880 2392.180 5.600 ;
  LAYER VI3 ;
  RECT 2361.260 3.880 2371.100 5.600 ;
  LAYER VI3 ;
  RECT 2340.180 3.880 2351.260 5.600 ;
  LAYER VI3 ;
  RECT 2320.340 3.880 2330.180 5.600 ;
  LAYER VI3 ;
  RECT 2299.260 3.880 2310.340 5.600 ;
  LAYER VI3 ;
  RECT 2279.420 3.880 2289.260 5.600 ;
  LAYER VI3 ;
  RECT 2258.340 3.880 2269.420 5.600 ;
  LAYER VI3 ;
  RECT 2238.500 3.880 2248.340 5.600 ;
  LAYER VI3 ;
  RECT 2217.420 3.880 2228.500 5.600 ;
  LAYER VI3 ;
  RECT 2197.580 3.880 2207.420 5.600 ;
  LAYER VI3 ;
  RECT 2176.500 3.880 2187.580 5.600 ;
  LAYER VI3 ;
  RECT 2156.660 3.880 2166.500 5.600 ;
  LAYER VI3 ;
  RECT 2135.580 3.880 2146.660 5.600 ;
  LAYER VI3 ;
  RECT 2115.740 3.880 2125.580 5.600 ;
  LAYER VI3 ;
  RECT 2094.660 3.880 2105.740 5.600 ;
  LAYER VI3 ;
  RECT 2074.820 3.880 2084.660 5.600 ;
  LAYER VI3 ;
  RECT 2053.740 3.880 2064.820 5.600 ;
  LAYER VI3 ;
  RECT 2033.900 3.880 2043.740 5.600 ;
  LAYER VI3 ;
  RECT 2012.820 3.880 2023.900 5.600 ;
  LAYER VI3 ;
  RECT 1992.980 3.880 2002.820 5.600 ;
  LAYER VI3 ;
  RECT 1971.900 3.880 1982.980 5.600 ;
  LAYER VI3 ;
  RECT 1952.060 3.880 1961.900 5.600 ;
  LAYER VI3 ;
  RECT 1930.980 3.880 1942.060 5.600 ;
  LAYER VI3 ;
  RECT 1911.140 3.880 1920.980 5.600 ;
  LAYER VI3 ;
  RECT 1890.060 3.880 1901.140 5.600 ;
  LAYER VI3 ;
  RECT 1870.220 3.880 1880.060 5.600 ;
  LAYER VI3 ;
  RECT 1849.140 3.880 1860.220 5.600 ;
  LAYER VI3 ;
  RECT 1829.300 3.880 1839.140 5.600 ;
  LAYER VI3 ;
  RECT 1808.220 3.880 1819.300 5.600 ;
  LAYER VI3 ;
  RECT 1788.380 3.880 1798.220 5.600 ;
  LAYER VI3 ;
  RECT 1767.300 3.880 1778.380 5.600 ;
  LAYER VI3 ;
  RECT 1747.460 3.880 1757.300 5.600 ;
  LAYER VI3 ;
  RECT 1726.380 3.880 1737.460 5.600 ;
  LAYER VI3 ;
  RECT 1706.540 3.880 1716.380 5.600 ;
  LAYER VI3 ;
  RECT 1685.460 3.880 1696.540 5.600 ;
  LAYER VI3 ;
  RECT 1665.620 3.880 1675.460 5.600 ;
  LAYER VI3 ;
  RECT 1644.540 3.880 1655.620 5.600 ;
  LAYER VI3 ;
  RECT 1624.700 3.880 1634.540 5.600 ;
  LAYER VI3 ;
  RECT 1603.620 3.880 1614.700 5.600 ;
  LAYER VI3 ;
  RECT 1583.780 3.880 1593.620 5.600 ;
  LAYER VI3 ;
  RECT 1562.700 3.880 1573.780 5.600 ;
  LAYER VI3 ;
  RECT 1542.860 3.880 1552.700 5.600 ;
  LAYER VI3 ;
  RECT 1521.780 3.880 1532.860 5.600 ;
  LAYER VI3 ;
  RECT 1501.940 3.880 1511.780 5.600 ;
  LAYER VI3 ;
  RECT 1480.860 3.880 1491.940 5.600 ;
  LAYER VI3 ;
  RECT 1461.020 3.880 1470.860 5.600 ;
  LAYER VI3 ;
  RECT 1439.940 3.880 1451.020 5.600 ;
  LAYER VI3 ;
  RECT 1420.100 3.880 1429.940 5.600 ;
  LAYER VI3 ;
  RECT 1399.020 3.880 1410.100 5.600 ;
  LAYER VI3 ;
  RECT 1379.180 3.880 1389.020 5.600 ;
  LAYER VI3 ;
  RECT 1351.210 3.880 1369.180 5.600 ;
  LAYER VI3 ;
  RECT 1339.890 3.880 1343.290 5.600 ;
  LAYER VI3 ;
  RECT 1329.920 3.880 1334.440 5.600 ;
  LAYER VI3 ;
  RECT 1324.580 3.880 1326.160 5.600 ;
  LAYER VI3 ;
  RECT 1305.720 3.880 1316.820 5.600 ;
  LAYER VI3 ;
  RECT 1285.880 3.880 1295.720 5.600 ;
  LAYER VI3 ;
  RECT 1264.800 3.880 1275.880 5.600 ;
  LAYER VI3 ;
  RECT 1244.960 3.880 1254.800 5.600 ;
  LAYER VI3 ;
  RECT 1223.880 3.880 1234.960 5.600 ;
  LAYER VI3 ;
  RECT 1204.040 3.880 1213.880 5.600 ;
  LAYER VI3 ;
  RECT 1182.960 3.880 1194.040 5.600 ;
  LAYER VI3 ;
  RECT 1163.120 3.880 1172.960 5.600 ;
  LAYER VI3 ;
  RECT 1142.040 3.880 1153.120 5.600 ;
  LAYER VI3 ;
  RECT 1122.200 3.880 1132.040 5.600 ;
  LAYER VI3 ;
  RECT 1101.120 3.880 1112.200 5.600 ;
  LAYER VI3 ;
  RECT 1081.280 3.880 1091.120 5.600 ;
  LAYER VI3 ;
  RECT 1060.200 3.880 1071.280 5.600 ;
  LAYER VI3 ;
  RECT 1040.360 3.880 1050.200 5.600 ;
  LAYER VI3 ;
  RECT 1019.280 3.880 1030.360 5.600 ;
  LAYER VI3 ;
  RECT 999.440 3.880 1009.280 5.600 ;
  LAYER VI3 ;
  RECT 978.360 3.880 989.440 5.600 ;
  LAYER VI3 ;
  RECT 958.520 3.880 968.360 5.600 ;
  LAYER VI3 ;
  RECT 937.440 3.880 948.520 5.600 ;
  LAYER VI3 ;
  RECT 917.600 3.880 927.440 5.600 ;
  LAYER VI3 ;
  RECT 896.520 3.880 907.600 5.600 ;
  LAYER VI3 ;
  RECT 876.680 3.880 886.520 5.600 ;
  LAYER VI3 ;
  RECT 855.600 3.880 866.680 5.600 ;
  LAYER VI3 ;
  RECT 835.760 3.880 845.600 5.600 ;
  LAYER VI3 ;
  RECT 814.680 3.880 825.760 5.600 ;
  LAYER VI3 ;
  RECT 794.840 3.880 804.680 5.600 ;
  LAYER VI3 ;
  RECT 773.760 3.880 784.840 5.600 ;
  LAYER VI3 ;
  RECT 753.920 3.880 763.760 5.600 ;
  LAYER VI3 ;
  RECT 732.840 3.880 743.920 5.600 ;
  LAYER VI3 ;
  RECT 713.000 3.880 722.840 5.600 ;
  LAYER VI3 ;
  RECT 691.920 3.880 703.000 5.600 ;
  LAYER VI3 ;
  RECT 672.080 3.880 681.920 5.600 ;
  LAYER VI3 ;
  RECT 651.000 3.880 662.080 5.600 ;
  LAYER VI3 ;
  RECT 631.160 3.880 641.000 5.600 ;
  LAYER VI3 ;
  RECT 610.080 3.880 621.160 5.600 ;
  LAYER VI3 ;
  RECT 590.240 3.880 600.080 5.600 ;
  LAYER VI3 ;
  RECT 569.160 3.880 580.240 5.600 ;
  LAYER VI3 ;
  RECT 549.320 3.880 559.160 5.600 ;
  LAYER VI3 ;
  RECT 528.240 3.880 539.320 5.600 ;
  LAYER VI3 ;
  RECT 508.400 3.880 518.240 5.600 ;
  LAYER VI3 ;
  RECT 487.320 3.880 498.400 5.600 ;
  LAYER VI3 ;
  RECT 467.480 3.880 477.320 5.600 ;
  LAYER VI3 ;
  RECT 446.400 3.880 457.480 5.600 ;
  LAYER VI3 ;
  RECT 426.560 3.880 436.400 5.600 ;
  LAYER VI3 ;
  RECT 405.480 3.880 416.560 5.600 ;
  LAYER VI3 ;
  RECT 385.640 3.880 395.480 5.600 ;
  LAYER VI3 ;
  RECT 364.560 3.880 375.640 5.600 ;
  LAYER VI3 ;
  RECT 344.720 3.880 354.560 5.600 ;
  LAYER VI3 ;
  RECT 323.640 3.880 334.720 5.600 ;
  LAYER VI3 ;
  RECT 303.800 3.880 313.640 5.600 ;
  LAYER VI3 ;
  RECT 282.720 3.880 293.800 5.600 ;
  LAYER VI3 ;
  RECT 262.880 3.880 272.720 5.600 ;
  LAYER VI3 ;
  RECT 241.800 3.880 252.880 5.600 ;
  LAYER VI3 ;
  RECT 221.960 3.880 231.800 5.600 ;
  LAYER VI3 ;
  RECT 200.880 3.880 211.960 5.600 ;
  LAYER VI3 ;
  RECT 181.040 3.880 190.880 5.600 ;
  LAYER VI3 ;
  RECT 159.960 3.880 171.040 5.600 ;
  LAYER VI3 ;
  RECT 140.120 3.880 149.960 5.600 ;
  LAYER VI3 ;
  RECT 119.040 3.880 130.120 5.600 ;
  LAYER VI3 ;
  RECT 99.200 3.880 109.040 5.600 ;
  LAYER VI3 ;
  RECT 78.120 3.880 89.200 5.600 ;
  LAYER VI3 ;
  RECT 58.280 3.880 68.120 5.600 ;
  LAYER VI3 ;
  RECT 37.200 3.880 48.280 5.600 ;
  LAYER VI3 ;
  RECT 17.360 3.880 27.200 5.600 ;
  LAYER VI2 ;
  RECT 2674.600 3.880 2677.380 5.600 ;
  LAYER VI2 ;
  RECT 2667.540 3.880 2672.280 5.600 ;
  LAYER VI2 ;
  RECT 2655.000 3.880 2657.540 5.600 ;
  LAYER VI2 ;
  RECT 2647.700 3.880 2652.440 5.600 ;
  LAYER VI2 ;
  RECT 2633.800 3.880 2637.700 5.600 ;
  LAYER VI2 ;
  RECT 2626.620 3.880 2631.360 5.600 ;
  LAYER VI2 ;
  RECT 2614.200 3.880 2616.620 5.600 ;
  LAYER VI2 ;
  RECT 2606.780 3.880 2611.520 5.600 ;
  LAYER VI2 ;
  RECT 2593.000 3.880 2596.780 5.600 ;
  LAYER VI2 ;
  RECT 2585.700 3.880 2590.440 5.600 ;
  LAYER VI2 ;
  RECT 2573.000 3.880 2575.700 5.600 ;
  LAYER VI2 ;
  RECT 2565.860 3.880 2570.600 5.600 ;
  LAYER VI2 ;
  RECT 2552.200 3.880 2555.860 5.600 ;
  LAYER VI2 ;
  RECT 2544.780 3.880 2549.520 5.600 ;
  LAYER VI2 ;
  RECT 2532.200 3.880 2534.780 5.600 ;
  LAYER VI2 ;
  RECT 2524.940 3.880 2529.680 5.600 ;
  LAYER VI2 ;
  RECT 2511.000 3.880 2514.940 5.600 ;
  LAYER VI2 ;
  RECT 2503.860 3.880 2508.600 5.600 ;
  LAYER VI2 ;
  RECT 2491.400 3.880 2493.860 5.600 ;
  LAYER VI2 ;
  RECT 2484.020 3.880 2488.760 5.600 ;
  LAYER VI2 ;
  RECT 2470.200 3.880 2474.020 5.600 ;
  LAYER VI2 ;
  RECT 2462.940 3.880 2467.680 5.600 ;
  LAYER VI2 ;
  RECT 2450.200 3.880 2452.940 5.600 ;
  LAYER VI2 ;
  RECT 2443.100 3.880 2447.840 5.600 ;
  LAYER VI2 ;
  RECT 2429.400 3.880 2433.100 5.600 ;
  LAYER VI2 ;
  RECT 2422.020 3.880 2426.760 5.600 ;
  LAYER VI2 ;
  RECT 2409.400 3.880 2412.020 5.600 ;
  LAYER VI2 ;
  RECT 2402.180 3.880 2406.920 5.600 ;
  LAYER VI2 ;
  RECT 2388.200 3.880 2392.180 5.600 ;
  LAYER VI2 ;
  RECT 2381.100 3.880 2385.840 5.600 ;
  LAYER VI2 ;
  RECT 2368.600 3.880 2371.100 5.600 ;
  LAYER VI2 ;
  RECT 2361.260 3.880 2366.000 5.600 ;
  LAYER VI2 ;
  RECT 2347.400 3.880 2351.260 5.600 ;
  LAYER VI2 ;
  RECT 2340.180 3.880 2344.920 5.600 ;
  LAYER VI2 ;
  RECT 2327.400 3.880 2330.180 5.600 ;
  LAYER VI2 ;
  RECT 2320.340 3.880 2325.080 5.600 ;
  LAYER VI2 ;
  RECT 2306.600 3.880 2310.340 5.600 ;
  LAYER VI2 ;
  RECT 2299.260 3.880 2304.000 5.600 ;
  LAYER VI2 ;
  RECT 2286.600 3.880 2289.260 5.600 ;
  LAYER VI2 ;
  RECT 2279.420 3.880 2284.160 5.600 ;
  LAYER VI2 ;
  RECT 2265.400 3.880 2269.420 5.600 ;
  LAYER VI2 ;
  RECT 2258.340 3.880 2263.080 5.600 ;
  LAYER VI2 ;
  RECT 2245.800 3.880 2248.340 5.600 ;
  LAYER VI2 ;
  RECT 2238.500 3.880 2243.240 5.600 ;
  LAYER VI2 ;
  RECT 2224.600 3.880 2228.500 5.600 ;
  LAYER VI2 ;
  RECT 2217.420 3.880 2222.160 5.600 ;
  LAYER VI2 ;
  RECT 2205.000 3.880 2207.420 5.600 ;
  LAYER VI2 ;
  RECT 2197.580 3.880 2202.320 5.600 ;
  LAYER VI2 ;
  RECT 2183.800 3.880 2187.580 5.600 ;
  LAYER VI2 ;
  RECT 2176.500 3.880 2181.240 5.600 ;
  LAYER VI2 ;
  RECT 2163.800 3.880 2166.500 5.600 ;
  LAYER VI2 ;
  RECT 2156.660 3.880 2161.400 5.600 ;
  LAYER VI2 ;
  RECT 2143.000 3.880 2146.660 5.600 ;
  LAYER VI2 ;
  RECT 2135.580 3.880 2140.320 5.600 ;
  LAYER VI2 ;
  RECT 2123.000 3.880 2125.580 5.600 ;
  LAYER VI2 ;
  RECT 2115.740 3.880 2120.480 5.600 ;
  LAYER VI2 ;
  RECT 2101.800 3.880 2105.740 5.600 ;
  LAYER VI2 ;
  RECT 2094.660 3.880 2099.400 5.600 ;
  LAYER VI2 ;
  RECT 2082.200 3.880 2084.660 5.600 ;
  LAYER VI2 ;
  RECT 2074.820 3.880 2079.560 5.600 ;
  LAYER VI2 ;
  RECT 2061.000 3.880 2064.820 5.600 ;
  LAYER VI2 ;
  RECT 2053.740 3.880 2058.480 5.600 ;
  LAYER VI2 ;
  RECT 2041.000 3.880 2043.740 5.600 ;
  LAYER VI2 ;
  RECT 2033.900 3.880 2038.640 5.600 ;
  LAYER VI2 ;
  RECT 2020.200 3.880 2023.900 5.600 ;
  LAYER VI2 ;
  RECT 2012.820 3.880 2017.560 5.600 ;
  LAYER VI2 ;
  RECT 2000.200 3.880 2002.820 5.600 ;
  LAYER VI2 ;
  RECT 1992.980 3.880 1997.720 5.600 ;
  LAYER VI2 ;
  RECT 1979.000 3.880 1982.980 5.600 ;
  LAYER VI2 ;
  RECT 1971.900 3.880 1976.640 5.600 ;
  LAYER VI2 ;
  RECT 1959.400 3.880 1961.900 5.600 ;
  LAYER VI2 ;
  RECT 1952.060 3.880 1956.800 5.600 ;
  LAYER VI2 ;
  RECT 1938.200 3.880 1942.060 5.600 ;
  LAYER VI2 ;
  RECT 1930.980 3.880 1935.720 5.600 ;
  LAYER VI2 ;
  RECT 1918.200 3.880 1920.980 5.600 ;
  LAYER VI2 ;
  RECT 1911.140 3.880 1915.880 5.600 ;
  LAYER VI2 ;
  RECT 1897.400 3.880 1901.140 5.600 ;
  LAYER VI2 ;
  RECT 1890.060 3.880 1894.800 5.600 ;
  LAYER VI2 ;
  RECT 1877.400 3.880 1880.060 5.600 ;
  LAYER VI2 ;
  RECT 1870.220 3.880 1874.960 5.600 ;
  LAYER VI2 ;
  RECT 1856.200 3.880 1860.220 5.600 ;
  LAYER VI2 ;
  RECT 1849.140 3.880 1853.880 5.600 ;
  LAYER VI2 ;
  RECT 1836.600 3.880 1839.140 5.600 ;
  LAYER VI2 ;
  RECT 1829.300 3.880 1834.040 5.600 ;
  LAYER VI2 ;
  RECT 1815.400 3.880 1819.300 5.600 ;
  LAYER VI2 ;
  RECT 1808.220 3.880 1812.960 5.600 ;
  LAYER VI2 ;
  RECT 1795.800 3.880 1798.220 5.600 ;
  LAYER VI2 ;
  RECT 1788.380 3.880 1793.120 5.600 ;
  LAYER VI2 ;
  RECT 1774.600 3.880 1778.380 5.600 ;
  LAYER VI2 ;
  RECT 1767.300 3.880 1772.040 5.600 ;
  LAYER VI2 ;
  RECT 1754.600 3.880 1757.300 5.600 ;
  LAYER VI2 ;
  RECT 1747.460 3.880 1752.200 5.600 ;
  LAYER VI2 ;
  RECT 1733.800 3.880 1737.460 5.600 ;
  LAYER VI2 ;
  RECT 1726.380 3.880 1731.120 5.600 ;
  LAYER VI2 ;
  RECT 1713.800 3.880 1716.380 5.600 ;
  LAYER VI2 ;
  RECT 1706.540 3.880 1711.280 5.600 ;
  LAYER VI2 ;
  RECT 1692.600 3.880 1696.540 5.600 ;
  LAYER VI2 ;
  RECT 1685.460 3.880 1690.200 5.600 ;
  LAYER VI2 ;
  RECT 1673.000 3.880 1675.460 5.600 ;
  LAYER VI2 ;
  RECT 1665.620 3.880 1670.360 5.600 ;
  LAYER VI2 ;
  RECT 1651.800 3.880 1655.620 5.600 ;
  LAYER VI2 ;
  RECT 1644.540 3.880 1649.280 5.600 ;
  LAYER VI2 ;
  RECT 1631.800 3.880 1634.540 5.600 ;
  LAYER VI2 ;
  RECT 1624.700 3.880 1629.440 5.600 ;
  LAYER VI2 ;
  RECT 1611.000 3.880 1614.700 5.600 ;
  LAYER VI2 ;
  RECT 1603.620 3.880 1608.360 5.600 ;
  LAYER VI2 ;
  RECT 1591.000 3.880 1593.620 5.600 ;
  LAYER VI2 ;
  RECT 1583.780 3.880 1588.520 5.600 ;
  LAYER VI2 ;
  RECT 1569.800 3.880 1573.780 5.600 ;
  LAYER VI2 ;
  RECT 1562.700 3.880 1567.440 5.600 ;
  LAYER VI2 ;
  RECT 1550.200 3.880 1552.700 5.600 ;
  LAYER VI2 ;
  RECT 1542.860 3.880 1547.600 5.600 ;
  LAYER VI2 ;
  RECT 1529.000 3.880 1532.860 5.600 ;
  LAYER VI2 ;
  RECT 1521.780 3.880 1526.520 5.600 ;
  LAYER VI2 ;
  RECT 1509.000 3.880 1511.780 5.600 ;
  LAYER VI2 ;
  RECT 1501.940 3.880 1506.680 5.600 ;
  LAYER VI2 ;
  RECT 1488.200 3.880 1491.940 5.600 ;
  LAYER VI2 ;
  RECT 1480.860 3.880 1485.600 5.600 ;
  LAYER VI2 ;
  RECT 1468.200 3.880 1470.860 5.600 ;
  LAYER VI2 ;
  RECT 1461.020 3.880 1465.760 5.600 ;
  LAYER VI2 ;
  RECT 1447.000 3.880 1451.020 5.600 ;
  LAYER VI2 ;
  RECT 1439.940 3.880 1444.680 5.600 ;
  LAYER VI2 ;
  RECT 1427.400 3.880 1429.940 5.600 ;
  LAYER VI2 ;
  RECT 1420.100 3.880 1424.840 5.600 ;
  LAYER VI2 ;
  RECT 1406.200 3.880 1410.100 5.600 ;
  LAYER VI2 ;
  RECT 1399.020 3.880 1403.760 5.600 ;
  LAYER VI2 ;
  RECT 1386.600 3.880 1389.020 5.600 ;
  LAYER VI2 ;
  RECT 1379.180 3.880 1383.920 5.600 ;
  LAYER VI2 ;
  RECT 1351.210 3.880 1369.180 5.600 ;
  LAYER VI2 ;
  RECT 1339.890 3.880 1342.450 5.600 ;
  LAYER VI2 ;
  RECT 1331.800 3.880 1334.440 5.600 ;
  LAYER VI2 ;
  RECT 1313.000 3.880 1316.820 5.600 ;
  LAYER VI2 ;
  RECT 1305.720 3.880 1310.460 5.600 ;
  LAYER VI2 ;
  RECT 1293.000 3.880 1295.720 5.600 ;
  LAYER VI2 ;
  RECT 1285.880 3.880 1290.620 5.600 ;
  LAYER VI2 ;
  RECT 1272.200 3.880 1275.880 5.600 ;
  LAYER VI2 ;
  RECT 1264.800 3.880 1269.540 5.600 ;
  LAYER VI2 ;
  RECT 1252.200 3.880 1254.800 5.600 ;
  LAYER VI2 ;
  RECT 1244.960 3.880 1249.700 5.600 ;
  LAYER VI2 ;
  RECT 1231.000 3.880 1234.960 5.600 ;
  LAYER VI2 ;
  RECT 1223.880 3.880 1228.620 5.600 ;
  LAYER VI2 ;
  RECT 1211.400 3.880 1213.880 5.600 ;
  LAYER VI2 ;
  RECT 1204.040 3.880 1208.780 5.600 ;
  LAYER VI2 ;
  RECT 1190.200 3.880 1194.040 5.600 ;
  LAYER VI2 ;
  RECT 1182.960 3.880 1187.700 5.600 ;
  LAYER VI2 ;
  RECT 1170.200 3.880 1172.960 5.600 ;
  LAYER VI2 ;
  RECT 1163.120 3.880 1167.860 5.600 ;
  LAYER VI2 ;
  RECT 1149.400 3.880 1153.120 5.600 ;
  LAYER VI2 ;
  RECT 1142.040 3.880 1146.780 5.600 ;
  LAYER VI2 ;
  RECT 1129.400 3.880 1132.040 5.600 ;
  LAYER VI2 ;
  RECT 1122.200 3.880 1126.940 5.600 ;
  LAYER VI2 ;
  RECT 1108.200 3.880 1112.200 5.600 ;
  LAYER VI2 ;
  RECT 1101.120 3.880 1105.860 5.600 ;
  LAYER VI2 ;
  RECT 1088.600 3.880 1091.120 5.600 ;
  LAYER VI2 ;
  RECT 1081.280 3.880 1086.020 5.600 ;
  LAYER VI2 ;
  RECT 1067.400 3.880 1071.280 5.600 ;
  LAYER VI2 ;
  RECT 1060.200 3.880 1064.940 5.600 ;
  LAYER VI2 ;
  RECT 1047.400 3.880 1050.200 5.600 ;
  LAYER VI2 ;
  RECT 1040.360 3.880 1045.100 5.600 ;
  LAYER VI2 ;
  RECT 1026.600 3.880 1030.360 5.600 ;
  LAYER VI2 ;
  RECT 1019.280 3.880 1024.020 5.600 ;
  LAYER VI2 ;
  RECT 1006.600 3.880 1009.280 5.600 ;
  LAYER VI2 ;
  RECT 999.440 3.880 1004.180 5.600 ;
  LAYER VI2 ;
  RECT 985.400 3.880 989.440 5.600 ;
  LAYER VI2 ;
  RECT 978.360 3.880 983.100 5.600 ;
  LAYER VI2 ;
  RECT 965.800 3.880 968.360 5.600 ;
  LAYER VI2 ;
  RECT 958.520 3.880 963.260 5.600 ;
  LAYER VI2 ;
  RECT 944.600 3.880 948.520 5.600 ;
  LAYER VI2 ;
  RECT 937.440 3.880 942.180 5.600 ;
  LAYER VI2 ;
  RECT 925.000 3.880 927.440 5.600 ;
  LAYER VI2 ;
  RECT 917.600 3.880 922.340 5.600 ;
  LAYER VI2 ;
  RECT 903.800 3.880 907.600 5.600 ;
  LAYER VI2 ;
  RECT 896.520 3.880 901.260 5.600 ;
  LAYER VI2 ;
  RECT 883.800 3.880 886.520 5.600 ;
  LAYER VI2 ;
  RECT 876.680 3.880 881.420 5.600 ;
  LAYER VI2 ;
  RECT 863.000 3.880 866.680 5.600 ;
  LAYER VI2 ;
  RECT 855.600 3.880 860.340 5.600 ;
  LAYER VI2 ;
  RECT 843.000 3.880 845.600 5.600 ;
  LAYER VI2 ;
  RECT 835.760 3.880 840.500 5.600 ;
  LAYER VI2 ;
  RECT 821.800 3.880 825.760 5.600 ;
  LAYER VI2 ;
  RECT 814.680 3.880 819.420 5.600 ;
  LAYER VI2 ;
  RECT 802.200 3.880 804.680 5.600 ;
  LAYER VI2 ;
  RECT 794.840 3.880 799.580 5.600 ;
  LAYER VI2 ;
  RECT 781.000 3.880 784.840 5.600 ;
  LAYER VI2 ;
  RECT 773.760 3.880 778.500 5.600 ;
  LAYER VI2 ;
  RECT 761.000 3.880 763.760 5.600 ;
  LAYER VI2 ;
  RECT 753.920 3.880 758.660 5.600 ;
  LAYER VI2 ;
  RECT 740.200 3.880 743.920 5.600 ;
  LAYER VI2 ;
  RECT 732.840 3.880 737.580 5.600 ;
  LAYER VI2 ;
  RECT 720.200 3.880 722.840 5.600 ;
  LAYER VI2 ;
  RECT 713.000 3.880 717.740 5.600 ;
  LAYER VI2 ;
  RECT 699.000 3.880 703.000 5.600 ;
  LAYER VI2 ;
  RECT 691.920 3.880 696.660 5.600 ;
  LAYER VI2 ;
  RECT 679.400 3.880 681.920 5.600 ;
  LAYER VI2 ;
  RECT 672.080 3.880 676.820 5.600 ;
  LAYER VI2 ;
  RECT 658.200 3.880 662.080 5.600 ;
  LAYER VI2 ;
  RECT 651.000 3.880 655.740 5.600 ;
  LAYER VI2 ;
  RECT 638.200 3.880 641.000 5.600 ;
  LAYER VI2 ;
  RECT 631.160 3.880 635.900 5.600 ;
  LAYER VI2 ;
  RECT 617.400 3.880 621.160 5.600 ;
  LAYER VI2 ;
  RECT 610.080 3.880 614.820 5.600 ;
  LAYER VI2 ;
  RECT 597.400 3.880 600.080 5.600 ;
  LAYER VI2 ;
  RECT 590.240 3.880 594.980 5.600 ;
  LAYER VI2 ;
  RECT 576.200 3.880 580.240 5.600 ;
  LAYER VI2 ;
  RECT 569.160 3.880 573.900 5.600 ;
  LAYER VI2 ;
  RECT 556.600 3.880 559.160 5.600 ;
  LAYER VI2 ;
  RECT 549.320 3.880 554.060 5.600 ;
  LAYER VI2 ;
  RECT 535.400 3.880 539.320 5.600 ;
  LAYER VI2 ;
  RECT 528.240 3.880 532.980 5.600 ;
  LAYER VI2 ;
  RECT 515.800 3.880 518.240 5.600 ;
  LAYER VI2 ;
  RECT 508.400 3.880 513.140 5.600 ;
  LAYER VI2 ;
  RECT 494.600 3.880 498.400 5.600 ;
  LAYER VI2 ;
  RECT 487.320 3.880 492.060 5.600 ;
  LAYER VI2 ;
  RECT 474.600 3.880 477.320 5.600 ;
  LAYER VI2 ;
  RECT 467.480 3.880 472.220 5.600 ;
  LAYER VI2 ;
  RECT 453.800 3.880 457.480 5.600 ;
  LAYER VI2 ;
  RECT 446.400 3.880 451.140 5.600 ;
  LAYER VI2 ;
  RECT 433.800 3.880 436.400 5.600 ;
  LAYER VI2 ;
  RECT 426.560 3.880 431.300 5.600 ;
  LAYER VI2 ;
  RECT 412.600 3.880 416.560 5.600 ;
  LAYER VI2 ;
  RECT 405.480 3.880 410.220 5.600 ;
  LAYER VI2 ;
  RECT 393.000 3.880 395.480 5.600 ;
  LAYER VI2 ;
  RECT 385.640 3.880 390.380 5.600 ;
  LAYER VI2 ;
  RECT 371.800 3.880 375.640 5.600 ;
  LAYER VI2 ;
  RECT 364.560 3.880 369.300 5.600 ;
  LAYER VI2 ;
  RECT 351.800 3.880 354.560 5.600 ;
  LAYER VI2 ;
  RECT 344.720 3.880 349.460 5.600 ;
  LAYER VI2 ;
  RECT 331.000 3.880 334.720 5.600 ;
  LAYER VI2 ;
  RECT 323.640 3.880 328.380 5.600 ;
  LAYER VI2 ;
  RECT 311.000 3.880 313.640 5.600 ;
  LAYER VI2 ;
  RECT 303.800 3.880 308.540 5.600 ;
  LAYER VI2 ;
  RECT 289.800 3.880 293.800 5.600 ;
  LAYER VI2 ;
  RECT 282.720 3.880 287.460 5.600 ;
  LAYER VI2 ;
  RECT 270.200 3.880 272.720 5.600 ;
  LAYER VI2 ;
  RECT 262.880 3.880 267.620 5.600 ;
  LAYER VI2 ;
  RECT 249.000 3.880 252.880 5.600 ;
  LAYER VI2 ;
  RECT 241.800 3.880 246.540 5.600 ;
  LAYER VI2 ;
  RECT 229.000 3.880 231.800 5.600 ;
  LAYER VI2 ;
  RECT 221.960 3.880 226.700 5.600 ;
  LAYER VI2 ;
  RECT 208.200 3.880 211.960 5.600 ;
  LAYER VI2 ;
  RECT 200.880 3.880 205.620 5.600 ;
  LAYER VI2 ;
  RECT 188.200 3.880 190.880 5.600 ;
  LAYER VI2 ;
  RECT 181.040 3.880 185.780 5.600 ;
  LAYER VI2 ;
  RECT 167.000 3.880 171.040 5.600 ;
  LAYER VI2 ;
  RECT 159.960 3.880 164.700 5.600 ;
  LAYER VI2 ;
  RECT 147.400 3.880 149.960 5.600 ;
  LAYER VI2 ;
  RECT 140.120 3.880 144.860 5.600 ;
  LAYER VI2 ;
  RECT 126.200 3.880 130.120 5.600 ;
  LAYER VI2 ;
  RECT 119.040 3.880 123.780 5.600 ;
  LAYER VI2 ;
  RECT 106.600 3.880 109.040 5.600 ;
  LAYER VI2 ;
  RECT 99.200 3.880 103.940 5.600 ;
  LAYER VI2 ;
  RECT 85.400 3.880 89.200 5.600 ;
  LAYER VI2 ;
  RECT 78.120 3.880 82.860 5.600 ;
  LAYER VI2 ;
  RECT 65.400 3.880 68.120 5.600 ;
  LAYER VI2 ;
  RECT 58.280 3.880 63.020 5.600 ;
  LAYER VI2 ;
  RECT 44.600 3.880 48.280 5.600 ;
  LAYER VI2 ;
  RECT 37.200 3.880 41.940 5.600 ;
  LAYER VI2 ;
  RECT 24.600 3.880 27.200 5.600 ;
  LAYER VI2 ;
  RECT 17.360 3.880 22.100 5.600 ;
  LAYER VI1 ;
  RECT 2674.600 3.740 2680.940 5.600 ;
  LAYER VI1 ;
  RECT 2660.200 3.740 2672.280 5.600 ;
  LAYER VI1 ;
  RECT 2655.000 3.740 2657.650 5.600 ;
  LAYER VI1 ;
  RECT 2640.200 3.740 2652.440 5.600 ;
  LAYER VI1 ;
  RECT 2633.800 3.740 2637.810 5.600 ;
  LAYER VI1 ;
  RECT 2619.400 3.740 2631.360 5.600 ;
  LAYER VI1 ;
  RECT 2614.200 3.740 2616.730 5.600 ;
  LAYER VI1 ;
  RECT 2599.400 3.740 2611.520 5.600 ;
  LAYER VI1 ;
  RECT 2593.000 3.740 2596.890 5.600 ;
  LAYER VI1 ;
  RECT 2578.200 3.740 2590.440 5.600 ;
  LAYER VI1 ;
  RECT 2573.000 3.740 2575.810 5.600 ;
  LAYER VI1 ;
  RECT 2558.600 3.740 2570.600 5.600 ;
  LAYER VI1 ;
  RECT 2552.200 3.740 2555.970 5.600 ;
  LAYER VI1 ;
  RECT 2537.400 3.740 2549.520 5.600 ;
  LAYER VI1 ;
  RECT 2532.200 3.740 2534.890 5.600 ;
  LAYER VI1 ;
  RECT 2517.400 3.740 2529.680 5.600 ;
  LAYER VI1 ;
  RECT 2511.000 3.740 2515.050 5.600 ;
  LAYER VI1 ;
  RECT 2496.600 3.740 2508.600 5.600 ;
  LAYER VI1 ;
  RECT 2491.400 3.740 2493.970 5.600 ;
  LAYER VI1 ;
  RECT 2476.600 3.740 2488.760 5.600 ;
  LAYER VI1 ;
  RECT 2470.200 3.740 2474.130 5.600 ;
  LAYER VI1 ;
  RECT 2455.400 3.740 2467.680 5.600 ;
  LAYER VI1 ;
  RECT 2450.200 3.740 2453.050 5.600 ;
  LAYER VI1 ;
  RECT 2435.800 3.740 2447.840 5.600 ;
  LAYER VI1 ;
  RECT 2429.400 3.740 2433.210 5.600 ;
  LAYER VI1 ;
  RECT 2414.600 3.740 2426.760 5.600 ;
  LAYER VI1 ;
  RECT 2409.400 3.740 2412.130 5.600 ;
  LAYER VI1 ;
  RECT 2394.600 3.740 2406.920 5.600 ;
  LAYER VI1 ;
  RECT 2388.200 3.740 2392.290 5.600 ;
  LAYER VI1 ;
  RECT 2373.800 3.740 2385.840 5.600 ;
  LAYER VI1 ;
  RECT 2368.600 3.740 2371.210 5.600 ;
  LAYER VI1 ;
  RECT 2355.400 3.740 2366.000 5.600 ;
  LAYER VI1 ;
  RECT 2347.400 3.740 2351.370 5.600 ;
  LAYER VI1 ;
  RECT 2332.600 3.740 2344.920 5.600 ;
  LAYER VI1 ;
  RECT 2327.400 3.740 2330.290 5.600 ;
  LAYER VI1 ;
  RECT 2313.000 3.740 2325.080 5.600 ;
  LAYER VI1 ;
  RECT 2306.600 3.740 2310.450 5.600 ;
  LAYER VI1 ;
  RECT 2291.800 3.740 2304.000 5.600 ;
  LAYER VI1 ;
  RECT 2286.600 3.740 2289.370 5.600 ;
  LAYER VI1 ;
  RECT 2272.200 3.740 2284.160 5.600 ;
  LAYER VI1 ;
  RECT 2265.400 3.740 2269.530 5.600 ;
  LAYER VI1 ;
  RECT 2251.000 3.740 2263.080 5.600 ;
  LAYER VI1 ;
  RECT 2245.800 3.740 2248.450 5.600 ;
  LAYER VI1 ;
  RECT 2231.000 3.740 2243.240 5.600 ;
  LAYER VI1 ;
  RECT 2224.600 3.740 2228.610 5.600 ;
  LAYER VI1 ;
  RECT 2210.200 3.740 2222.160 5.600 ;
  LAYER VI1 ;
  RECT 2205.000 3.740 2207.530 5.600 ;
  LAYER VI1 ;
  RECT 2190.200 3.740 2202.320 5.600 ;
  LAYER VI1 ;
  RECT 2183.800 3.740 2187.690 5.600 ;
  LAYER VI1 ;
  RECT 2169.000 3.740 2181.240 5.600 ;
  LAYER VI1 ;
  RECT 2163.800 3.740 2166.610 5.600 ;
  LAYER VI1 ;
  RECT 2149.400 3.740 2161.400 5.600 ;
  LAYER VI1 ;
  RECT 2143.000 3.740 2146.770 5.600 ;
  LAYER VI1 ;
  RECT 2128.200 3.740 2140.320 5.600 ;
  LAYER VI1 ;
  RECT 2123.000 3.740 2125.690 5.600 ;
  LAYER VI1 ;
  RECT 2108.200 3.740 2120.480 5.600 ;
  LAYER VI1 ;
  RECT 2101.800 3.740 2105.850 5.600 ;
  LAYER VI1 ;
  RECT 2087.400 3.740 2099.400 5.600 ;
  LAYER VI1 ;
  RECT 2082.200 3.740 2084.770 5.600 ;
  LAYER VI1 ;
  RECT 2067.400 3.740 2079.560 5.600 ;
  LAYER VI1 ;
  RECT 2061.000 3.740 2064.930 5.600 ;
  LAYER VI1 ;
  RECT 2046.200 3.740 2058.480 5.600 ;
  LAYER VI1 ;
  RECT 2041.000 3.740 2043.850 5.600 ;
  LAYER VI1 ;
  RECT 2028.200 3.740 2038.640 5.600 ;
  LAYER VI1 ;
  RECT 2020.200 3.740 2024.010 5.600 ;
  LAYER VI1 ;
  RECT 2005.400 3.740 2017.560 5.600 ;
  LAYER VI1 ;
  RECT 2000.200 3.740 2002.930 5.600 ;
  LAYER VI1 ;
  RECT 1985.400 3.740 1997.720 5.600 ;
  LAYER VI1 ;
  RECT 1979.000 3.740 1983.090 5.600 ;
  LAYER VI1 ;
  RECT 1964.600 3.740 1976.640 5.600 ;
  LAYER VI1 ;
  RECT 1959.400 3.740 1962.010 5.600 ;
  LAYER VI1 ;
  RECT 1944.600 3.740 1956.800 5.600 ;
  LAYER VI1 ;
  RECT 1938.200 3.740 1942.170 5.600 ;
  LAYER VI1 ;
  RECT 1923.400 3.740 1935.720 5.600 ;
  LAYER VI1 ;
  RECT 1918.200 3.740 1921.090 5.600 ;
  LAYER VI1 ;
  RECT 1903.800 3.740 1915.880 5.600 ;
  LAYER VI1 ;
  RECT 1897.400 3.740 1901.250 5.600 ;
  LAYER VI1 ;
  RECT 1882.600 3.740 1894.800 5.600 ;
  LAYER VI1 ;
  RECT 1877.400 3.740 1880.170 5.600 ;
  LAYER VI1 ;
  RECT 1863.000 3.740 1874.960 5.600 ;
  LAYER VI1 ;
  RECT 1856.200 3.740 1860.330 5.600 ;
  LAYER VI1 ;
  RECT 1841.800 3.740 1853.880 5.600 ;
  LAYER VI1 ;
  RECT 1836.600 3.740 1839.250 5.600 ;
  LAYER VI1 ;
  RECT 1821.800 3.740 1834.040 5.600 ;
  LAYER VI1 ;
  RECT 1815.400 3.740 1819.410 5.600 ;
  LAYER VI1 ;
  RECT 1801.000 3.740 1812.960 5.600 ;
  LAYER VI1 ;
  RECT 1795.800 3.740 1798.330 5.600 ;
  LAYER VI1 ;
  RECT 1781.000 3.740 1793.120 5.600 ;
  LAYER VI1 ;
  RECT 1774.600 3.740 1778.490 5.600 ;
  LAYER VI1 ;
  RECT 1759.800 3.740 1772.040 5.600 ;
  LAYER VI1 ;
  RECT 1754.600 3.740 1757.410 5.600 ;
  LAYER VI1 ;
  RECT 1740.200 3.740 1752.200 5.600 ;
  LAYER VI1 ;
  RECT 1733.800 3.740 1737.570 5.600 ;
  LAYER VI1 ;
  RECT 1719.000 3.740 1731.120 5.600 ;
  LAYER VI1 ;
  RECT 1713.800 3.740 1716.490 5.600 ;
  LAYER VI1 ;
  RECT 1701.000 3.740 1711.280 5.600 ;
  LAYER VI1 ;
  RECT 1692.600 3.740 1696.650 5.600 ;
  LAYER VI1 ;
  RECT 1678.200 3.740 1690.200 5.600 ;
  LAYER VI1 ;
  RECT 1673.000 3.740 1675.570 5.600 ;
  LAYER VI1 ;
  RECT 1658.200 3.740 1670.360 5.600 ;
  LAYER VI1 ;
  RECT 1651.800 3.740 1655.730 5.600 ;
  LAYER VI1 ;
  RECT 1637.000 3.740 1649.280 5.600 ;
  LAYER VI1 ;
  RECT 1631.800 3.740 1634.650 5.600 ;
  LAYER VI1 ;
  RECT 1617.400 3.740 1629.440 5.600 ;
  LAYER VI1 ;
  RECT 1611.000 3.740 1614.810 5.600 ;
  LAYER VI1 ;
  RECT 1596.200 3.740 1608.360 5.600 ;
  LAYER VI1 ;
  RECT 1591.000 3.740 1593.730 5.600 ;
  LAYER VI1 ;
  RECT 1576.200 3.740 1588.520 5.600 ;
  LAYER VI1 ;
  RECT 1569.800 3.740 1573.890 5.600 ;
  LAYER VI1 ;
  RECT 1555.400 3.740 1567.440 5.600 ;
  LAYER VI1 ;
  RECT 1550.200 3.740 1552.810 5.600 ;
  LAYER VI1 ;
  RECT 1535.400 3.740 1547.600 5.600 ;
  LAYER VI1 ;
  RECT 1529.000 3.740 1532.970 5.600 ;
  LAYER VI1 ;
  RECT 1514.200 3.740 1526.520 5.600 ;
  LAYER VI1 ;
  RECT 1509.000 3.740 1511.890 5.600 ;
  LAYER VI1 ;
  RECT 1494.600 3.740 1506.680 5.600 ;
  LAYER VI1 ;
  RECT 1488.200 3.740 1492.050 5.600 ;
  LAYER VI1 ;
  RECT 1473.400 3.740 1485.600 5.600 ;
  LAYER VI1 ;
  RECT 1468.200 3.740 1470.970 5.600 ;
  LAYER VI1 ;
  RECT 1453.800 3.740 1465.760 5.600 ;
  LAYER VI1 ;
  RECT 1447.000 3.740 1451.130 5.600 ;
  LAYER VI1 ;
  RECT 1432.600 3.740 1444.680 5.600 ;
  LAYER VI1 ;
  RECT 1427.400 3.740 1430.050 5.600 ;
  LAYER VI1 ;
  RECT 1412.600 3.740 1424.840 5.600 ;
  LAYER VI1 ;
  RECT 1406.200 3.740 1410.210 5.600 ;
  LAYER VI1 ;
  RECT 1391.800 3.740 1403.760 5.600 ;
  LAYER VI1 ;
  RECT 1386.600 3.740 1389.130 5.600 ;
  LAYER VI1 ;
  RECT 1373.400 3.740 1383.920 5.600 ;
  LAYER VI1 ;
  RECT 1351.000 3.740 1369.290 5.600 ;
  LAYER VI1 ;
  RECT 1339.000 3.740 1342.450 5.600 ;
  LAYER VI1 ;
  RECT 1331.800 3.740 1336.480 5.600 ;
  LAYER VI1 ;
  RECT 1313.000 3.740 1317.360 5.600 ;
  LAYER VI1 ;
  RECT 1298.200 3.740 1310.460 5.600 ;
  LAYER VI1 ;
  RECT 1293.000 3.740 1295.830 5.600 ;
  LAYER VI1 ;
  RECT 1278.600 3.740 1290.620 5.600 ;
  LAYER VI1 ;
  RECT 1272.200 3.740 1275.990 5.600 ;
  LAYER VI1 ;
  RECT 1257.400 3.740 1269.540 5.600 ;
  LAYER VI1 ;
  RECT 1252.200 3.740 1254.910 5.600 ;
  LAYER VI1 ;
  RECT 1237.400 3.740 1249.700 5.600 ;
  LAYER VI1 ;
  RECT 1231.000 3.740 1235.070 5.600 ;
  LAYER VI1 ;
  RECT 1216.600 3.740 1228.620 5.600 ;
  LAYER VI1 ;
  RECT 1211.400 3.740 1213.990 5.600 ;
  LAYER VI1 ;
  RECT 1196.600 3.740 1208.780 5.600 ;
  LAYER VI1 ;
  RECT 1190.200 3.740 1194.150 5.600 ;
  LAYER VI1 ;
  RECT 1175.400 3.740 1187.700 5.600 ;
  LAYER VI1 ;
  RECT 1170.200 3.740 1173.070 5.600 ;
  LAYER VI1 ;
  RECT 1155.800 3.740 1167.860 5.600 ;
  LAYER VI1 ;
  RECT 1149.400 3.740 1153.230 5.600 ;
  LAYER VI1 ;
  RECT 1134.600 3.740 1146.780 5.600 ;
  LAYER VI1 ;
  RECT 1129.400 3.740 1132.150 5.600 ;
  LAYER VI1 ;
  RECT 1115.000 3.740 1126.940 5.600 ;
  LAYER VI1 ;
  RECT 1108.200 3.740 1112.310 5.600 ;
  LAYER VI1 ;
  RECT 1093.800 3.740 1105.860 5.600 ;
  LAYER VI1 ;
  RECT 1088.600 3.740 1091.230 5.600 ;
  LAYER VI1 ;
  RECT 1073.800 3.740 1086.020 5.600 ;
  LAYER VI1 ;
  RECT 1067.400 3.740 1071.390 5.600 ;
  LAYER VI1 ;
  RECT 1053.000 3.740 1064.940 5.600 ;
  LAYER VI1 ;
  RECT 1047.400 3.740 1050.310 5.600 ;
  LAYER VI1 ;
  RECT 1033.000 3.740 1045.100 5.600 ;
  LAYER VI1 ;
  RECT 1026.600 3.740 1030.470 5.600 ;
  LAYER VI1 ;
  RECT 1011.800 3.740 1024.020 5.600 ;
  LAYER VI1 ;
  RECT 1006.600 3.740 1009.390 5.600 ;
  LAYER VI1 ;
  RECT 993.800 3.740 1004.180 5.600 ;
  LAYER VI1 ;
  RECT 985.400 3.740 989.550 5.600 ;
  LAYER VI1 ;
  RECT 971.000 3.740 983.100 5.600 ;
  LAYER VI1 ;
  RECT 965.800 3.740 968.470 5.600 ;
  LAYER VI1 ;
  RECT 951.000 3.740 963.260 5.600 ;
  LAYER VI1 ;
  RECT 944.600 3.740 948.630 5.600 ;
  LAYER VI1 ;
  RECT 930.200 3.740 942.180 5.600 ;
  LAYER VI1 ;
  RECT 925.000 3.740 927.550 5.600 ;
  LAYER VI1 ;
  RECT 910.200 3.740 922.340 5.600 ;
  LAYER VI1 ;
  RECT 903.800 3.740 907.710 5.600 ;
  LAYER VI1 ;
  RECT 889.000 3.740 901.260 5.600 ;
  LAYER VI1 ;
  RECT 883.800 3.740 886.630 5.600 ;
  LAYER VI1 ;
  RECT 869.400 3.740 881.420 5.600 ;
  LAYER VI1 ;
  RECT 863.000 3.740 866.790 5.600 ;
  LAYER VI1 ;
  RECT 848.200 3.740 860.340 5.600 ;
  LAYER VI1 ;
  RECT 843.000 3.740 845.710 5.600 ;
  LAYER VI1 ;
  RECT 828.200 3.740 840.500 5.600 ;
  LAYER VI1 ;
  RECT 821.800 3.740 825.870 5.600 ;
  LAYER VI1 ;
  RECT 807.400 3.740 819.420 5.600 ;
  LAYER VI1 ;
  RECT 802.200 3.740 804.790 5.600 ;
  LAYER VI1 ;
  RECT 787.400 3.740 799.580 5.600 ;
  LAYER VI1 ;
  RECT 781.000 3.740 784.950 5.600 ;
  LAYER VI1 ;
  RECT 766.200 3.740 778.500 5.600 ;
  LAYER VI1 ;
  RECT 761.000 3.740 763.870 5.600 ;
  LAYER VI1 ;
  RECT 746.600 3.740 758.660 5.600 ;
  LAYER VI1 ;
  RECT 740.200 3.740 744.030 5.600 ;
  LAYER VI1 ;
  RECT 725.400 3.740 737.580 5.600 ;
  LAYER VI1 ;
  RECT 720.200 3.740 722.950 5.600 ;
  LAYER VI1 ;
  RECT 705.800 3.740 717.740 5.600 ;
  LAYER VI1 ;
  RECT 699.000 3.740 703.110 5.600 ;
  LAYER VI1 ;
  RECT 684.600 3.740 696.660 5.600 ;
  LAYER VI1 ;
  RECT 679.400 3.740 682.030 5.600 ;
  LAYER VI1 ;
  RECT 666.600 3.740 676.820 5.600 ;
  LAYER VI1 ;
  RECT 658.200 3.740 662.190 5.600 ;
  LAYER VI1 ;
  RECT 643.800 3.740 655.740 5.600 ;
  LAYER VI1 ;
  RECT 638.200 3.740 641.110 5.600 ;
  LAYER VI1 ;
  RECT 623.800 3.740 635.900 5.600 ;
  LAYER VI1 ;
  RECT 617.400 3.740 621.270 5.600 ;
  LAYER VI1 ;
  RECT 602.600 3.740 614.820 5.600 ;
  LAYER VI1 ;
  RECT 597.400 3.740 600.190 5.600 ;
  LAYER VI1 ;
  RECT 583.000 3.740 594.980 5.600 ;
  LAYER VI1 ;
  RECT 576.200 3.740 580.350 5.600 ;
  LAYER VI1 ;
  RECT 561.800 3.740 573.900 5.600 ;
  LAYER VI1 ;
  RECT 556.600 3.740 559.270 5.600 ;
  LAYER VI1 ;
  RECT 541.800 3.740 554.060 5.600 ;
  LAYER VI1 ;
  RECT 535.400 3.740 539.430 5.600 ;
  LAYER VI1 ;
  RECT 521.000 3.740 532.980 5.600 ;
  LAYER VI1 ;
  RECT 515.800 3.740 518.350 5.600 ;
  LAYER VI1 ;
  RECT 501.000 3.740 513.140 5.600 ;
  LAYER VI1 ;
  RECT 494.600 3.740 498.510 5.600 ;
  LAYER VI1 ;
  RECT 479.800 3.740 492.060 5.600 ;
  LAYER VI1 ;
  RECT 474.600 3.740 477.430 5.600 ;
  LAYER VI1 ;
  RECT 460.200 3.740 472.220 5.600 ;
  LAYER VI1 ;
  RECT 453.800 3.740 457.590 5.600 ;
  LAYER VI1 ;
  RECT 439.000 3.740 451.140 5.600 ;
  LAYER VI1 ;
  RECT 433.800 3.740 436.510 5.600 ;
  LAYER VI1 ;
  RECT 419.000 3.740 431.300 5.600 ;
  LAYER VI1 ;
  RECT 412.600 3.740 416.670 5.600 ;
  LAYER VI1 ;
  RECT 398.200 3.740 410.220 5.600 ;
  LAYER VI1 ;
  RECT 393.000 3.740 395.590 5.600 ;
  LAYER VI1 ;
  RECT 378.200 3.740 390.380 5.600 ;
  LAYER VI1 ;
  RECT 371.800 3.740 375.750 5.600 ;
  LAYER VI1 ;
  RECT 357.000 3.740 369.300 5.600 ;
  LAYER VI1 ;
  RECT 351.800 3.740 354.670 5.600 ;
  LAYER VI1 ;
  RECT 339.000 3.740 349.460 5.600 ;
  LAYER VI1 ;
  RECT 331.000 3.740 334.830 5.600 ;
  LAYER VI1 ;
  RECT 316.200 3.740 328.380 5.600 ;
  LAYER VI1 ;
  RECT 311.000 3.740 313.750 5.600 ;
  LAYER VI1 ;
  RECT 296.600 3.740 308.540 5.600 ;
  LAYER VI1 ;
  RECT 289.800 3.740 293.910 5.600 ;
  LAYER VI1 ;
  RECT 275.400 3.740 287.460 5.600 ;
  LAYER VI1 ;
  RECT 270.200 3.740 272.830 5.600 ;
  LAYER VI1 ;
  RECT 255.400 3.740 267.620 5.600 ;
  LAYER VI1 ;
  RECT 249.000 3.740 252.990 5.600 ;
  LAYER VI1 ;
  RECT 234.600 3.740 246.540 5.600 ;
  LAYER VI1 ;
  RECT 229.000 3.740 231.910 5.600 ;
  LAYER VI1 ;
  RECT 214.600 3.740 226.700 5.600 ;
  LAYER VI1 ;
  RECT 208.200 3.740 212.070 5.600 ;
  LAYER VI1 ;
  RECT 193.400 3.740 205.620 5.600 ;
  LAYER VI1 ;
  RECT 188.200 3.740 190.990 5.600 ;
  LAYER VI1 ;
  RECT 173.800 3.740 185.780 5.600 ;
  LAYER VI1 ;
  RECT 167.000 3.740 171.150 5.600 ;
  LAYER VI1 ;
  RECT 152.600 3.740 164.700 5.600 ;
  LAYER VI1 ;
  RECT 147.400 3.740 150.070 5.600 ;
  LAYER VI1 ;
  RECT 132.600 3.740 144.860 5.600 ;
  LAYER VI1 ;
  RECT 126.200 3.740 130.230 5.600 ;
  LAYER VI1 ;
  RECT 111.800 3.740 123.780 5.600 ;
  LAYER VI1 ;
  RECT 106.600 3.740 109.150 5.600 ;
  LAYER VI1 ;
  RECT 91.800 3.740 103.940 5.600 ;
  LAYER VI1 ;
  RECT 85.400 3.740 89.310 5.600 ;
  LAYER VI1 ;
  RECT 70.600 3.740 82.860 5.600 ;
  LAYER VI1 ;
  RECT 65.400 3.740 68.230 5.600 ;
  LAYER VI1 ;
  RECT 51.000 3.740 63.020 5.600 ;
  LAYER VI1 ;
  RECT 44.600 3.740 48.390 5.600 ;
  LAYER VI1 ;
  RECT 29.800 3.740 41.940 5.600 ;
  LAYER VI1 ;
  RECT 24.600 3.740 27.310 5.600 ;
  LAYER VI1 ;
  RECT 11.800 3.740 22.100 5.600 ;
  LAYER VI1 ;
  RECT 4.000 3.740 7.470 5.600 ;
  LAYER VI3 ;
  RECT 2.280 193.930 4.000 195.650 ;
  LAYER VI2 ;
  RECT 2.280 193.930 4.000 195.650 ;
  LAYER VI1 ;
  RECT 2.140 193.930 4.000 195.790 ;
  LAYER VI2 ;
  RECT 0.000 196.070 1.860 197.930 ;
  LAYER VI1 ;
  RECT 0.000 196.070 1.860 197.930 ;
  LAYER VI3 ;
  RECT 2680.940 3.880 2682.660 5.600 ;
  LAYER VI2 ;
  RECT 2680.940 3.880 2682.660 5.600 ;
  LAYER VI1 ;
  RECT 2680.940 3.740 2682.800 5.600 ;
  LAYER VI2 ;
  RECT 2683.080 1.600 2684.940 3.460 ;
  LAYER VI1 ;
  RECT 2683.080 1.600 2684.940 3.460 ;
  LAYER VI3 ;
  RECT 2680.940 193.930 2682.660 195.650 ;
  LAYER VI2 ;
  RECT 2680.940 193.930 2682.660 195.650 ;
  LAYER VI1 ;
  RECT 2680.940 193.930 2682.800 195.790 ;
  LAYER VI2 ;
  RECT 2683.080 196.070 2684.940 197.930 ;
  LAYER VI1 ;
  RECT 2683.080 196.070 2684.940 197.930 ;
  LAYER VI3 ;
  RECT 2.280 3.880 4.000 5.600 ;
  LAYER VI2 ;
  RECT 2.280 3.880 4.000 5.600 ;
  LAYER VI1 ;
  RECT 2.140 3.740 4.000 5.600 ;
  LAYER VI2 ;
  RECT 0.000 1.600 1.860 3.460 ;
  LAYER VI1 ;
  RECT 0.000 1.600 1.860 3.460 ;
  LAYER VI1 ;
  RECT 2672.800 0.200 2673.600 1.000 ;
  LAYER VI2 ;
  RECT 2672.800 0.200 2673.600 1.000 ;
  LAYER VI3 ;
  RECT 2672.800 0.200 2673.600 1.000 ;
  LAYER VI1 ;
  RECT 2658.400 0.200 2659.200 1.000 ;
  LAYER VI2 ;
  RECT 2658.400 0.200 2659.200 1.000 ;
  LAYER VI3 ;
  RECT 2658.400 0.200 2659.200 1.000 ;
  LAYER VI1 ;
  RECT 2653.200 0.200 2654.000 1.000 ;
  LAYER VI2 ;
  RECT 2653.200 0.200 2654.000 1.000 ;
  LAYER VI3 ;
  RECT 2653.200 0.200 2654.000 1.000 ;
  LAYER VI1 ;
  RECT 2638.400 0.200 2639.200 1.000 ;
  LAYER VI2 ;
  RECT 2638.400 0.200 2639.200 1.000 ;
  LAYER VI3 ;
  RECT 2638.400 0.200 2639.200 1.000 ;
  LAYER VI1 ;
  RECT 2632.000 0.200 2632.800 1.000 ;
  LAYER VI2 ;
  RECT 2632.000 0.200 2632.800 1.000 ;
  LAYER VI3 ;
  RECT 2632.000 0.200 2632.800 1.000 ;
  LAYER VI1 ;
  RECT 2617.600 0.200 2618.400 1.000 ;
  LAYER VI2 ;
  RECT 2617.600 0.200 2618.400 1.000 ;
  LAYER VI3 ;
  RECT 2617.600 0.200 2618.400 1.000 ;
  LAYER VI1 ;
  RECT 2612.400 0.200 2613.200 1.000 ;
  LAYER VI2 ;
  RECT 2612.400 0.200 2613.200 1.000 ;
  LAYER VI3 ;
  RECT 2612.400 0.200 2613.200 1.000 ;
  LAYER VI1 ;
  RECT 2597.600 0.200 2598.400 1.000 ;
  LAYER VI2 ;
  RECT 2597.600 0.200 2598.400 1.000 ;
  LAYER VI3 ;
  RECT 2597.600 0.200 2598.400 1.000 ;
  LAYER VI1 ;
  RECT 2591.200 0.200 2592.000 1.000 ;
  LAYER VI2 ;
  RECT 2591.200 0.200 2592.000 1.000 ;
  LAYER VI3 ;
  RECT 2591.200 0.200 2592.000 1.000 ;
  LAYER VI1 ;
  RECT 2576.400 0.200 2577.200 1.000 ;
  LAYER VI2 ;
  RECT 2576.400 0.200 2577.200 1.000 ;
  LAYER VI3 ;
  RECT 2576.400 0.200 2577.200 1.000 ;
  LAYER VI1 ;
  RECT 2571.200 0.200 2572.000 1.000 ;
  LAYER VI2 ;
  RECT 2571.200 0.200 2572.000 1.000 ;
  LAYER VI3 ;
  RECT 2571.200 0.200 2572.000 1.000 ;
  LAYER VI1 ;
  RECT 2556.800 0.200 2557.600 1.000 ;
  LAYER VI2 ;
  RECT 2556.800 0.200 2557.600 1.000 ;
  LAYER VI3 ;
  RECT 2556.800 0.200 2557.600 1.000 ;
  LAYER VI1 ;
  RECT 2550.400 0.200 2551.200 1.000 ;
  LAYER VI2 ;
  RECT 2550.400 0.200 2551.200 1.000 ;
  LAYER VI3 ;
  RECT 2550.400 0.200 2551.200 1.000 ;
  LAYER VI1 ;
  RECT 2535.600 0.200 2536.400 1.000 ;
  LAYER VI2 ;
  RECT 2535.600 0.200 2536.400 1.000 ;
  LAYER VI3 ;
  RECT 2535.600 0.200 2536.400 1.000 ;
  LAYER VI1 ;
  RECT 2530.400 0.200 2531.200 1.000 ;
  LAYER VI2 ;
  RECT 2530.400 0.200 2531.200 1.000 ;
  LAYER VI3 ;
  RECT 2530.400 0.200 2531.200 1.000 ;
  LAYER VI1 ;
  RECT 2515.600 0.200 2516.400 1.000 ;
  LAYER VI2 ;
  RECT 2515.600 0.200 2516.400 1.000 ;
  LAYER VI3 ;
  RECT 2515.600 0.200 2516.400 1.000 ;
  LAYER VI1 ;
  RECT 2509.200 0.200 2510.000 1.000 ;
  LAYER VI2 ;
  RECT 2509.200 0.200 2510.000 1.000 ;
  LAYER VI3 ;
  RECT 2509.200 0.200 2510.000 1.000 ;
  LAYER VI1 ;
  RECT 2494.800 0.200 2495.600 1.000 ;
  LAYER VI2 ;
  RECT 2494.800 0.200 2495.600 1.000 ;
  LAYER VI3 ;
  RECT 2494.800 0.200 2495.600 1.000 ;
  LAYER VI1 ;
  RECT 2489.600 0.200 2490.400 1.000 ;
  LAYER VI2 ;
  RECT 2489.600 0.200 2490.400 1.000 ;
  LAYER VI3 ;
  RECT 2489.600 0.200 2490.400 1.000 ;
  LAYER VI1 ;
  RECT 2474.800 0.200 2475.600 1.000 ;
  LAYER VI2 ;
  RECT 2474.800 0.200 2475.600 1.000 ;
  LAYER VI3 ;
  RECT 2474.800 0.200 2475.600 1.000 ;
  LAYER VI1 ;
  RECT 2468.400 0.200 2469.200 1.000 ;
  LAYER VI2 ;
  RECT 2468.400 0.200 2469.200 1.000 ;
  LAYER VI3 ;
  RECT 2468.400 0.200 2469.200 1.000 ;
  LAYER VI1 ;
  RECT 2453.600 0.200 2454.400 1.000 ;
  LAYER VI2 ;
  RECT 2453.600 0.200 2454.400 1.000 ;
  LAYER VI3 ;
  RECT 2453.600 0.200 2454.400 1.000 ;
  LAYER VI1 ;
  RECT 2448.400 0.200 2449.200 1.000 ;
  LAYER VI2 ;
  RECT 2448.400 0.200 2449.200 1.000 ;
  LAYER VI3 ;
  RECT 2448.400 0.200 2449.200 1.000 ;
  LAYER VI1 ;
  RECT 2434.000 0.200 2434.800 1.000 ;
  LAYER VI2 ;
  RECT 2434.000 0.200 2434.800 1.000 ;
  LAYER VI3 ;
  RECT 2434.000 0.200 2434.800 1.000 ;
  LAYER VI1 ;
  RECT 2427.600 0.200 2428.400 1.000 ;
  LAYER VI2 ;
  RECT 2427.600 0.200 2428.400 1.000 ;
  LAYER VI3 ;
  RECT 2427.600 0.200 2428.400 1.000 ;
  LAYER VI1 ;
  RECT 2412.800 0.200 2413.600 1.000 ;
  LAYER VI2 ;
  RECT 2412.800 0.200 2413.600 1.000 ;
  LAYER VI3 ;
  RECT 2412.800 0.200 2413.600 1.000 ;
  LAYER VI1 ;
  RECT 2407.600 0.200 2408.400 1.000 ;
  LAYER VI2 ;
  RECT 2407.600 0.200 2408.400 1.000 ;
  LAYER VI3 ;
  RECT 2407.600 0.200 2408.400 1.000 ;
  LAYER VI1 ;
  RECT 2392.800 0.200 2393.600 1.000 ;
  LAYER VI2 ;
  RECT 2392.800 0.200 2393.600 1.000 ;
  LAYER VI3 ;
  RECT 2392.800 0.200 2393.600 1.000 ;
  LAYER VI1 ;
  RECT 2386.400 0.200 2387.200 1.000 ;
  LAYER VI2 ;
  RECT 2386.400 0.200 2387.200 1.000 ;
  LAYER VI3 ;
  RECT 2386.400 0.200 2387.200 1.000 ;
  LAYER VI1 ;
  RECT 2372.000 0.200 2372.800 1.000 ;
  LAYER VI2 ;
  RECT 2372.000 0.200 2372.800 1.000 ;
  LAYER VI3 ;
  RECT 2372.000 0.200 2372.800 1.000 ;
  LAYER VI1 ;
  RECT 2366.800 0.200 2367.600 1.000 ;
  LAYER VI2 ;
  RECT 2366.800 0.200 2367.600 1.000 ;
  LAYER VI3 ;
  RECT 2366.800 0.200 2367.600 1.000 ;
  LAYER VI1 ;
  RECT 2353.600 0.200 2354.400 1.000 ;
  LAYER VI2 ;
  RECT 2353.600 0.200 2354.400 1.000 ;
  LAYER VI3 ;
  RECT 2353.600 0.200 2354.400 1.000 ;
  LAYER VI1 ;
  RECT 2352.000 0.200 2352.800 1.000 ;
  LAYER VI2 ;
  RECT 2352.000 0.200 2352.800 1.000 ;
  LAYER VI3 ;
  RECT 2352.000 0.200 2352.800 1.000 ;
  LAYER VI1 ;
  RECT 2345.600 0.200 2346.400 1.000 ;
  LAYER VI2 ;
  RECT 2345.600 0.200 2346.400 1.000 ;
  LAYER VI3 ;
  RECT 2345.600 0.200 2346.400 1.000 ;
  LAYER VI1 ;
  RECT 2330.800 0.200 2331.600 1.000 ;
  LAYER VI2 ;
  RECT 2330.800 0.200 2331.600 1.000 ;
  LAYER VI3 ;
  RECT 2330.800 0.200 2331.600 1.000 ;
  LAYER VI1 ;
  RECT 2325.600 0.200 2326.400 1.000 ;
  LAYER VI2 ;
  RECT 2325.600 0.200 2326.400 1.000 ;
  LAYER VI3 ;
  RECT 2325.600 0.200 2326.400 1.000 ;
  LAYER VI1 ;
  RECT 2311.200 0.200 2312.000 1.000 ;
  LAYER VI2 ;
  RECT 2311.200 0.200 2312.000 1.000 ;
  LAYER VI3 ;
  RECT 2311.200 0.200 2312.000 1.000 ;
  LAYER VI1 ;
  RECT 2304.800 0.200 2305.600 1.000 ;
  LAYER VI2 ;
  RECT 2304.800 0.200 2305.600 1.000 ;
  LAYER VI3 ;
  RECT 2304.800 0.200 2305.600 1.000 ;
  LAYER VI1 ;
  RECT 2290.000 0.200 2290.800 1.000 ;
  LAYER VI2 ;
  RECT 2290.000 0.200 2290.800 1.000 ;
  LAYER VI3 ;
  RECT 2290.000 0.200 2290.800 1.000 ;
  LAYER VI1 ;
  RECT 2284.800 0.200 2285.600 1.000 ;
  LAYER VI2 ;
  RECT 2284.800 0.200 2285.600 1.000 ;
  LAYER VI3 ;
  RECT 2284.800 0.200 2285.600 1.000 ;
  LAYER VI1 ;
  RECT 2270.400 0.200 2271.200 1.000 ;
  LAYER VI2 ;
  RECT 2270.400 0.200 2271.200 1.000 ;
  LAYER VI3 ;
  RECT 2270.400 0.200 2271.200 1.000 ;
  LAYER VI1 ;
  RECT 2263.600 0.200 2264.400 1.000 ;
  LAYER VI2 ;
  RECT 2263.600 0.200 2264.400 1.000 ;
  LAYER VI3 ;
  RECT 2263.600 0.200 2264.400 1.000 ;
  LAYER VI1 ;
  RECT 2249.200 0.200 2250.000 1.000 ;
  LAYER VI2 ;
  RECT 2249.200 0.200 2250.000 1.000 ;
  LAYER VI3 ;
  RECT 2249.200 0.200 2250.000 1.000 ;
  LAYER VI1 ;
  RECT 2244.000 0.200 2244.800 1.000 ;
  LAYER VI2 ;
  RECT 2244.000 0.200 2244.800 1.000 ;
  LAYER VI3 ;
  RECT 2244.000 0.200 2244.800 1.000 ;
  LAYER VI1 ;
  RECT 2229.200 0.200 2230.000 1.000 ;
  LAYER VI2 ;
  RECT 2229.200 0.200 2230.000 1.000 ;
  LAYER VI3 ;
  RECT 2229.200 0.200 2230.000 1.000 ;
  LAYER VI1 ;
  RECT 2222.800 0.200 2223.600 1.000 ;
  LAYER VI2 ;
  RECT 2222.800 0.200 2223.600 1.000 ;
  LAYER VI3 ;
  RECT 2222.800 0.200 2223.600 1.000 ;
  LAYER VI1 ;
  RECT 2208.400 0.200 2209.200 1.000 ;
  LAYER VI2 ;
  RECT 2208.400 0.200 2209.200 1.000 ;
  LAYER VI3 ;
  RECT 2208.400 0.200 2209.200 1.000 ;
  LAYER VI1 ;
  RECT 2203.200 0.200 2204.000 1.000 ;
  LAYER VI2 ;
  RECT 2203.200 0.200 2204.000 1.000 ;
  LAYER VI3 ;
  RECT 2203.200 0.200 2204.000 1.000 ;
  LAYER VI1 ;
  RECT 2188.400 0.200 2189.200 1.000 ;
  LAYER VI2 ;
  RECT 2188.400 0.200 2189.200 1.000 ;
  LAYER VI3 ;
  RECT 2188.400 0.200 2189.200 1.000 ;
  LAYER VI1 ;
  RECT 2182.000 0.200 2182.800 1.000 ;
  LAYER VI2 ;
  RECT 2182.000 0.200 2182.800 1.000 ;
  LAYER VI3 ;
  RECT 2182.000 0.200 2182.800 1.000 ;
  LAYER VI1 ;
  RECT 2167.200 0.200 2168.000 1.000 ;
  LAYER VI2 ;
  RECT 2167.200 0.200 2168.000 1.000 ;
  LAYER VI3 ;
  RECT 2167.200 0.200 2168.000 1.000 ;
  LAYER VI1 ;
  RECT 2162.000 0.200 2162.800 1.000 ;
  LAYER VI2 ;
  RECT 2162.000 0.200 2162.800 1.000 ;
  LAYER VI3 ;
  RECT 2162.000 0.200 2162.800 1.000 ;
  LAYER VI1 ;
  RECT 2147.600 0.200 2148.400 1.000 ;
  LAYER VI2 ;
  RECT 2147.600 0.200 2148.400 1.000 ;
  LAYER VI3 ;
  RECT 2147.600 0.200 2148.400 1.000 ;
  LAYER VI1 ;
  RECT 2141.200 0.200 2142.000 1.000 ;
  LAYER VI2 ;
  RECT 2141.200 0.200 2142.000 1.000 ;
  LAYER VI3 ;
  RECT 2141.200 0.200 2142.000 1.000 ;
  LAYER VI1 ;
  RECT 2126.400 0.200 2127.200 1.000 ;
  LAYER VI2 ;
  RECT 2126.400 0.200 2127.200 1.000 ;
  LAYER VI3 ;
  RECT 2126.400 0.200 2127.200 1.000 ;
  LAYER VI1 ;
  RECT 2121.200 0.200 2122.000 1.000 ;
  LAYER VI2 ;
  RECT 2121.200 0.200 2122.000 1.000 ;
  LAYER VI3 ;
  RECT 2121.200 0.200 2122.000 1.000 ;
  LAYER VI1 ;
  RECT 2106.400 0.200 2107.200 1.000 ;
  LAYER VI2 ;
  RECT 2106.400 0.200 2107.200 1.000 ;
  LAYER VI3 ;
  RECT 2106.400 0.200 2107.200 1.000 ;
  LAYER VI1 ;
  RECT 2100.000 0.200 2100.800 1.000 ;
  LAYER VI2 ;
  RECT 2100.000 0.200 2100.800 1.000 ;
  LAYER VI3 ;
  RECT 2100.000 0.200 2100.800 1.000 ;
  LAYER VI1 ;
  RECT 2085.600 0.200 2086.400 1.000 ;
  LAYER VI2 ;
  RECT 2085.600 0.200 2086.400 1.000 ;
  LAYER VI3 ;
  RECT 2085.600 0.200 2086.400 1.000 ;
  LAYER VI1 ;
  RECT 2080.400 0.200 2081.200 1.000 ;
  LAYER VI2 ;
  RECT 2080.400 0.200 2081.200 1.000 ;
  LAYER VI3 ;
  RECT 2080.400 0.200 2081.200 1.000 ;
  LAYER VI1 ;
  RECT 2065.600 0.200 2066.400 1.000 ;
  LAYER VI2 ;
  RECT 2065.600 0.200 2066.400 1.000 ;
  LAYER VI3 ;
  RECT 2065.600 0.200 2066.400 1.000 ;
  LAYER VI1 ;
  RECT 2059.200 0.200 2060.000 1.000 ;
  LAYER VI2 ;
  RECT 2059.200 0.200 2060.000 1.000 ;
  LAYER VI3 ;
  RECT 2059.200 0.200 2060.000 1.000 ;
  LAYER VI1 ;
  RECT 2044.400 0.200 2045.200 1.000 ;
  LAYER VI2 ;
  RECT 2044.400 0.200 2045.200 1.000 ;
  LAYER VI3 ;
  RECT 2044.400 0.200 2045.200 1.000 ;
  LAYER VI1 ;
  RECT 2039.200 0.200 2040.000 1.000 ;
  LAYER VI2 ;
  RECT 2039.200 0.200 2040.000 1.000 ;
  LAYER VI3 ;
  RECT 2039.200 0.200 2040.000 1.000 ;
  LAYER VI1 ;
  RECT 2026.400 0.200 2027.200 1.000 ;
  LAYER VI2 ;
  RECT 2026.400 0.200 2027.200 1.000 ;
  LAYER VI3 ;
  RECT 2026.400 0.200 2027.200 1.000 ;
  LAYER VI1 ;
  RECT 2024.800 0.200 2025.600 1.000 ;
  LAYER VI2 ;
  RECT 2024.800 0.200 2025.600 1.000 ;
  LAYER VI3 ;
  RECT 2024.800 0.200 2025.600 1.000 ;
  LAYER VI1 ;
  RECT 2018.400 0.200 2019.200 1.000 ;
  LAYER VI2 ;
  RECT 2018.400 0.200 2019.200 1.000 ;
  LAYER VI3 ;
  RECT 2018.400 0.200 2019.200 1.000 ;
  LAYER VI1 ;
  RECT 2003.600 0.200 2004.400 1.000 ;
  LAYER VI2 ;
  RECT 2003.600 0.200 2004.400 1.000 ;
  LAYER VI3 ;
  RECT 2003.600 0.200 2004.400 1.000 ;
  LAYER VI1 ;
  RECT 1998.400 0.200 1999.200 1.000 ;
  LAYER VI2 ;
  RECT 1998.400 0.200 1999.200 1.000 ;
  LAYER VI3 ;
  RECT 1998.400 0.200 1999.200 1.000 ;
  LAYER VI1 ;
  RECT 1983.600 0.200 1984.400 1.000 ;
  LAYER VI2 ;
  RECT 1983.600 0.200 1984.400 1.000 ;
  LAYER VI3 ;
  RECT 1983.600 0.200 1984.400 1.000 ;
  LAYER VI1 ;
  RECT 1977.200 0.200 1978.000 1.000 ;
  LAYER VI2 ;
  RECT 1977.200 0.200 1978.000 1.000 ;
  LAYER VI3 ;
  RECT 1977.200 0.200 1978.000 1.000 ;
  LAYER VI1 ;
  RECT 1962.800 0.200 1963.600 1.000 ;
  LAYER VI2 ;
  RECT 1962.800 0.200 1963.600 1.000 ;
  LAYER VI3 ;
  RECT 1962.800 0.200 1963.600 1.000 ;
  LAYER VI1 ;
  RECT 1957.600 0.200 1958.400 1.000 ;
  LAYER VI2 ;
  RECT 1957.600 0.200 1958.400 1.000 ;
  LAYER VI3 ;
  RECT 1957.600 0.200 1958.400 1.000 ;
  LAYER VI1 ;
  RECT 1942.800 0.200 1943.600 1.000 ;
  LAYER VI2 ;
  RECT 1942.800 0.200 1943.600 1.000 ;
  LAYER VI3 ;
  RECT 1942.800 0.200 1943.600 1.000 ;
  LAYER VI1 ;
  RECT 1936.400 0.200 1937.200 1.000 ;
  LAYER VI2 ;
  RECT 1936.400 0.200 1937.200 1.000 ;
  LAYER VI3 ;
  RECT 1936.400 0.200 1937.200 1.000 ;
  LAYER VI1 ;
  RECT 1921.600 0.200 1922.400 1.000 ;
  LAYER VI2 ;
  RECT 1921.600 0.200 1922.400 1.000 ;
  LAYER VI3 ;
  RECT 1921.600 0.200 1922.400 1.000 ;
  LAYER VI1 ;
  RECT 1916.400 0.200 1917.200 1.000 ;
  LAYER VI2 ;
  RECT 1916.400 0.200 1917.200 1.000 ;
  LAYER VI3 ;
  RECT 1916.400 0.200 1917.200 1.000 ;
  LAYER VI1 ;
  RECT 1902.000 0.200 1902.800 1.000 ;
  LAYER VI2 ;
  RECT 1902.000 0.200 1902.800 1.000 ;
  LAYER VI3 ;
  RECT 1902.000 0.200 1902.800 1.000 ;
  LAYER VI1 ;
  RECT 1895.600 0.200 1896.400 1.000 ;
  LAYER VI2 ;
  RECT 1895.600 0.200 1896.400 1.000 ;
  LAYER VI3 ;
  RECT 1895.600 0.200 1896.400 1.000 ;
  LAYER VI1 ;
  RECT 1880.800 0.200 1881.600 1.000 ;
  LAYER VI2 ;
  RECT 1880.800 0.200 1881.600 1.000 ;
  LAYER VI3 ;
  RECT 1880.800 0.200 1881.600 1.000 ;
  LAYER VI1 ;
  RECT 1875.600 0.200 1876.400 1.000 ;
  LAYER VI2 ;
  RECT 1875.600 0.200 1876.400 1.000 ;
  LAYER VI3 ;
  RECT 1875.600 0.200 1876.400 1.000 ;
  LAYER VI1 ;
  RECT 1861.200 0.200 1862.000 1.000 ;
  LAYER VI2 ;
  RECT 1861.200 0.200 1862.000 1.000 ;
  LAYER VI3 ;
  RECT 1861.200 0.200 1862.000 1.000 ;
  LAYER VI1 ;
  RECT 1854.400 0.200 1855.200 1.000 ;
  LAYER VI2 ;
  RECT 1854.400 0.200 1855.200 1.000 ;
  LAYER VI3 ;
  RECT 1854.400 0.200 1855.200 1.000 ;
  LAYER VI1 ;
  RECT 1840.000 0.200 1840.800 1.000 ;
  LAYER VI2 ;
  RECT 1840.000 0.200 1840.800 1.000 ;
  LAYER VI3 ;
  RECT 1840.000 0.200 1840.800 1.000 ;
  LAYER VI1 ;
  RECT 1834.800 0.200 1835.600 1.000 ;
  LAYER VI2 ;
  RECT 1834.800 0.200 1835.600 1.000 ;
  LAYER VI3 ;
  RECT 1834.800 0.200 1835.600 1.000 ;
  LAYER VI1 ;
  RECT 1820.000 0.200 1820.800 1.000 ;
  LAYER VI2 ;
  RECT 1820.000 0.200 1820.800 1.000 ;
  LAYER VI3 ;
  RECT 1820.000 0.200 1820.800 1.000 ;
  LAYER VI1 ;
  RECT 1813.600 0.200 1814.400 1.000 ;
  LAYER VI2 ;
  RECT 1813.600 0.200 1814.400 1.000 ;
  LAYER VI3 ;
  RECT 1813.600 0.200 1814.400 1.000 ;
  LAYER VI1 ;
  RECT 1799.200 0.200 1800.000 1.000 ;
  LAYER VI2 ;
  RECT 1799.200 0.200 1800.000 1.000 ;
  LAYER VI3 ;
  RECT 1799.200 0.200 1800.000 1.000 ;
  LAYER VI1 ;
  RECT 1794.000 0.200 1794.800 1.000 ;
  LAYER VI2 ;
  RECT 1794.000 0.200 1794.800 1.000 ;
  LAYER VI3 ;
  RECT 1794.000 0.200 1794.800 1.000 ;
  LAYER VI1 ;
  RECT 1779.200 0.200 1780.000 1.000 ;
  LAYER VI2 ;
  RECT 1779.200 0.200 1780.000 1.000 ;
  LAYER VI3 ;
  RECT 1779.200 0.200 1780.000 1.000 ;
  LAYER VI1 ;
  RECT 1772.800 0.200 1773.600 1.000 ;
  LAYER VI2 ;
  RECT 1772.800 0.200 1773.600 1.000 ;
  LAYER VI3 ;
  RECT 1772.800 0.200 1773.600 1.000 ;
  LAYER VI1 ;
  RECT 1758.000 0.200 1758.800 1.000 ;
  LAYER VI2 ;
  RECT 1758.000 0.200 1758.800 1.000 ;
  LAYER VI3 ;
  RECT 1758.000 0.200 1758.800 1.000 ;
  LAYER VI1 ;
  RECT 1752.800 0.200 1753.600 1.000 ;
  LAYER VI2 ;
  RECT 1752.800 0.200 1753.600 1.000 ;
  LAYER VI3 ;
  RECT 1752.800 0.200 1753.600 1.000 ;
  LAYER VI1 ;
  RECT 1738.400 0.200 1739.200 1.000 ;
  LAYER VI2 ;
  RECT 1738.400 0.200 1739.200 1.000 ;
  LAYER VI3 ;
  RECT 1738.400 0.200 1739.200 1.000 ;
  LAYER VI1 ;
  RECT 1732.000 0.200 1732.800 1.000 ;
  LAYER VI2 ;
  RECT 1732.000 0.200 1732.800 1.000 ;
  LAYER VI3 ;
  RECT 1732.000 0.200 1732.800 1.000 ;
  LAYER VI1 ;
  RECT 1717.200 0.200 1718.000 1.000 ;
  LAYER VI2 ;
  RECT 1717.200 0.200 1718.000 1.000 ;
  LAYER VI3 ;
  RECT 1717.200 0.200 1718.000 1.000 ;
  LAYER VI1 ;
  RECT 1712.000 0.200 1712.800 1.000 ;
  LAYER VI2 ;
  RECT 1712.000 0.200 1712.800 1.000 ;
  LAYER VI3 ;
  RECT 1712.000 0.200 1712.800 1.000 ;
  LAYER VI1 ;
  RECT 1699.200 0.200 1700.000 1.000 ;
  LAYER VI2 ;
  RECT 1699.200 0.200 1700.000 1.000 ;
  LAYER VI3 ;
  RECT 1699.200 0.200 1700.000 1.000 ;
  LAYER VI1 ;
  RECT 1697.200 0.200 1698.000 1.000 ;
  LAYER VI2 ;
  RECT 1697.200 0.200 1698.000 1.000 ;
  LAYER VI3 ;
  RECT 1697.200 0.200 1698.000 1.000 ;
  LAYER VI1 ;
  RECT 1690.800 0.200 1691.600 1.000 ;
  LAYER VI2 ;
  RECT 1690.800 0.200 1691.600 1.000 ;
  LAYER VI3 ;
  RECT 1690.800 0.200 1691.600 1.000 ;
  LAYER VI1 ;
  RECT 1676.400 0.200 1677.200 1.000 ;
  LAYER VI2 ;
  RECT 1676.400 0.200 1677.200 1.000 ;
  LAYER VI3 ;
  RECT 1676.400 0.200 1677.200 1.000 ;
  LAYER VI1 ;
  RECT 1671.200 0.200 1672.000 1.000 ;
  LAYER VI2 ;
  RECT 1671.200 0.200 1672.000 1.000 ;
  LAYER VI3 ;
  RECT 1671.200 0.200 1672.000 1.000 ;
  LAYER VI1 ;
  RECT 1656.400 0.200 1657.200 1.000 ;
  LAYER VI2 ;
  RECT 1656.400 0.200 1657.200 1.000 ;
  LAYER VI3 ;
  RECT 1656.400 0.200 1657.200 1.000 ;
  LAYER VI1 ;
  RECT 1650.000 0.200 1650.800 1.000 ;
  LAYER VI2 ;
  RECT 1650.000 0.200 1650.800 1.000 ;
  LAYER VI3 ;
  RECT 1650.000 0.200 1650.800 1.000 ;
  LAYER VI1 ;
  RECT 1635.200 0.200 1636.000 1.000 ;
  LAYER VI2 ;
  RECT 1635.200 0.200 1636.000 1.000 ;
  LAYER VI3 ;
  RECT 1635.200 0.200 1636.000 1.000 ;
  LAYER VI1 ;
  RECT 1630.000 0.200 1630.800 1.000 ;
  LAYER VI2 ;
  RECT 1630.000 0.200 1630.800 1.000 ;
  LAYER VI3 ;
  RECT 1630.000 0.200 1630.800 1.000 ;
  LAYER VI1 ;
  RECT 1615.600 0.200 1616.400 1.000 ;
  LAYER VI2 ;
  RECT 1615.600 0.200 1616.400 1.000 ;
  LAYER VI3 ;
  RECT 1615.600 0.200 1616.400 1.000 ;
  LAYER VI1 ;
  RECT 1609.200 0.200 1610.000 1.000 ;
  LAYER VI2 ;
  RECT 1609.200 0.200 1610.000 1.000 ;
  LAYER VI3 ;
  RECT 1609.200 0.200 1610.000 1.000 ;
  LAYER VI1 ;
  RECT 1594.400 0.200 1595.200 1.000 ;
  LAYER VI2 ;
  RECT 1594.400 0.200 1595.200 1.000 ;
  LAYER VI3 ;
  RECT 1594.400 0.200 1595.200 1.000 ;
  LAYER VI1 ;
  RECT 1589.200 0.200 1590.000 1.000 ;
  LAYER VI2 ;
  RECT 1589.200 0.200 1590.000 1.000 ;
  LAYER VI3 ;
  RECT 1589.200 0.200 1590.000 1.000 ;
  LAYER VI1 ;
  RECT 1574.400 0.200 1575.200 1.000 ;
  LAYER VI2 ;
  RECT 1574.400 0.200 1575.200 1.000 ;
  LAYER VI3 ;
  RECT 1574.400 0.200 1575.200 1.000 ;
  LAYER VI1 ;
  RECT 1568.000 0.200 1568.800 1.000 ;
  LAYER VI2 ;
  RECT 1568.000 0.200 1568.800 1.000 ;
  LAYER VI3 ;
  RECT 1568.000 0.200 1568.800 1.000 ;
  LAYER VI1 ;
  RECT 1553.600 0.200 1554.400 1.000 ;
  LAYER VI2 ;
  RECT 1553.600 0.200 1554.400 1.000 ;
  LAYER VI3 ;
  RECT 1553.600 0.200 1554.400 1.000 ;
  LAYER VI1 ;
  RECT 1548.400 0.200 1549.200 1.000 ;
  LAYER VI2 ;
  RECT 1548.400 0.200 1549.200 1.000 ;
  LAYER VI3 ;
  RECT 1548.400 0.200 1549.200 1.000 ;
  LAYER VI1 ;
  RECT 1533.600 0.200 1534.400 1.000 ;
  LAYER VI2 ;
  RECT 1533.600 0.200 1534.400 1.000 ;
  LAYER VI3 ;
  RECT 1533.600 0.200 1534.400 1.000 ;
  LAYER VI1 ;
  RECT 1527.200 0.200 1528.000 1.000 ;
  LAYER VI2 ;
  RECT 1527.200 0.200 1528.000 1.000 ;
  LAYER VI3 ;
  RECT 1527.200 0.200 1528.000 1.000 ;
  LAYER VI1 ;
  RECT 1512.400 0.200 1513.200 1.000 ;
  LAYER VI2 ;
  RECT 1512.400 0.200 1513.200 1.000 ;
  LAYER VI3 ;
  RECT 1512.400 0.200 1513.200 1.000 ;
  LAYER VI1 ;
  RECT 1507.200 0.200 1508.000 1.000 ;
  LAYER VI2 ;
  RECT 1507.200 0.200 1508.000 1.000 ;
  LAYER VI3 ;
  RECT 1507.200 0.200 1508.000 1.000 ;
  LAYER VI1 ;
  RECT 1492.800 0.200 1493.600 1.000 ;
  LAYER VI2 ;
  RECT 1492.800 0.200 1493.600 1.000 ;
  LAYER VI3 ;
  RECT 1492.800 0.200 1493.600 1.000 ;
  LAYER VI1 ;
  RECT 1486.400 0.200 1487.200 1.000 ;
  LAYER VI2 ;
  RECT 1486.400 0.200 1487.200 1.000 ;
  LAYER VI3 ;
  RECT 1486.400 0.200 1487.200 1.000 ;
  LAYER VI1 ;
  RECT 1471.600 0.200 1472.400 1.000 ;
  LAYER VI2 ;
  RECT 1471.600 0.200 1472.400 1.000 ;
  LAYER VI3 ;
  RECT 1471.600 0.200 1472.400 1.000 ;
  LAYER VI1 ;
  RECT 1466.400 0.200 1467.200 1.000 ;
  LAYER VI2 ;
  RECT 1466.400 0.200 1467.200 1.000 ;
  LAYER VI3 ;
  RECT 1466.400 0.200 1467.200 1.000 ;
  LAYER VI1 ;
  RECT 1452.000 0.200 1452.800 1.000 ;
  LAYER VI2 ;
  RECT 1452.000 0.200 1452.800 1.000 ;
  LAYER VI3 ;
  RECT 1452.000 0.200 1452.800 1.000 ;
  LAYER VI1 ;
  RECT 1445.200 0.200 1446.000 1.000 ;
  LAYER VI2 ;
  RECT 1445.200 0.200 1446.000 1.000 ;
  LAYER VI3 ;
  RECT 1445.200 0.200 1446.000 1.000 ;
  LAYER VI1 ;
  RECT 1430.800 0.200 1431.600 1.000 ;
  LAYER VI2 ;
  RECT 1430.800 0.200 1431.600 1.000 ;
  LAYER VI3 ;
  RECT 1430.800 0.200 1431.600 1.000 ;
  LAYER VI1 ;
  RECT 1425.600 0.200 1426.400 1.000 ;
  LAYER VI2 ;
  RECT 1425.600 0.200 1426.400 1.000 ;
  LAYER VI3 ;
  RECT 1425.600 0.200 1426.400 1.000 ;
  LAYER VI1 ;
  RECT 1410.800 0.200 1411.600 1.000 ;
  LAYER VI2 ;
  RECT 1410.800 0.200 1411.600 1.000 ;
  LAYER VI3 ;
  RECT 1410.800 0.200 1411.600 1.000 ;
  LAYER VI1 ;
  RECT 1404.400 0.200 1405.200 1.000 ;
  LAYER VI2 ;
  RECT 1404.400 0.200 1405.200 1.000 ;
  LAYER VI3 ;
  RECT 1404.400 0.200 1405.200 1.000 ;
  LAYER VI1 ;
  RECT 1390.000 0.200 1390.800 1.000 ;
  LAYER VI2 ;
  RECT 1390.000 0.200 1390.800 1.000 ;
  LAYER VI3 ;
  RECT 1390.000 0.200 1390.800 1.000 ;
  LAYER VI1 ;
  RECT 1384.800 0.200 1385.600 1.000 ;
  LAYER VI2 ;
  RECT 1384.800 0.200 1385.600 1.000 ;
  LAYER VI3 ;
  RECT 1384.800 0.200 1385.600 1.000 ;
  LAYER VI1 ;
  RECT 1371.600 0.200 1372.400 1.000 ;
  LAYER VI2 ;
  RECT 1371.600 0.200 1372.400 1.000 ;
  LAYER VI3 ;
  RECT 1371.600 0.200 1372.400 1.000 ;
  LAYER VI1 ;
  RECT 1370.000 0.200 1370.800 1.000 ;
  LAYER VI2 ;
  RECT 1370.000 0.200 1370.800 1.000 ;
  LAYER VI3 ;
  RECT 1370.000 0.200 1370.800 1.000 ;
  LAYER VI1 ;
  RECT 1349.200 0.200 1350.000 1.000 ;
  LAYER VI2 ;
  RECT 1349.200 0.200 1350.000 1.000 ;
  LAYER VI3 ;
  RECT 1349.200 0.200 1350.000 1.000 ;
  LAYER VI1 ;
  RECT 1348.000 0.200 1348.800 1.000 ;
  LAYER VI2 ;
  RECT 1348.000 0.200 1348.800 1.000 ;
  LAYER VI3 ;
  RECT 1348.000 0.200 1348.800 1.000 ;
  LAYER VI1 ;
  RECT 1346.800 0.200 1347.600 1.000 ;
  LAYER VI2 ;
  RECT 1346.800 0.200 1347.600 1.000 ;
  LAYER VI3 ;
  RECT 1346.800 0.200 1347.600 1.000 ;
  LAYER VI1 ;
  RECT 1345.600 0.200 1346.400 1.000 ;
  LAYER VI2 ;
  RECT 1345.600 0.200 1346.400 1.000 ;
  LAYER VI3 ;
  RECT 1345.600 0.200 1346.400 1.000 ;
  LAYER VI1 ;
  RECT 1344.400 0.200 1345.200 1.000 ;
  LAYER VI2 ;
  RECT 1344.400 0.200 1345.200 1.000 ;
  LAYER VI3 ;
  RECT 1344.400 0.200 1345.200 1.000 ;
  LAYER VI1 ;
  RECT 1343.200 0.200 1344.000 1.000 ;
  LAYER VI2 ;
  RECT 1343.200 0.200 1344.000 1.000 ;
  LAYER VI3 ;
  RECT 1343.200 0.200 1344.000 1.000 ;
  LAYER VI1 ;
  RECT 1337.200 0.200 1338.000 1.000 ;
  LAYER VI2 ;
  RECT 1337.200 0.200 1338.000 1.000 ;
  LAYER VI3 ;
  RECT 1337.200 0.200 1338.000 1.000 ;
  LAYER VI1 ;
  RECT 1330.000 0.200 1330.800 1.000 ;
  LAYER VI2 ;
  RECT 1330.000 0.200 1330.800 1.000 ;
  LAYER VI3 ;
  RECT 1330.000 0.200 1330.800 1.000 ;
  LAYER VI1 ;
  RECT 1327.200 0.200 1328.000 1.000 ;
  LAYER VI2 ;
  RECT 1327.200 0.200 1328.000 1.000 ;
  LAYER VI3 ;
  RECT 1327.200 0.200 1328.000 1.000 ;
  LAYER VI1 ;
  RECT 1324.400 0.200 1325.200 1.000 ;
  LAYER VI2 ;
  RECT 1324.400 0.200 1325.200 1.000 ;
  LAYER VI3 ;
  RECT 1324.400 0.200 1325.200 1.000 ;
  LAYER VI1 ;
  RECT 1322.000 0.200 1322.800 1.000 ;
  LAYER VI2 ;
  RECT 1322.000 0.200 1322.800 1.000 ;
  LAYER VI3 ;
  RECT 1322.000 0.200 1322.800 1.000 ;
  LAYER VI1 ;
  RECT 1320.400 0.200 1321.200 1.000 ;
  LAYER VI2 ;
  RECT 1320.400 0.200 1321.200 1.000 ;
  LAYER VI3 ;
  RECT 1320.400 0.200 1321.200 1.000 ;
  LAYER VI1 ;
  RECT 1318.000 0.200 1318.800 1.000 ;
  LAYER VI2 ;
  RECT 1318.000 0.200 1318.800 1.000 ;
  LAYER VI3 ;
  RECT 1318.000 0.200 1318.800 1.000 ;
  LAYER VI1 ;
  RECT 1311.200 0.200 1312.000 1.000 ;
  LAYER VI2 ;
  RECT 1311.200 0.200 1312.000 1.000 ;
  LAYER VI3 ;
  RECT 1311.200 0.200 1312.000 1.000 ;
  LAYER VI1 ;
  RECT 1296.400 0.200 1297.200 1.000 ;
  LAYER VI2 ;
  RECT 1296.400 0.200 1297.200 1.000 ;
  LAYER VI3 ;
  RECT 1296.400 0.200 1297.200 1.000 ;
  LAYER VI1 ;
  RECT 1291.200 0.200 1292.000 1.000 ;
  LAYER VI2 ;
  RECT 1291.200 0.200 1292.000 1.000 ;
  LAYER VI3 ;
  RECT 1291.200 0.200 1292.000 1.000 ;
  LAYER VI1 ;
  RECT 1276.800 0.200 1277.600 1.000 ;
  LAYER VI2 ;
  RECT 1276.800 0.200 1277.600 1.000 ;
  LAYER VI3 ;
  RECT 1276.800 0.200 1277.600 1.000 ;
  LAYER VI1 ;
  RECT 1270.400 0.200 1271.200 1.000 ;
  LAYER VI2 ;
  RECT 1270.400 0.200 1271.200 1.000 ;
  LAYER VI3 ;
  RECT 1270.400 0.200 1271.200 1.000 ;
  LAYER VI1 ;
  RECT 1255.600 0.200 1256.400 1.000 ;
  LAYER VI2 ;
  RECT 1255.600 0.200 1256.400 1.000 ;
  LAYER VI3 ;
  RECT 1255.600 0.200 1256.400 1.000 ;
  LAYER VI1 ;
  RECT 1250.400 0.200 1251.200 1.000 ;
  LAYER VI2 ;
  RECT 1250.400 0.200 1251.200 1.000 ;
  LAYER VI3 ;
  RECT 1250.400 0.200 1251.200 1.000 ;
  LAYER VI1 ;
  RECT 1235.600 0.200 1236.400 1.000 ;
  LAYER VI2 ;
  RECT 1235.600 0.200 1236.400 1.000 ;
  LAYER VI3 ;
  RECT 1235.600 0.200 1236.400 1.000 ;
  LAYER VI1 ;
  RECT 1229.200 0.200 1230.000 1.000 ;
  LAYER VI2 ;
  RECT 1229.200 0.200 1230.000 1.000 ;
  LAYER VI3 ;
  RECT 1229.200 0.200 1230.000 1.000 ;
  LAYER VI1 ;
  RECT 1214.800 0.200 1215.600 1.000 ;
  LAYER VI2 ;
  RECT 1214.800 0.200 1215.600 1.000 ;
  LAYER VI3 ;
  RECT 1214.800 0.200 1215.600 1.000 ;
  LAYER VI1 ;
  RECT 1209.600 0.200 1210.400 1.000 ;
  LAYER VI2 ;
  RECT 1209.600 0.200 1210.400 1.000 ;
  LAYER VI3 ;
  RECT 1209.600 0.200 1210.400 1.000 ;
  LAYER VI1 ;
  RECT 1194.800 0.200 1195.600 1.000 ;
  LAYER VI2 ;
  RECT 1194.800 0.200 1195.600 1.000 ;
  LAYER VI3 ;
  RECT 1194.800 0.200 1195.600 1.000 ;
  LAYER VI1 ;
  RECT 1188.400 0.200 1189.200 1.000 ;
  LAYER VI2 ;
  RECT 1188.400 0.200 1189.200 1.000 ;
  LAYER VI3 ;
  RECT 1188.400 0.200 1189.200 1.000 ;
  LAYER VI1 ;
  RECT 1173.600 0.200 1174.400 1.000 ;
  LAYER VI2 ;
  RECT 1173.600 0.200 1174.400 1.000 ;
  LAYER VI3 ;
  RECT 1173.600 0.200 1174.400 1.000 ;
  LAYER VI1 ;
  RECT 1168.400 0.200 1169.200 1.000 ;
  LAYER VI2 ;
  RECT 1168.400 0.200 1169.200 1.000 ;
  LAYER VI3 ;
  RECT 1168.400 0.200 1169.200 1.000 ;
  LAYER VI1 ;
  RECT 1154.000 0.200 1154.800 1.000 ;
  LAYER VI2 ;
  RECT 1154.000 0.200 1154.800 1.000 ;
  LAYER VI3 ;
  RECT 1154.000 0.200 1154.800 1.000 ;
  LAYER VI1 ;
  RECT 1147.600 0.200 1148.400 1.000 ;
  LAYER VI2 ;
  RECT 1147.600 0.200 1148.400 1.000 ;
  LAYER VI3 ;
  RECT 1147.600 0.200 1148.400 1.000 ;
  LAYER VI1 ;
  RECT 1132.800 0.200 1133.600 1.000 ;
  LAYER VI2 ;
  RECT 1132.800 0.200 1133.600 1.000 ;
  LAYER VI3 ;
  RECT 1132.800 0.200 1133.600 1.000 ;
  LAYER VI1 ;
  RECT 1127.600 0.200 1128.400 1.000 ;
  LAYER VI2 ;
  RECT 1127.600 0.200 1128.400 1.000 ;
  LAYER VI3 ;
  RECT 1127.600 0.200 1128.400 1.000 ;
  LAYER VI1 ;
  RECT 1113.200 0.200 1114.000 1.000 ;
  LAYER VI2 ;
  RECT 1113.200 0.200 1114.000 1.000 ;
  LAYER VI3 ;
  RECT 1113.200 0.200 1114.000 1.000 ;
  LAYER VI1 ;
  RECT 1106.400 0.200 1107.200 1.000 ;
  LAYER VI2 ;
  RECT 1106.400 0.200 1107.200 1.000 ;
  LAYER VI3 ;
  RECT 1106.400 0.200 1107.200 1.000 ;
  LAYER VI1 ;
  RECT 1092.000 0.200 1092.800 1.000 ;
  LAYER VI2 ;
  RECT 1092.000 0.200 1092.800 1.000 ;
  LAYER VI3 ;
  RECT 1092.000 0.200 1092.800 1.000 ;
  LAYER VI1 ;
  RECT 1086.800 0.200 1087.600 1.000 ;
  LAYER VI2 ;
  RECT 1086.800 0.200 1087.600 1.000 ;
  LAYER VI3 ;
  RECT 1086.800 0.200 1087.600 1.000 ;
  LAYER VI1 ;
  RECT 1072.000 0.200 1072.800 1.000 ;
  LAYER VI2 ;
  RECT 1072.000 0.200 1072.800 1.000 ;
  LAYER VI3 ;
  RECT 1072.000 0.200 1072.800 1.000 ;
  LAYER VI1 ;
  RECT 1065.600 0.200 1066.400 1.000 ;
  LAYER VI2 ;
  RECT 1065.600 0.200 1066.400 1.000 ;
  LAYER VI3 ;
  RECT 1065.600 0.200 1066.400 1.000 ;
  LAYER VI1 ;
  RECT 1051.200 0.200 1052.000 1.000 ;
  LAYER VI2 ;
  RECT 1051.200 0.200 1052.000 1.000 ;
  LAYER VI3 ;
  RECT 1051.200 0.200 1052.000 1.000 ;
  LAYER VI1 ;
  RECT 1045.600 0.200 1046.400 1.000 ;
  LAYER VI2 ;
  RECT 1045.600 0.200 1046.400 1.000 ;
  LAYER VI3 ;
  RECT 1045.600 0.200 1046.400 1.000 ;
  LAYER VI1 ;
  RECT 1031.200 0.200 1032.000 1.000 ;
  LAYER VI2 ;
  RECT 1031.200 0.200 1032.000 1.000 ;
  LAYER VI3 ;
  RECT 1031.200 0.200 1032.000 1.000 ;
  LAYER VI1 ;
  RECT 1024.800 0.200 1025.600 1.000 ;
  LAYER VI2 ;
  RECT 1024.800 0.200 1025.600 1.000 ;
  LAYER VI3 ;
  RECT 1024.800 0.200 1025.600 1.000 ;
  LAYER VI1 ;
  RECT 1010.000 0.200 1010.800 1.000 ;
  LAYER VI2 ;
  RECT 1010.000 0.200 1010.800 1.000 ;
  LAYER VI3 ;
  RECT 1010.000 0.200 1010.800 1.000 ;
  LAYER VI1 ;
  RECT 1004.800 0.200 1005.600 1.000 ;
  LAYER VI2 ;
  RECT 1004.800 0.200 1005.600 1.000 ;
  LAYER VI3 ;
  RECT 1004.800 0.200 1005.600 1.000 ;
  LAYER VI1 ;
  RECT 992.000 0.200 992.800 1.000 ;
  LAYER VI2 ;
  RECT 992.000 0.200 992.800 1.000 ;
  LAYER VI3 ;
  RECT 992.000 0.200 992.800 1.000 ;
  LAYER VI1 ;
  RECT 990.400 0.200 991.200 1.000 ;
  LAYER VI2 ;
  RECT 990.400 0.200 991.200 1.000 ;
  LAYER VI3 ;
  RECT 990.400 0.200 991.200 1.000 ;
  LAYER VI1 ;
  RECT 983.600 0.200 984.400 1.000 ;
  LAYER VI2 ;
  RECT 983.600 0.200 984.400 1.000 ;
  LAYER VI3 ;
  RECT 983.600 0.200 984.400 1.000 ;
  LAYER VI1 ;
  RECT 969.200 0.200 970.000 1.000 ;
  LAYER VI2 ;
  RECT 969.200 0.200 970.000 1.000 ;
  LAYER VI3 ;
  RECT 969.200 0.200 970.000 1.000 ;
  LAYER VI1 ;
  RECT 964.000 0.200 964.800 1.000 ;
  LAYER VI2 ;
  RECT 964.000 0.200 964.800 1.000 ;
  LAYER VI3 ;
  RECT 964.000 0.200 964.800 1.000 ;
  LAYER VI1 ;
  RECT 949.200 0.200 950.000 1.000 ;
  LAYER VI2 ;
  RECT 949.200 0.200 950.000 1.000 ;
  LAYER VI3 ;
  RECT 949.200 0.200 950.000 1.000 ;
  LAYER VI1 ;
  RECT 942.800 0.200 943.600 1.000 ;
  LAYER VI2 ;
  RECT 942.800 0.200 943.600 1.000 ;
  LAYER VI3 ;
  RECT 942.800 0.200 943.600 1.000 ;
  LAYER VI1 ;
  RECT 928.400 0.200 929.200 1.000 ;
  LAYER VI2 ;
  RECT 928.400 0.200 929.200 1.000 ;
  LAYER VI3 ;
  RECT 928.400 0.200 929.200 1.000 ;
  LAYER VI1 ;
  RECT 923.200 0.200 924.000 1.000 ;
  LAYER VI2 ;
  RECT 923.200 0.200 924.000 1.000 ;
  LAYER VI3 ;
  RECT 923.200 0.200 924.000 1.000 ;
  LAYER VI1 ;
  RECT 908.400 0.200 909.200 1.000 ;
  LAYER VI2 ;
  RECT 908.400 0.200 909.200 1.000 ;
  LAYER VI3 ;
  RECT 908.400 0.200 909.200 1.000 ;
  LAYER VI1 ;
  RECT 902.000 0.200 902.800 1.000 ;
  LAYER VI2 ;
  RECT 902.000 0.200 902.800 1.000 ;
  LAYER VI3 ;
  RECT 902.000 0.200 902.800 1.000 ;
  LAYER VI1 ;
  RECT 887.200 0.200 888.000 1.000 ;
  LAYER VI2 ;
  RECT 887.200 0.200 888.000 1.000 ;
  LAYER VI3 ;
  RECT 887.200 0.200 888.000 1.000 ;
  LAYER VI1 ;
  RECT 882.000 0.200 882.800 1.000 ;
  LAYER VI2 ;
  RECT 882.000 0.200 882.800 1.000 ;
  LAYER VI3 ;
  RECT 882.000 0.200 882.800 1.000 ;
  LAYER VI1 ;
  RECT 867.600 0.200 868.400 1.000 ;
  LAYER VI2 ;
  RECT 867.600 0.200 868.400 1.000 ;
  LAYER VI3 ;
  RECT 867.600 0.200 868.400 1.000 ;
  LAYER VI1 ;
  RECT 861.200 0.200 862.000 1.000 ;
  LAYER VI2 ;
  RECT 861.200 0.200 862.000 1.000 ;
  LAYER VI3 ;
  RECT 861.200 0.200 862.000 1.000 ;
  LAYER VI1 ;
  RECT 846.400 0.200 847.200 1.000 ;
  LAYER VI2 ;
  RECT 846.400 0.200 847.200 1.000 ;
  LAYER VI3 ;
  RECT 846.400 0.200 847.200 1.000 ;
  LAYER VI1 ;
  RECT 841.200 0.200 842.000 1.000 ;
  LAYER VI2 ;
  RECT 841.200 0.200 842.000 1.000 ;
  LAYER VI3 ;
  RECT 841.200 0.200 842.000 1.000 ;
  LAYER VI1 ;
  RECT 826.400 0.200 827.200 1.000 ;
  LAYER VI2 ;
  RECT 826.400 0.200 827.200 1.000 ;
  LAYER VI3 ;
  RECT 826.400 0.200 827.200 1.000 ;
  LAYER VI1 ;
  RECT 820.000 0.200 820.800 1.000 ;
  LAYER VI2 ;
  RECT 820.000 0.200 820.800 1.000 ;
  LAYER VI3 ;
  RECT 820.000 0.200 820.800 1.000 ;
  LAYER VI1 ;
  RECT 805.600 0.200 806.400 1.000 ;
  LAYER VI2 ;
  RECT 805.600 0.200 806.400 1.000 ;
  LAYER VI3 ;
  RECT 805.600 0.200 806.400 1.000 ;
  LAYER VI1 ;
  RECT 800.400 0.200 801.200 1.000 ;
  LAYER VI2 ;
  RECT 800.400 0.200 801.200 1.000 ;
  LAYER VI3 ;
  RECT 800.400 0.200 801.200 1.000 ;
  LAYER VI1 ;
  RECT 785.600 0.200 786.400 1.000 ;
  LAYER VI2 ;
  RECT 785.600 0.200 786.400 1.000 ;
  LAYER VI3 ;
  RECT 785.600 0.200 786.400 1.000 ;
  LAYER VI1 ;
  RECT 779.200 0.200 780.000 1.000 ;
  LAYER VI2 ;
  RECT 779.200 0.200 780.000 1.000 ;
  LAYER VI3 ;
  RECT 779.200 0.200 780.000 1.000 ;
  LAYER VI1 ;
  RECT 764.400 0.200 765.200 1.000 ;
  LAYER VI2 ;
  RECT 764.400 0.200 765.200 1.000 ;
  LAYER VI3 ;
  RECT 764.400 0.200 765.200 1.000 ;
  LAYER VI1 ;
  RECT 759.200 0.200 760.000 1.000 ;
  LAYER VI2 ;
  RECT 759.200 0.200 760.000 1.000 ;
  LAYER VI3 ;
  RECT 759.200 0.200 760.000 1.000 ;
  LAYER VI1 ;
  RECT 744.800 0.200 745.600 1.000 ;
  LAYER VI2 ;
  RECT 744.800 0.200 745.600 1.000 ;
  LAYER VI3 ;
  RECT 744.800 0.200 745.600 1.000 ;
  LAYER VI1 ;
  RECT 738.400 0.200 739.200 1.000 ;
  LAYER VI2 ;
  RECT 738.400 0.200 739.200 1.000 ;
  LAYER VI3 ;
  RECT 738.400 0.200 739.200 1.000 ;
  LAYER VI1 ;
  RECT 723.600 0.200 724.400 1.000 ;
  LAYER VI2 ;
  RECT 723.600 0.200 724.400 1.000 ;
  LAYER VI3 ;
  RECT 723.600 0.200 724.400 1.000 ;
  LAYER VI1 ;
  RECT 718.400 0.200 719.200 1.000 ;
  LAYER VI2 ;
  RECT 718.400 0.200 719.200 1.000 ;
  LAYER VI3 ;
  RECT 718.400 0.200 719.200 1.000 ;
  LAYER VI1 ;
  RECT 704.000 0.200 704.800 1.000 ;
  LAYER VI2 ;
  RECT 704.000 0.200 704.800 1.000 ;
  LAYER VI3 ;
  RECT 704.000 0.200 704.800 1.000 ;
  LAYER VI1 ;
  RECT 697.200 0.200 698.000 1.000 ;
  LAYER VI2 ;
  RECT 697.200 0.200 698.000 1.000 ;
  LAYER VI3 ;
  RECT 697.200 0.200 698.000 1.000 ;
  LAYER VI1 ;
  RECT 682.800 0.200 683.600 1.000 ;
  LAYER VI2 ;
  RECT 682.800 0.200 683.600 1.000 ;
  LAYER VI3 ;
  RECT 682.800 0.200 683.600 1.000 ;
  LAYER VI1 ;
  RECT 677.600 0.200 678.400 1.000 ;
  LAYER VI2 ;
  RECT 677.600 0.200 678.400 1.000 ;
  LAYER VI3 ;
  RECT 677.600 0.200 678.400 1.000 ;
  LAYER VI1 ;
  RECT 664.800 0.200 665.600 1.000 ;
  LAYER VI2 ;
  RECT 664.800 0.200 665.600 1.000 ;
  LAYER VI3 ;
  RECT 664.800 0.200 665.600 1.000 ;
  LAYER VI1 ;
  RECT 662.800 0.200 663.600 1.000 ;
  LAYER VI2 ;
  RECT 662.800 0.200 663.600 1.000 ;
  LAYER VI3 ;
  RECT 662.800 0.200 663.600 1.000 ;
  LAYER VI1 ;
  RECT 656.400 0.200 657.200 1.000 ;
  LAYER VI2 ;
  RECT 656.400 0.200 657.200 1.000 ;
  LAYER VI3 ;
  RECT 656.400 0.200 657.200 1.000 ;
  LAYER VI1 ;
  RECT 642.000 0.200 642.800 1.000 ;
  LAYER VI2 ;
  RECT 642.000 0.200 642.800 1.000 ;
  LAYER VI3 ;
  RECT 642.000 0.200 642.800 1.000 ;
  LAYER VI1 ;
  RECT 636.400 0.200 637.200 1.000 ;
  LAYER VI2 ;
  RECT 636.400 0.200 637.200 1.000 ;
  LAYER VI3 ;
  RECT 636.400 0.200 637.200 1.000 ;
  LAYER VI1 ;
  RECT 622.000 0.200 622.800 1.000 ;
  LAYER VI2 ;
  RECT 622.000 0.200 622.800 1.000 ;
  LAYER VI3 ;
  RECT 622.000 0.200 622.800 1.000 ;
  LAYER VI1 ;
  RECT 615.600 0.200 616.400 1.000 ;
  LAYER VI2 ;
  RECT 615.600 0.200 616.400 1.000 ;
  LAYER VI3 ;
  RECT 615.600 0.200 616.400 1.000 ;
  LAYER VI1 ;
  RECT 600.800 0.200 601.600 1.000 ;
  LAYER VI2 ;
  RECT 600.800 0.200 601.600 1.000 ;
  LAYER VI3 ;
  RECT 600.800 0.200 601.600 1.000 ;
  LAYER VI1 ;
  RECT 595.600 0.200 596.400 1.000 ;
  LAYER VI2 ;
  RECT 595.600 0.200 596.400 1.000 ;
  LAYER VI3 ;
  RECT 595.600 0.200 596.400 1.000 ;
  LAYER VI1 ;
  RECT 581.200 0.200 582.000 1.000 ;
  LAYER VI2 ;
  RECT 581.200 0.200 582.000 1.000 ;
  LAYER VI3 ;
  RECT 581.200 0.200 582.000 1.000 ;
  LAYER VI1 ;
  RECT 574.400 0.200 575.200 1.000 ;
  LAYER VI2 ;
  RECT 574.400 0.200 575.200 1.000 ;
  LAYER VI3 ;
  RECT 574.400 0.200 575.200 1.000 ;
  LAYER VI1 ;
  RECT 560.000 0.200 560.800 1.000 ;
  LAYER VI2 ;
  RECT 560.000 0.200 560.800 1.000 ;
  LAYER VI3 ;
  RECT 560.000 0.200 560.800 1.000 ;
  LAYER VI1 ;
  RECT 554.800 0.200 555.600 1.000 ;
  LAYER VI2 ;
  RECT 554.800 0.200 555.600 1.000 ;
  LAYER VI3 ;
  RECT 554.800 0.200 555.600 1.000 ;
  LAYER VI1 ;
  RECT 540.000 0.200 540.800 1.000 ;
  LAYER VI2 ;
  RECT 540.000 0.200 540.800 1.000 ;
  LAYER VI3 ;
  RECT 540.000 0.200 540.800 1.000 ;
  LAYER VI1 ;
  RECT 533.600 0.200 534.400 1.000 ;
  LAYER VI2 ;
  RECT 533.600 0.200 534.400 1.000 ;
  LAYER VI3 ;
  RECT 533.600 0.200 534.400 1.000 ;
  LAYER VI1 ;
  RECT 519.200 0.200 520.000 1.000 ;
  LAYER VI2 ;
  RECT 519.200 0.200 520.000 1.000 ;
  LAYER VI3 ;
  RECT 519.200 0.200 520.000 1.000 ;
  LAYER VI1 ;
  RECT 514.000 0.200 514.800 1.000 ;
  LAYER VI2 ;
  RECT 514.000 0.200 514.800 1.000 ;
  LAYER VI3 ;
  RECT 514.000 0.200 514.800 1.000 ;
  LAYER VI1 ;
  RECT 499.200 0.200 500.000 1.000 ;
  LAYER VI2 ;
  RECT 499.200 0.200 500.000 1.000 ;
  LAYER VI3 ;
  RECT 499.200 0.200 500.000 1.000 ;
  LAYER VI1 ;
  RECT 492.800 0.200 493.600 1.000 ;
  LAYER VI2 ;
  RECT 492.800 0.200 493.600 1.000 ;
  LAYER VI3 ;
  RECT 492.800 0.200 493.600 1.000 ;
  LAYER VI1 ;
  RECT 478.000 0.200 478.800 1.000 ;
  LAYER VI2 ;
  RECT 478.000 0.200 478.800 1.000 ;
  LAYER VI3 ;
  RECT 478.000 0.200 478.800 1.000 ;
  LAYER VI1 ;
  RECT 472.800 0.200 473.600 1.000 ;
  LAYER VI2 ;
  RECT 472.800 0.200 473.600 1.000 ;
  LAYER VI3 ;
  RECT 472.800 0.200 473.600 1.000 ;
  LAYER VI1 ;
  RECT 458.400 0.200 459.200 1.000 ;
  LAYER VI2 ;
  RECT 458.400 0.200 459.200 1.000 ;
  LAYER VI3 ;
  RECT 458.400 0.200 459.200 1.000 ;
  LAYER VI1 ;
  RECT 452.000 0.200 452.800 1.000 ;
  LAYER VI2 ;
  RECT 452.000 0.200 452.800 1.000 ;
  LAYER VI3 ;
  RECT 452.000 0.200 452.800 1.000 ;
  LAYER VI1 ;
  RECT 437.200 0.200 438.000 1.000 ;
  LAYER VI2 ;
  RECT 437.200 0.200 438.000 1.000 ;
  LAYER VI3 ;
  RECT 437.200 0.200 438.000 1.000 ;
  LAYER VI1 ;
  RECT 432.000 0.200 432.800 1.000 ;
  LAYER VI2 ;
  RECT 432.000 0.200 432.800 1.000 ;
  LAYER VI3 ;
  RECT 432.000 0.200 432.800 1.000 ;
  LAYER VI1 ;
  RECT 417.200 0.200 418.000 1.000 ;
  LAYER VI2 ;
  RECT 417.200 0.200 418.000 1.000 ;
  LAYER VI3 ;
  RECT 417.200 0.200 418.000 1.000 ;
  LAYER VI1 ;
  RECT 410.800 0.200 411.600 1.000 ;
  LAYER VI2 ;
  RECT 410.800 0.200 411.600 1.000 ;
  LAYER VI3 ;
  RECT 410.800 0.200 411.600 1.000 ;
  LAYER VI1 ;
  RECT 396.400 0.200 397.200 1.000 ;
  LAYER VI2 ;
  RECT 396.400 0.200 397.200 1.000 ;
  LAYER VI3 ;
  RECT 396.400 0.200 397.200 1.000 ;
  LAYER VI1 ;
  RECT 391.200 0.200 392.000 1.000 ;
  LAYER VI2 ;
  RECT 391.200 0.200 392.000 1.000 ;
  LAYER VI3 ;
  RECT 391.200 0.200 392.000 1.000 ;
  LAYER VI1 ;
  RECT 376.400 0.200 377.200 1.000 ;
  LAYER VI2 ;
  RECT 376.400 0.200 377.200 1.000 ;
  LAYER VI3 ;
  RECT 376.400 0.200 377.200 1.000 ;
  LAYER VI1 ;
  RECT 370.000 0.200 370.800 1.000 ;
  LAYER VI2 ;
  RECT 370.000 0.200 370.800 1.000 ;
  LAYER VI3 ;
  RECT 370.000 0.200 370.800 1.000 ;
  LAYER VI1 ;
  RECT 355.200 0.200 356.000 1.000 ;
  LAYER VI2 ;
  RECT 355.200 0.200 356.000 1.000 ;
  LAYER VI3 ;
  RECT 355.200 0.200 356.000 1.000 ;
  LAYER VI1 ;
  RECT 350.000 0.200 350.800 1.000 ;
  LAYER VI2 ;
  RECT 350.000 0.200 350.800 1.000 ;
  LAYER VI3 ;
  RECT 350.000 0.200 350.800 1.000 ;
  LAYER VI1 ;
  RECT 337.200 0.200 338.000 1.000 ;
  LAYER VI2 ;
  RECT 337.200 0.200 338.000 1.000 ;
  LAYER VI3 ;
  RECT 337.200 0.200 338.000 1.000 ;
  LAYER VI1 ;
  RECT 335.600 0.200 336.400 1.000 ;
  LAYER VI2 ;
  RECT 335.600 0.200 336.400 1.000 ;
  LAYER VI3 ;
  RECT 335.600 0.200 336.400 1.000 ;
  LAYER VI1 ;
  RECT 329.200 0.200 330.000 1.000 ;
  LAYER VI2 ;
  RECT 329.200 0.200 330.000 1.000 ;
  LAYER VI3 ;
  RECT 329.200 0.200 330.000 1.000 ;
  LAYER VI1 ;
  RECT 314.400 0.200 315.200 1.000 ;
  LAYER VI2 ;
  RECT 314.400 0.200 315.200 1.000 ;
  LAYER VI3 ;
  RECT 314.400 0.200 315.200 1.000 ;
  LAYER VI1 ;
  RECT 309.200 0.200 310.000 1.000 ;
  LAYER VI2 ;
  RECT 309.200 0.200 310.000 1.000 ;
  LAYER VI3 ;
  RECT 309.200 0.200 310.000 1.000 ;
  LAYER VI1 ;
  RECT 294.800 0.200 295.600 1.000 ;
  LAYER VI2 ;
  RECT 294.800 0.200 295.600 1.000 ;
  LAYER VI3 ;
  RECT 294.800 0.200 295.600 1.000 ;
  LAYER VI1 ;
  RECT 288.000 0.200 288.800 1.000 ;
  LAYER VI2 ;
  RECT 288.000 0.200 288.800 1.000 ;
  LAYER VI3 ;
  RECT 288.000 0.200 288.800 1.000 ;
  LAYER VI1 ;
  RECT 273.600 0.200 274.400 1.000 ;
  LAYER VI2 ;
  RECT 273.600 0.200 274.400 1.000 ;
  LAYER VI3 ;
  RECT 273.600 0.200 274.400 1.000 ;
  LAYER VI1 ;
  RECT 268.400 0.200 269.200 1.000 ;
  LAYER VI2 ;
  RECT 268.400 0.200 269.200 1.000 ;
  LAYER VI3 ;
  RECT 268.400 0.200 269.200 1.000 ;
  LAYER VI1 ;
  RECT 253.600 0.200 254.400 1.000 ;
  LAYER VI2 ;
  RECT 253.600 0.200 254.400 1.000 ;
  LAYER VI3 ;
  RECT 253.600 0.200 254.400 1.000 ;
  LAYER VI1 ;
  RECT 247.200 0.200 248.000 1.000 ;
  LAYER VI2 ;
  RECT 247.200 0.200 248.000 1.000 ;
  LAYER VI3 ;
  RECT 247.200 0.200 248.000 1.000 ;
  LAYER VI1 ;
  RECT 232.800 0.200 233.600 1.000 ;
  LAYER VI2 ;
  RECT 232.800 0.200 233.600 1.000 ;
  LAYER VI3 ;
  RECT 232.800 0.200 233.600 1.000 ;
  LAYER VI1 ;
  RECT 227.200 0.200 228.000 1.000 ;
  LAYER VI2 ;
  RECT 227.200 0.200 228.000 1.000 ;
  LAYER VI3 ;
  RECT 227.200 0.200 228.000 1.000 ;
  LAYER VI1 ;
  RECT 212.800 0.200 213.600 1.000 ;
  LAYER VI2 ;
  RECT 212.800 0.200 213.600 1.000 ;
  LAYER VI3 ;
  RECT 212.800 0.200 213.600 1.000 ;
  LAYER VI1 ;
  RECT 206.400 0.200 207.200 1.000 ;
  LAYER VI2 ;
  RECT 206.400 0.200 207.200 1.000 ;
  LAYER VI3 ;
  RECT 206.400 0.200 207.200 1.000 ;
  LAYER VI1 ;
  RECT 191.600 0.200 192.400 1.000 ;
  LAYER VI2 ;
  RECT 191.600 0.200 192.400 1.000 ;
  LAYER VI3 ;
  RECT 191.600 0.200 192.400 1.000 ;
  LAYER VI1 ;
  RECT 186.400 0.200 187.200 1.000 ;
  LAYER VI2 ;
  RECT 186.400 0.200 187.200 1.000 ;
  LAYER VI3 ;
  RECT 186.400 0.200 187.200 1.000 ;
  LAYER VI1 ;
  RECT 172.000 0.200 172.800 1.000 ;
  LAYER VI2 ;
  RECT 172.000 0.200 172.800 1.000 ;
  LAYER VI3 ;
  RECT 172.000 0.200 172.800 1.000 ;
  LAYER VI1 ;
  RECT 165.200 0.200 166.000 1.000 ;
  LAYER VI2 ;
  RECT 165.200 0.200 166.000 1.000 ;
  LAYER VI3 ;
  RECT 165.200 0.200 166.000 1.000 ;
  LAYER VI1 ;
  RECT 150.800 0.200 151.600 1.000 ;
  LAYER VI2 ;
  RECT 150.800 0.200 151.600 1.000 ;
  LAYER VI3 ;
  RECT 150.800 0.200 151.600 1.000 ;
  LAYER VI1 ;
  RECT 145.600 0.200 146.400 1.000 ;
  LAYER VI2 ;
  RECT 145.600 0.200 146.400 1.000 ;
  LAYER VI3 ;
  RECT 145.600 0.200 146.400 1.000 ;
  LAYER VI1 ;
  RECT 130.800 0.200 131.600 1.000 ;
  LAYER VI2 ;
  RECT 130.800 0.200 131.600 1.000 ;
  LAYER VI3 ;
  RECT 130.800 0.200 131.600 1.000 ;
  LAYER VI1 ;
  RECT 124.400 0.200 125.200 1.000 ;
  LAYER VI2 ;
  RECT 124.400 0.200 125.200 1.000 ;
  LAYER VI3 ;
  RECT 124.400 0.200 125.200 1.000 ;
  LAYER VI1 ;
  RECT 110.000 0.200 110.800 1.000 ;
  LAYER VI2 ;
  RECT 110.000 0.200 110.800 1.000 ;
  LAYER VI3 ;
  RECT 110.000 0.200 110.800 1.000 ;
  LAYER VI1 ;
  RECT 104.800 0.200 105.600 1.000 ;
  LAYER VI2 ;
  RECT 104.800 0.200 105.600 1.000 ;
  LAYER VI3 ;
  RECT 104.800 0.200 105.600 1.000 ;
  LAYER VI1 ;
  RECT 90.000 0.200 90.800 1.000 ;
  LAYER VI2 ;
  RECT 90.000 0.200 90.800 1.000 ;
  LAYER VI3 ;
  RECT 90.000 0.200 90.800 1.000 ;
  LAYER VI1 ;
  RECT 83.600 0.200 84.400 1.000 ;
  LAYER VI2 ;
  RECT 83.600 0.200 84.400 1.000 ;
  LAYER VI3 ;
  RECT 83.600 0.200 84.400 1.000 ;
  LAYER VI1 ;
  RECT 68.800 0.200 69.600 1.000 ;
  LAYER VI2 ;
  RECT 68.800 0.200 69.600 1.000 ;
  LAYER VI3 ;
  RECT 68.800 0.200 69.600 1.000 ;
  LAYER VI1 ;
  RECT 63.600 0.200 64.400 1.000 ;
  LAYER VI2 ;
  RECT 63.600 0.200 64.400 1.000 ;
  LAYER VI3 ;
  RECT 63.600 0.200 64.400 1.000 ;
  LAYER VI1 ;
  RECT 49.200 0.200 50.000 1.000 ;
  LAYER VI2 ;
  RECT 49.200 0.200 50.000 1.000 ;
  LAYER VI3 ;
  RECT 49.200 0.200 50.000 1.000 ;
  LAYER VI1 ;
  RECT 42.800 0.200 43.600 1.000 ;
  LAYER VI2 ;
  RECT 42.800 0.200 43.600 1.000 ;
  LAYER VI3 ;
  RECT 42.800 0.200 43.600 1.000 ;
  LAYER VI1 ;
  RECT 28.000 0.200 28.800 1.000 ;
  LAYER VI2 ;
  RECT 28.000 0.200 28.800 1.000 ;
  LAYER VI3 ;
  RECT 28.000 0.200 28.800 1.000 ;
  LAYER VI1 ;
  RECT 22.800 0.200 23.600 1.000 ;
  LAYER VI2 ;
  RECT 22.800 0.200 23.600 1.000 ;
  LAYER VI3 ;
  RECT 22.800 0.200 23.600 1.000 ;
  LAYER VI1 ;
  RECT 10.000 0.200 10.800 1.000 ;
  LAYER VI2 ;
  RECT 10.000 0.200 10.800 1.000 ;
  LAYER VI3 ;
  RECT 10.000 0.200 10.800 1.000 ;
  LAYER VI1 ;
  RECT 8.000 0.200 8.800 1.000 ;
  LAYER VI2 ;
  RECT 8.000 0.200 8.800 1.000 ;
  LAYER VI3 ;
  RECT 8.000 0.200 8.800 1.000 ;
  LAYER VI3 ;
  RECT 2679.800 9.570 2680.660 11.170 ;
  LAYER VI3 ;
  RECT 2680.260 10.770 2680.460 10.970 ;
  LAYER VI3 ;
  RECT 2680.260 10.370 2680.460 10.570 ;
  LAYER VI3 ;
  RECT 2680.260 9.970 2680.460 10.170 ;
  LAYER VI3 ;
  RECT 2680.260 9.570 2680.460 9.770 ;
  LAYER VI3 ;
  RECT 2679.860 10.770 2680.060 10.970 ;
  LAYER VI3 ;
  RECT 2679.860 10.370 2680.060 10.570 ;
  LAYER VI3 ;
  RECT 2679.860 9.970 2680.060 10.170 ;
  LAYER VI3 ;
  RECT 2679.860 9.570 2680.060 9.770 ;
  LAYER VI2 ;
  RECT 2679.800 9.570 2680.660 11.170 ;
  LAYER VI2 ;
  RECT 2680.260 10.770 2680.460 10.970 ;
  LAYER VI2 ;
  RECT 2680.260 10.370 2680.460 10.570 ;
  LAYER VI2 ;
  RECT 2680.260 9.970 2680.460 10.170 ;
  LAYER VI2 ;
  RECT 2680.260 9.570 2680.460 9.770 ;
  LAYER VI2 ;
  RECT 2679.860 10.770 2680.060 10.970 ;
  LAYER VI2 ;
  RECT 2679.860 10.370 2680.060 10.570 ;
  LAYER VI2 ;
  RECT 2679.860 9.970 2680.060 10.170 ;
  LAYER VI2 ;
  RECT 2679.860 9.570 2680.060 9.770 ;
  LAYER VI3 ;
  RECT 2679.800 14.200 2680.660 15.200 ;
  LAYER VI3 ;
  RECT 2680.260 14.600 2680.460 14.800 ;
  LAYER VI3 ;
  RECT 2680.260 14.200 2680.460 14.400 ;
  LAYER VI3 ;
  RECT 2679.860 14.600 2680.060 14.800 ;
  LAYER VI3 ;
  RECT 2679.860 14.200 2680.060 14.400 ;
  LAYER VI2 ;
  RECT 2679.800 14.200 2680.660 15.200 ;
  LAYER VI2 ;
  RECT 2680.260 14.600 2680.460 14.800 ;
  LAYER VI2 ;
  RECT 2680.260 14.200 2680.460 14.400 ;
  LAYER VI2 ;
  RECT 2679.860 14.600 2680.060 14.800 ;
  LAYER VI2 ;
  RECT 2679.860 14.200 2680.060 14.400 ;
  LAYER VI3 ;
  RECT 2679.800 18.730 2680.660 19.730 ;
  LAYER VI3 ;
  RECT 2680.260 19.130 2680.460 19.330 ;
  LAYER VI3 ;
  RECT 2680.260 18.730 2680.460 18.930 ;
  LAYER VI3 ;
  RECT 2679.860 19.130 2680.060 19.330 ;
  LAYER VI3 ;
  RECT 2679.860 18.730 2680.060 18.930 ;
  LAYER VI2 ;
  RECT 2679.800 18.730 2680.660 19.730 ;
  LAYER VI2 ;
  RECT 2680.260 19.130 2680.460 19.330 ;
  LAYER VI2 ;
  RECT 2680.260 18.730 2680.460 18.930 ;
  LAYER VI2 ;
  RECT 2679.860 19.130 2680.060 19.330 ;
  LAYER VI2 ;
  RECT 2679.860 18.730 2680.060 18.930 ;
  LAYER VI3 ;
  RECT 2679.800 21.230 2680.660 22.070 ;
  LAYER VI3 ;
  RECT 2680.200 21.690 2680.400 21.890 ;
  LAYER VI3 ;
  RECT 2680.200 21.290 2680.400 21.490 ;
  LAYER VI3 ;
  RECT 2679.800 21.690 2680.000 21.890 ;
  LAYER VI3 ;
  RECT 2679.800 21.290 2680.000 21.490 ;
  LAYER VI2 ;
  RECT 2679.800 21.230 2680.660 22.070 ;
  LAYER VI2 ;
  RECT 2680.200 21.690 2680.400 21.890 ;
  LAYER VI2 ;
  RECT 2680.200 21.290 2680.400 21.490 ;
  LAYER VI2 ;
  RECT 2679.800 21.690 2680.000 21.890 ;
  LAYER VI2 ;
  RECT 2679.800 21.290 2680.000 21.490 ;
  LAYER VI3 ;
  RECT 2679.800 24.170 2680.660 25.170 ;
  LAYER VI3 ;
  RECT 2680.260 24.570 2680.460 24.770 ;
  LAYER VI3 ;
  RECT 2680.260 24.170 2680.460 24.370 ;
  LAYER VI3 ;
  RECT 2679.860 24.570 2680.060 24.770 ;
  LAYER VI3 ;
  RECT 2679.860 24.170 2680.060 24.370 ;
  LAYER VI2 ;
  RECT 2679.800 24.170 2680.660 25.170 ;
  LAYER VI2 ;
  RECT 2680.260 24.570 2680.460 24.770 ;
  LAYER VI2 ;
  RECT 2680.260 24.170 2680.460 24.370 ;
  LAYER VI2 ;
  RECT 2679.860 24.570 2680.060 24.770 ;
  LAYER VI2 ;
  RECT 2679.860 24.170 2680.060 24.370 ;
  LAYER VI3 ;
  RECT 2679.800 36.320 2680.660 37.320 ;
  LAYER VI3 ;
  RECT 2680.260 36.720 2680.460 36.920 ;
  LAYER VI3 ;
  RECT 2680.260 36.320 2680.460 36.520 ;
  LAYER VI3 ;
  RECT 2679.860 36.720 2680.060 36.920 ;
  LAYER VI3 ;
  RECT 2679.860 36.320 2680.060 36.520 ;
  LAYER VI2 ;
  RECT 2679.800 36.320 2680.660 37.320 ;
  LAYER VI2 ;
  RECT 2680.260 36.720 2680.460 36.920 ;
  LAYER VI2 ;
  RECT 2680.260 36.320 2680.460 36.520 ;
  LAYER VI2 ;
  RECT 2679.860 36.720 2680.060 36.920 ;
  LAYER VI2 ;
  RECT 2679.860 36.320 2680.060 36.520 ;
  LAYER VI3 ;
  RECT 2679.800 39.480 2680.660 40.080 ;
  LAYER VI3 ;
  RECT 2680.200 39.540 2680.400 39.740 ;
  LAYER VI3 ;
  RECT 2679.800 39.540 2680.000 39.740 ;
  LAYER VI2 ;
  RECT 2679.800 39.480 2680.660 40.080 ;
  LAYER VI2 ;
  RECT 2680.200 39.540 2680.400 39.740 ;
  LAYER VI2 ;
  RECT 2679.800 39.540 2680.000 39.740 ;
  LAYER VI3 ;
  RECT 2679.800 45.560 2680.660 46.160 ;
  LAYER VI3 ;
  RECT 2680.200 45.620 2680.400 45.820 ;
  LAYER VI3 ;
  RECT 2679.800 45.620 2680.000 45.820 ;
  LAYER VI2 ;
  RECT 2679.800 45.560 2680.660 46.160 ;
  LAYER VI2 ;
  RECT 2680.200 45.620 2680.400 45.820 ;
  LAYER VI2 ;
  RECT 2679.800 45.620 2680.000 45.820 ;
  LAYER VI3 ;
  RECT 2679.800 57.100 2680.660 61.420 ;
  LAYER VI3 ;
  RECT 2680.260 61.100 2680.460 61.300 ;
  LAYER VI3 ;
  RECT 2680.260 60.700 2680.460 60.900 ;
  LAYER VI3 ;
  RECT 2680.260 60.300 2680.460 60.500 ;
  LAYER VI3 ;
  RECT 2680.260 59.900 2680.460 60.100 ;
  LAYER VI3 ;
  RECT 2680.260 59.500 2680.460 59.700 ;
  LAYER VI3 ;
  RECT 2680.260 59.100 2680.460 59.300 ;
  LAYER VI3 ;
  RECT 2680.260 58.700 2680.460 58.900 ;
  LAYER VI3 ;
  RECT 2680.260 58.300 2680.460 58.500 ;
  LAYER VI3 ;
  RECT 2680.260 57.900 2680.460 58.100 ;
  LAYER VI3 ;
  RECT 2680.260 57.500 2680.460 57.700 ;
  LAYER VI3 ;
  RECT 2680.260 57.100 2680.460 57.300 ;
  LAYER VI3 ;
  RECT 2679.860 61.100 2680.060 61.300 ;
  LAYER VI3 ;
  RECT 2679.860 60.700 2680.060 60.900 ;
  LAYER VI3 ;
  RECT 2679.860 60.300 2680.060 60.500 ;
  LAYER VI3 ;
  RECT 2679.860 59.900 2680.060 60.100 ;
  LAYER VI3 ;
  RECT 2679.860 59.500 2680.060 59.700 ;
  LAYER VI3 ;
  RECT 2679.860 59.100 2680.060 59.300 ;
  LAYER VI3 ;
  RECT 2679.860 58.700 2680.060 58.900 ;
  LAYER VI3 ;
  RECT 2679.860 58.300 2680.060 58.500 ;
  LAYER VI3 ;
  RECT 2679.860 57.900 2680.060 58.100 ;
  LAYER VI3 ;
  RECT 2679.860 57.500 2680.060 57.700 ;
  LAYER VI3 ;
  RECT 2679.860 57.100 2680.060 57.300 ;
  LAYER VI2 ;
  RECT 2679.800 57.100 2680.660 61.420 ;
  LAYER VI2 ;
  RECT 2680.260 61.100 2680.460 61.300 ;
  LAYER VI2 ;
  RECT 2680.260 60.700 2680.460 60.900 ;
  LAYER VI2 ;
  RECT 2680.260 60.300 2680.460 60.500 ;
  LAYER VI2 ;
  RECT 2680.260 59.900 2680.460 60.100 ;
  LAYER VI2 ;
  RECT 2680.260 59.500 2680.460 59.700 ;
  LAYER VI2 ;
  RECT 2680.260 59.100 2680.460 59.300 ;
  LAYER VI2 ;
  RECT 2680.260 58.700 2680.460 58.900 ;
  LAYER VI2 ;
  RECT 2680.260 58.300 2680.460 58.500 ;
  LAYER VI2 ;
  RECT 2680.260 57.900 2680.460 58.100 ;
  LAYER VI2 ;
  RECT 2680.260 57.500 2680.460 57.700 ;
  LAYER VI2 ;
  RECT 2680.260 57.100 2680.460 57.300 ;
  LAYER VI2 ;
  RECT 2679.860 61.100 2680.060 61.300 ;
  LAYER VI2 ;
  RECT 2679.860 60.700 2680.060 60.900 ;
  LAYER VI2 ;
  RECT 2679.860 60.300 2680.060 60.500 ;
  LAYER VI2 ;
  RECT 2679.860 59.900 2680.060 60.100 ;
  LAYER VI2 ;
  RECT 2679.860 59.500 2680.060 59.700 ;
  LAYER VI2 ;
  RECT 2679.860 59.100 2680.060 59.300 ;
  LAYER VI2 ;
  RECT 2679.860 58.700 2680.060 58.900 ;
  LAYER VI2 ;
  RECT 2679.860 58.300 2680.060 58.500 ;
  LAYER VI2 ;
  RECT 2679.860 57.900 2680.060 58.100 ;
  LAYER VI2 ;
  RECT 2679.860 57.500 2680.060 57.700 ;
  LAYER VI2 ;
  RECT 2679.860 57.100 2680.060 57.300 ;
  LAYER VI3 ;
  RECT 2678.380 5.880 2679.520 6.740 ;
  LAYER VI3 ;
  RECT 2679.180 6.340 2679.380 6.540 ;
  LAYER VI3 ;
  RECT 2679.180 5.940 2679.380 6.140 ;
  LAYER VI3 ;
  RECT 2678.780 6.340 2678.980 6.540 ;
  LAYER VI3 ;
  RECT 2678.780 5.940 2678.980 6.140 ;
  LAYER VI3 ;
  RECT 2678.380 6.340 2678.580 6.540 ;
  LAYER VI3 ;
  RECT 2678.380 5.940 2678.580 6.140 ;
  LAYER VI3 ;
  RECT 1370.180 5.880 1378.180 6.740 ;
  LAYER VI3 ;
  RECT 1377.780 6.340 1377.980 6.540 ;
  LAYER VI3 ;
  RECT 1377.780 5.940 1377.980 6.140 ;
  LAYER VI3 ;
  RECT 1377.380 6.340 1377.580 6.540 ;
  LAYER VI3 ;
  RECT 1377.380 5.940 1377.580 6.140 ;
  LAYER VI3 ;
  RECT 1376.980 6.340 1377.180 6.540 ;
  LAYER VI3 ;
  RECT 1376.980 5.940 1377.180 6.140 ;
  LAYER VI3 ;
  RECT 1376.580 6.340 1376.780 6.540 ;
  LAYER VI3 ;
  RECT 1376.580 5.940 1376.780 6.140 ;
  LAYER VI3 ;
  RECT 1376.180 6.340 1376.380 6.540 ;
  LAYER VI3 ;
  RECT 1376.180 5.940 1376.380 6.140 ;
  LAYER VI3 ;
  RECT 1375.780 6.340 1375.980 6.540 ;
  LAYER VI3 ;
  RECT 1375.780 5.940 1375.980 6.140 ;
  LAYER VI3 ;
  RECT 1375.380 6.340 1375.580 6.540 ;
  LAYER VI3 ;
  RECT 1375.380 5.940 1375.580 6.140 ;
  LAYER VI3 ;
  RECT 1374.980 6.340 1375.180 6.540 ;
  LAYER VI3 ;
  RECT 1374.980 5.940 1375.180 6.140 ;
  LAYER VI3 ;
  RECT 1374.580 6.340 1374.780 6.540 ;
  LAYER VI3 ;
  RECT 1374.580 5.940 1374.780 6.140 ;
  LAYER VI3 ;
  RECT 1374.180 6.340 1374.380 6.540 ;
  LAYER VI3 ;
  RECT 1374.180 5.940 1374.380 6.140 ;
  LAYER VI3 ;
  RECT 1373.780 6.340 1373.980 6.540 ;
  LAYER VI3 ;
  RECT 1373.780 5.940 1373.980 6.140 ;
  LAYER VI3 ;
  RECT 1373.380 6.340 1373.580 6.540 ;
  LAYER VI3 ;
  RECT 1373.380 5.940 1373.580 6.140 ;
  LAYER VI3 ;
  RECT 1372.980 6.340 1373.180 6.540 ;
  LAYER VI3 ;
  RECT 1372.980 5.940 1373.180 6.140 ;
  LAYER VI3 ;
  RECT 1372.580 6.340 1372.780 6.540 ;
  LAYER VI3 ;
  RECT 1372.580 5.940 1372.780 6.140 ;
  LAYER VI3 ;
  RECT 1372.180 6.340 1372.380 6.540 ;
  LAYER VI3 ;
  RECT 1372.180 5.940 1372.380 6.140 ;
  LAYER VI3 ;
  RECT 1371.780 6.340 1371.980 6.540 ;
  LAYER VI3 ;
  RECT 1371.780 5.940 1371.980 6.140 ;
  LAYER VI3 ;
  RECT 1371.380 6.340 1371.580 6.540 ;
  LAYER VI3 ;
  RECT 1371.380 5.940 1371.580 6.140 ;
  LAYER VI3 ;
  RECT 1370.980 6.340 1371.180 6.540 ;
  LAYER VI3 ;
  RECT 1370.980 5.940 1371.180 6.140 ;
  LAYER VI3 ;
  RECT 1370.580 6.340 1370.780 6.540 ;
  LAYER VI3 ;
  RECT 1370.580 5.940 1370.780 6.140 ;
  LAYER VI3 ;
  RECT 1370.180 6.340 1370.380 6.540 ;
  LAYER VI3 ;
  RECT 1370.180 5.940 1370.380 6.140 ;
  LAYER VI3 ;
  RECT 1390.020 5.880 1398.020 6.740 ;
  LAYER VI3 ;
  RECT 1397.620 6.340 1397.820 6.540 ;
  LAYER VI3 ;
  RECT 1397.620 5.940 1397.820 6.140 ;
  LAYER VI3 ;
  RECT 1397.220 6.340 1397.420 6.540 ;
  LAYER VI3 ;
  RECT 1397.220 5.940 1397.420 6.140 ;
  LAYER VI3 ;
  RECT 1396.820 6.340 1397.020 6.540 ;
  LAYER VI3 ;
  RECT 1396.820 5.940 1397.020 6.140 ;
  LAYER VI3 ;
  RECT 1396.420 6.340 1396.620 6.540 ;
  LAYER VI3 ;
  RECT 1396.420 5.940 1396.620 6.140 ;
  LAYER VI3 ;
  RECT 1396.020 6.340 1396.220 6.540 ;
  LAYER VI3 ;
  RECT 1396.020 5.940 1396.220 6.140 ;
  LAYER VI3 ;
  RECT 1395.620 6.340 1395.820 6.540 ;
  LAYER VI3 ;
  RECT 1395.620 5.940 1395.820 6.140 ;
  LAYER VI3 ;
  RECT 1395.220 6.340 1395.420 6.540 ;
  LAYER VI3 ;
  RECT 1395.220 5.940 1395.420 6.140 ;
  LAYER VI3 ;
  RECT 1394.820 6.340 1395.020 6.540 ;
  LAYER VI3 ;
  RECT 1394.820 5.940 1395.020 6.140 ;
  LAYER VI3 ;
  RECT 1394.420 6.340 1394.620 6.540 ;
  LAYER VI3 ;
  RECT 1394.420 5.940 1394.620 6.140 ;
  LAYER VI3 ;
  RECT 1394.020 6.340 1394.220 6.540 ;
  LAYER VI3 ;
  RECT 1394.020 5.940 1394.220 6.140 ;
  LAYER VI3 ;
  RECT 1393.620 6.340 1393.820 6.540 ;
  LAYER VI3 ;
  RECT 1393.620 5.940 1393.820 6.140 ;
  LAYER VI3 ;
  RECT 1393.220 6.340 1393.420 6.540 ;
  LAYER VI3 ;
  RECT 1393.220 5.940 1393.420 6.140 ;
  LAYER VI3 ;
  RECT 1392.820 6.340 1393.020 6.540 ;
  LAYER VI3 ;
  RECT 1392.820 5.940 1393.020 6.140 ;
  LAYER VI3 ;
  RECT 1392.420 6.340 1392.620 6.540 ;
  LAYER VI3 ;
  RECT 1392.420 5.940 1392.620 6.140 ;
  LAYER VI3 ;
  RECT 1392.020 6.340 1392.220 6.540 ;
  LAYER VI3 ;
  RECT 1392.020 5.940 1392.220 6.140 ;
  LAYER VI3 ;
  RECT 1391.620 6.340 1391.820 6.540 ;
  LAYER VI3 ;
  RECT 1391.620 5.940 1391.820 6.140 ;
  LAYER VI3 ;
  RECT 1391.220 6.340 1391.420 6.540 ;
  LAYER VI3 ;
  RECT 1391.220 5.940 1391.420 6.140 ;
  LAYER VI3 ;
  RECT 1390.820 6.340 1391.020 6.540 ;
  LAYER VI3 ;
  RECT 1390.820 5.940 1391.020 6.140 ;
  LAYER VI3 ;
  RECT 1390.420 6.340 1390.620 6.540 ;
  LAYER VI3 ;
  RECT 1390.420 5.940 1390.620 6.140 ;
  LAYER VI3 ;
  RECT 1390.020 6.340 1390.220 6.540 ;
  LAYER VI3 ;
  RECT 1390.020 5.940 1390.220 6.140 ;
  LAYER VI3 ;
  RECT 1411.100 5.880 1419.100 6.740 ;
  LAYER VI3 ;
  RECT 1418.700 6.340 1418.900 6.540 ;
  LAYER VI3 ;
  RECT 1418.700 5.940 1418.900 6.140 ;
  LAYER VI3 ;
  RECT 1418.300 6.340 1418.500 6.540 ;
  LAYER VI3 ;
  RECT 1418.300 5.940 1418.500 6.140 ;
  LAYER VI3 ;
  RECT 1417.900 6.340 1418.100 6.540 ;
  LAYER VI3 ;
  RECT 1417.900 5.940 1418.100 6.140 ;
  LAYER VI3 ;
  RECT 1417.500 6.340 1417.700 6.540 ;
  LAYER VI3 ;
  RECT 1417.500 5.940 1417.700 6.140 ;
  LAYER VI3 ;
  RECT 1417.100 6.340 1417.300 6.540 ;
  LAYER VI3 ;
  RECT 1417.100 5.940 1417.300 6.140 ;
  LAYER VI3 ;
  RECT 1416.700 6.340 1416.900 6.540 ;
  LAYER VI3 ;
  RECT 1416.700 5.940 1416.900 6.140 ;
  LAYER VI3 ;
  RECT 1416.300 6.340 1416.500 6.540 ;
  LAYER VI3 ;
  RECT 1416.300 5.940 1416.500 6.140 ;
  LAYER VI3 ;
  RECT 1415.900 6.340 1416.100 6.540 ;
  LAYER VI3 ;
  RECT 1415.900 5.940 1416.100 6.140 ;
  LAYER VI3 ;
  RECT 1415.500 6.340 1415.700 6.540 ;
  LAYER VI3 ;
  RECT 1415.500 5.940 1415.700 6.140 ;
  LAYER VI3 ;
  RECT 1415.100 6.340 1415.300 6.540 ;
  LAYER VI3 ;
  RECT 1415.100 5.940 1415.300 6.140 ;
  LAYER VI3 ;
  RECT 1414.700 6.340 1414.900 6.540 ;
  LAYER VI3 ;
  RECT 1414.700 5.940 1414.900 6.140 ;
  LAYER VI3 ;
  RECT 1414.300 6.340 1414.500 6.540 ;
  LAYER VI3 ;
  RECT 1414.300 5.940 1414.500 6.140 ;
  LAYER VI3 ;
  RECT 1413.900 6.340 1414.100 6.540 ;
  LAYER VI3 ;
  RECT 1413.900 5.940 1414.100 6.140 ;
  LAYER VI3 ;
  RECT 1413.500 6.340 1413.700 6.540 ;
  LAYER VI3 ;
  RECT 1413.500 5.940 1413.700 6.140 ;
  LAYER VI3 ;
  RECT 1413.100 6.340 1413.300 6.540 ;
  LAYER VI3 ;
  RECT 1413.100 5.940 1413.300 6.140 ;
  LAYER VI3 ;
  RECT 1412.700 6.340 1412.900 6.540 ;
  LAYER VI3 ;
  RECT 1412.700 5.940 1412.900 6.140 ;
  LAYER VI3 ;
  RECT 1412.300 6.340 1412.500 6.540 ;
  LAYER VI3 ;
  RECT 1412.300 5.940 1412.500 6.140 ;
  LAYER VI3 ;
  RECT 1411.900 6.340 1412.100 6.540 ;
  LAYER VI3 ;
  RECT 1411.900 5.940 1412.100 6.140 ;
  LAYER VI3 ;
  RECT 1411.500 6.340 1411.700 6.540 ;
  LAYER VI3 ;
  RECT 1411.500 5.940 1411.700 6.140 ;
  LAYER VI3 ;
  RECT 1411.100 6.340 1411.300 6.540 ;
  LAYER VI3 ;
  RECT 1411.100 5.940 1411.300 6.140 ;
  LAYER VI3 ;
  RECT 1430.940 5.880 1438.940 6.740 ;
  LAYER VI3 ;
  RECT 1438.540 6.340 1438.740 6.540 ;
  LAYER VI3 ;
  RECT 1438.540 5.940 1438.740 6.140 ;
  LAYER VI3 ;
  RECT 1438.140 6.340 1438.340 6.540 ;
  LAYER VI3 ;
  RECT 1438.140 5.940 1438.340 6.140 ;
  LAYER VI3 ;
  RECT 1437.740 6.340 1437.940 6.540 ;
  LAYER VI3 ;
  RECT 1437.740 5.940 1437.940 6.140 ;
  LAYER VI3 ;
  RECT 1437.340 6.340 1437.540 6.540 ;
  LAYER VI3 ;
  RECT 1437.340 5.940 1437.540 6.140 ;
  LAYER VI3 ;
  RECT 1436.940 6.340 1437.140 6.540 ;
  LAYER VI3 ;
  RECT 1436.940 5.940 1437.140 6.140 ;
  LAYER VI3 ;
  RECT 1436.540 6.340 1436.740 6.540 ;
  LAYER VI3 ;
  RECT 1436.540 5.940 1436.740 6.140 ;
  LAYER VI3 ;
  RECT 1436.140 6.340 1436.340 6.540 ;
  LAYER VI3 ;
  RECT 1436.140 5.940 1436.340 6.140 ;
  LAYER VI3 ;
  RECT 1435.740 6.340 1435.940 6.540 ;
  LAYER VI3 ;
  RECT 1435.740 5.940 1435.940 6.140 ;
  LAYER VI3 ;
  RECT 1435.340 6.340 1435.540 6.540 ;
  LAYER VI3 ;
  RECT 1435.340 5.940 1435.540 6.140 ;
  LAYER VI3 ;
  RECT 1434.940 6.340 1435.140 6.540 ;
  LAYER VI3 ;
  RECT 1434.940 5.940 1435.140 6.140 ;
  LAYER VI3 ;
  RECT 1434.540 6.340 1434.740 6.540 ;
  LAYER VI3 ;
  RECT 1434.540 5.940 1434.740 6.140 ;
  LAYER VI3 ;
  RECT 1434.140 6.340 1434.340 6.540 ;
  LAYER VI3 ;
  RECT 1434.140 5.940 1434.340 6.140 ;
  LAYER VI3 ;
  RECT 1433.740 6.340 1433.940 6.540 ;
  LAYER VI3 ;
  RECT 1433.740 5.940 1433.940 6.140 ;
  LAYER VI3 ;
  RECT 1433.340 6.340 1433.540 6.540 ;
  LAYER VI3 ;
  RECT 1433.340 5.940 1433.540 6.140 ;
  LAYER VI3 ;
  RECT 1432.940 6.340 1433.140 6.540 ;
  LAYER VI3 ;
  RECT 1432.940 5.940 1433.140 6.140 ;
  LAYER VI3 ;
  RECT 1432.540 6.340 1432.740 6.540 ;
  LAYER VI3 ;
  RECT 1432.540 5.940 1432.740 6.140 ;
  LAYER VI3 ;
  RECT 1432.140 6.340 1432.340 6.540 ;
  LAYER VI3 ;
  RECT 1432.140 5.940 1432.340 6.140 ;
  LAYER VI3 ;
  RECT 1431.740 6.340 1431.940 6.540 ;
  LAYER VI3 ;
  RECT 1431.740 5.940 1431.940 6.140 ;
  LAYER VI3 ;
  RECT 1431.340 6.340 1431.540 6.540 ;
  LAYER VI3 ;
  RECT 1431.340 5.940 1431.540 6.140 ;
  LAYER VI3 ;
  RECT 1430.940 6.340 1431.140 6.540 ;
  LAYER VI3 ;
  RECT 1430.940 5.940 1431.140 6.140 ;
  LAYER VI3 ;
  RECT 1452.020 5.880 1460.020 6.740 ;
  LAYER VI3 ;
  RECT 1459.620 6.340 1459.820 6.540 ;
  LAYER VI3 ;
  RECT 1459.620 5.940 1459.820 6.140 ;
  LAYER VI3 ;
  RECT 1459.220 6.340 1459.420 6.540 ;
  LAYER VI3 ;
  RECT 1459.220 5.940 1459.420 6.140 ;
  LAYER VI3 ;
  RECT 1458.820 6.340 1459.020 6.540 ;
  LAYER VI3 ;
  RECT 1458.820 5.940 1459.020 6.140 ;
  LAYER VI3 ;
  RECT 1458.420 6.340 1458.620 6.540 ;
  LAYER VI3 ;
  RECT 1458.420 5.940 1458.620 6.140 ;
  LAYER VI3 ;
  RECT 1458.020 6.340 1458.220 6.540 ;
  LAYER VI3 ;
  RECT 1458.020 5.940 1458.220 6.140 ;
  LAYER VI3 ;
  RECT 1457.620 6.340 1457.820 6.540 ;
  LAYER VI3 ;
  RECT 1457.620 5.940 1457.820 6.140 ;
  LAYER VI3 ;
  RECT 1457.220 6.340 1457.420 6.540 ;
  LAYER VI3 ;
  RECT 1457.220 5.940 1457.420 6.140 ;
  LAYER VI3 ;
  RECT 1456.820 6.340 1457.020 6.540 ;
  LAYER VI3 ;
  RECT 1456.820 5.940 1457.020 6.140 ;
  LAYER VI3 ;
  RECT 1456.420 6.340 1456.620 6.540 ;
  LAYER VI3 ;
  RECT 1456.420 5.940 1456.620 6.140 ;
  LAYER VI3 ;
  RECT 1456.020 6.340 1456.220 6.540 ;
  LAYER VI3 ;
  RECT 1456.020 5.940 1456.220 6.140 ;
  LAYER VI3 ;
  RECT 1455.620 6.340 1455.820 6.540 ;
  LAYER VI3 ;
  RECT 1455.620 5.940 1455.820 6.140 ;
  LAYER VI3 ;
  RECT 1455.220 6.340 1455.420 6.540 ;
  LAYER VI3 ;
  RECT 1455.220 5.940 1455.420 6.140 ;
  LAYER VI3 ;
  RECT 1454.820 6.340 1455.020 6.540 ;
  LAYER VI3 ;
  RECT 1454.820 5.940 1455.020 6.140 ;
  LAYER VI3 ;
  RECT 1454.420 6.340 1454.620 6.540 ;
  LAYER VI3 ;
  RECT 1454.420 5.940 1454.620 6.140 ;
  LAYER VI3 ;
  RECT 1454.020 6.340 1454.220 6.540 ;
  LAYER VI3 ;
  RECT 1454.020 5.940 1454.220 6.140 ;
  LAYER VI3 ;
  RECT 1453.620 6.340 1453.820 6.540 ;
  LAYER VI3 ;
  RECT 1453.620 5.940 1453.820 6.140 ;
  LAYER VI3 ;
  RECT 1453.220 6.340 1453.420 6.540 ;
  LAYER VI3 ;
  RECT 1453.220 5.940 1453.420 6.140 ;
  LAYER VI3 ;
  RECT 1452.820 6.340 1453.020 6.540 ;
  LAYER VI3 ;
  RECT 1452.820 5.940 1453.020 6.140 ;
  LAYER VI3 ;
  RECT 1452.420 6.340 1452.620 6.540 ;
  LAYER VI3 ;
  RECT 1452.420 5.940 1452.620 6.140 ;
  LAYER VI3 ;
  RECT 1452.020 6.340 1452.220 6.540 ;
  LAYER VI3 ;
  RECT 1452.020 5.940 1452.220 6.140 ;
  LAYER VI3 ;
  RECT 1471.860 5.880 1479.860 6.740 ;
  LAYER VI3 ;
  RECT 1479.460 6.340 1479.660 6.540 ;
  LAYER VI3 ;
  RECT 1479.460 5.940 1479.660 6.140 ;
  LAYER VI3 ;
  RECT 1479.060 6.340 1479.260 6.540 ;
  LAYER VI3 ;
  RECT 1479.060 5.940 1479.260 6.140 ;
  LAYER VI3 ;
  RECT 1478.660 6.340 1478.860 6.540 ;
  LAYER VI3 ;
  RECT 1478.660 5.940 1478.860 6.140 ;
  LAYER VI3 ;
  RECT 1478.260 6.340 1478.460 6.540 ;
  LAYER VI3 ;
  RECT 1478.260 5.940 1478.460 6.140 ;
  LAYER VI3 ;
  RECT 1477.860 6.340 1478.060 6.540 ;
  LAYER VI3 ;
  RECT 1477.860 5.940 1478.060 6.140 ;
  LAYER VI3 ;
  RECT 1477.460 6.340 1477.660 6.540 ;
  LAYER VI3 ;
  RECT 1477.460 5.940 1477.660 6.140 ;
  LAYER VI3 ;
  RECT 1477.060 6.340 1477.260 6.540 ;
  LAYER VI3 ;
  RECT 1477.060 5.940 1477.260 6.140 ;
  LAYER VI3 ;
  RECT 1476.660 6.340 1476.860 6.540 ;
  LAYER VI3 ;
  RECT 1476.660 5.940 1476.860 6.140 ;
  LAYER VI3 ;
  RECT 1476.260 6.340 1476.460 6.540 ;
  LAYER VI3 ;
  RECT 1476.260 5.940 1476.460 6.140 ;
  LAYER VI3 ;
  RECT 1475.860 6.340 1476.060 6.540 ;
  LAYER VI3 ;
  RECT 1475.860 5.940 1476.060 6.140 ;
  LAYER VI3 ;
  RECT 1475.460 6.340 1475.660 6.540 ;
  LAYER VI3 ;
  RECT 1475.460 5.940 1475.660 6.140 ;
  LAYER VI3 ;
  RECT 1475.060 6.340 1475.260 6.540 ;
  LAYER VI3 ;
  RECT 1475.060 5.940 1475.260 6.140 ;
  LAYER VI3 ;
  RECT 1474.660 6.340 1474.860 6.540 ;
  LAYER VI3 ;
  RECT 1474.660 5.940 1474.860 6.140 ;
  LAYER VI3 ;
  RECT 1474.260 6.340 1474.460 6.540 ;
  LAYER VI3 ;
  RECT 1474.260 5.940 1474.460 6.140 ;
  LAYER VI3 ;
  RECT 1473.860 6.340 1474.060 6.540 ;
  LAYER VI3 ;
  RECT 1473.860 5.940 1474.060 6.140 ;
  LAYER VI3 ;
  RECT 1473.460 6.340 1473.660 6.540 ;
  LAYER VI3 ;
  RECT 1473.460 5.940 1473.660 6.140 ;
  LAYER VI3 ;
  RECT 1473.060 6.340 1473.260 6.540 ;
  LAYER VI3 ;
  RECT 1473.060 5.940 1473.260 6.140 ;
  LAYER VI3 ;
  RECT 1472.660 6.340 1472.860 6.540 ;
  LAYER VI3 ;
  RECT 1472.660 5.940 1472.860 6.140 ;
  LAYER VI3 ;
  RECT 1472.260 6.340 1472.460 6.540 ;
  LAYER VI3 ;
  RECT 1472.260 5.940 1472.460 6.140 ;
  LAYER VI3 ;
  RECT 1471.860 6.340 1472.060 6.540 ;
  LAYER VI3 ;
  RECT 1471.860 5.940 1472.060 6.140 ;
  LAYER VI3 ;
  RECT 1492.940 5.880 1500.940 6.740 ;
  LAYER VI3 ;
  RECT 1500.540 6.340 1500.740 6.540 ;
  LAYER VI3 ;
  RECT 1500.540 5.940 1500.740 6.140 ;
  LAYER VI3 ;
  RECT 1500.140 6.340 1500.340 6.540 ;
  LAYER VI3 ;
  RECT 1500.140 5.940 1500.340 6.140 ;
  LAYER VI3 ;
  RECT 1499.740 6.340 1499.940 6.540 ;
  LAYER VI3 ;
  RECT 1499.740 5.940 1499.940 6.140 ;
  LAYER VI3 ;
  RECT 1499.340 6.340 1499.540 6.540 ;
  LAYER VI3 ;
  RECT 1499.340 5.940 1499.540 6.140 ;
  LAYER VI3 ;
  RECT 1498.940 6.340 1499.140 6.540 ;
  LAYER VI3 ;
  RECT 1498.940 5.940 1499.140 6.140 ;
  LAYER VI3 ;
  RECT 1498.540 6.340 1498.740 6.540 ;
  LAYER VI3 ;
  RECT 1498.540 5.940 1498.740 6.140 ;
  LAYER VI3 ;
  RECT 1498.140 6.340 1498.340 6.540 ;
  LAYER VI3 ;
  RECT 1498.140 5.940 1498.340 6.140 ;
  LAYER VI3 ;
  RECT 1497.740 6.340 1497.940 6.540 ;
  LAYER VI3 ;
  RECT 1497.740 5.940 1497.940 6.140 ;
  LAYER VI3 ;
  RECT 1497.340 6.340 1497.540 6.540 ;
  LAYER VI3 ;
  RECT 1497.340 5.940 1497.540 6.140 ;
  LAYER VI3 ;
  RECT 1496.940 6.340 1497.140 6.540 ;
  LAYER VI3 ;
  RECT 1496.940 5.940 1497.140 6.140 ;
  LAYER VI3 ;
  RECT 1496.540 6.340 1496.740 6.540 ;
  LAYER VI3 ;
  RECT 1496.540 5.940 1496.740 6.140 ;
  LAYER VI3 ;
  RECT 1496.140 6.340 1496.340 6.540 ;
  LAYER VI3 ;
  RECT 1496.140 5.940 1496.340 6.140 ;
  LAYER VI3 ;
  RECT 1495.740 6.340 1495.940 6.540 ;
  LAYER VI3 ;
  RECT 1495.740 5.940 1495.940 6.140 ;
  LAYER VI3 ;
  RECT 1495.340 6.340 1495.540 6.540 ;
  LAYER VI3 ;
  RECT 1495.340 5.940 1495.540 6.140 ;
  LAYER VI3 ;
  RECT 1494.940 6.340 1495.140 6.540 ;
  LAYER VI3 ;
  RECT 1494.940 5.940 1495.140 6.140 ;
  LAYER VI3 ;
  RECT 1494.540 6.340 1494.740 6.540 ;
  LAYER VI3 ;
  RECT 1494.540 5.940 1494.740 6.140 ;
  LAYER VI3 ;
  RECT 1494.140 6.340 1494.340 6.540 ;
  LAYER VI3 ;
  RECT 1494.140 5.940 1494.340 6.140 ;
  LAYER VI3 ;
  RECT 1493.740 6.340 1493.940 6.540 ;
  LAYER VI3 ;
  RECT 1493.740 5.940 1493.940 6.140 ;
  LAYER VI3 ;
  RECT 1493.340 6.340 1493.540 6.540 ;
  LAYER VI3 ;
  RECT 1493.340 5.940 1493.540 6.140 ;
  LAYER VI3 ;
  RECT 1492.940 6.340 1493.140 6.540 ;
  LAYER VI3 ;
  RECT 1492.940 5.940 1493.140 6.140 ;
  LAYER VI3 ;
  RECT 1512.780 5.880 1520.780 6.740 ;
  LAYER VI3 ;
  RECT 1520.380 6.340 1520.580 6.540 ;
  LAYER VI3 ;
  RECT 1520.380 5.940 1520.580 6.140 ;
  LAYER VI3 ;
  RECT 1519.980 6.340 1520.180 6.540 ;
  LAYER VI3 ;
  RECT 1519.980 5.940 1520.180 6.140 ;
  LAYER VI3 ;
  RECT 1519.580 6.340 1519.780 6.540 ;
  LAYER VI3 ;
  RECT 1519.580 5.940 1519.780 6.140 ;
  LAYER VI3 ;
  RECT 1519.180 6.340 1519.380 6.540 ;
  LAYER VI3 ;
  RECT 1519.180 5.940 1519.380 6.140 ;
  LAYER VI3 ;
  RECT 1518.780 6.340 1518.980 6.540 ;
  LAYER VI3 ;
  RECT 1518.780 5.940 1518.980 6.140 ;
  LAYER VI3 ;
  RECT 1518.380 6.340 1518.580 6.540 ;
  LAYER VI3 ;
  RECT 1518.380 5.940 1518.580 6.140 ;
  LAYER VI3 ;
  RECT 1517.980 6.340 1518.180 6.540 ;
  LAYER VI3 ;
  RECT 1517.980 5.940 1518.180 6.140 ;
  LAYER VI3 ;
  RECT 1517.580 6.340 1517.780 6.540 ;
  LAYER VI3 ;
  RECT 1517.580 5.940 1517.780 6.140 ;
  LAYER VI3 ;
  RECT 1517.180 6.340 1517.380 6.540 ;
  LAYER VI3 ;
  RECT 1517.180 5.940 1517.380 6.140 ;
  LAYER VI3 ;
  RECT 1516.780 6.340 1516.980 6.540 ;
  LAYER VI3 ;
  RECT 1516.780 5.940 1516.980 6.140 ;
  LAYER VI3 ;
  RECT 1516.380 6.340 1516.580 6.540 ;
  LAYER VI3 ;
  RECT 1516.380 5.940 1516.580 6.140 ;
  LAYER VI3 ;
  RECT 1515.980 6.340 1516.180 6.540 ;
  LAYER VI3 ;
  RECT 1515.980 5.940 1516.180 6.140 ;
  LAYER VI3 ;
  RECT 1515.580 6.340 1515.780 6.540 ;
  LAYER VI3 ;
  RECT 1515.580 5.940 1515.780 6.140 ;
  LAYER VI3 ;
  RECT 1515.180 6.340 1515.380 6.540 ;
  LAYER VI3 ;
  RECT 1515.180 5.940 1515.380 6.140 ;
  LAYER VI3 ;
  RECT 1514.780 6.340 1514.980 6.540 ;
  LAYER VI3 ;
  RECT 1514.780 5.940 1514.980 6.140 ;
  LAYER VI3 ;
  RECT 1514.380 6.340 1514.580 6.540 ;
  LAYER VI3 ;
  RECT 1514.380 5.940 1514.580 6.140 ;
  LAYER VI3 ;
  RECT 1513.980 6.340 1514.180 6.540 ;
  LAYER VI3 ;
  RECT 1513.980 5.940 1514.180 6.140 ;
  LAYER VI3 ;
  RECT 1513.580 6.340 1513.780 6.540 ;
  LAYER VI3 ;
  RECT 1513.580 5.940 1513.780 6.140 ;
  LAYER VI3 ;
  RECT 1513.180 6.340 1513.380 6.540 ;
  LAYER VI3 ;
  RECT 1513.180 5.940 1513.380 6.140 ;
  LAYER VI3 ;
  RECT 1512.780 6.340 1512.980 6.540 ;
  LAYER VI3 ;
  RECT 1512.780 5.940 1512.980 6.140 ;
  LAYER VI3 ;
  RECT 1533.860 5.880 1541.860 6.740 ;
  LAYER VI3 ;
  RECT 1541.460 6.340 1541.660 6.540 ;
  LAYER VI3 ;
  RECT 1541.460 5.940 1541.660 6.140 ;
  LAYER VI3 ;
  RECT 1541.060 6.340 1541.260 6.540 ;
  LAYER VI3 ;
  RECT 1541.060 5.940 1541.260 6.140 ;
  LAYER VI3 ;
  RECT 1540.660 6.340 1540.860 6.540 ;
  LAYER VI3 ;
  RECT 1540.660 5.940 1540.860 6.140 ;
  LAYER VI3 ;
  RECT 1540.260 6.340 1540.460 6.540 ;
  LAYER VI3 ;
  RECT 1540.260 5.940 1540.460 6.140 ;
  LAYER VI3 ;
  RECT 1539.860 6.340 1540.060 6.540 ;
  LAYER VI3 ;
  RECT 1539.860 5.940 1540.060 6.140 ;
  LAYER VI3 ;
  RECT 1539.460 6.340 1539.660 6.540 ;
  LAYER VI3 ;
  RECT 1539.460 5.940 1539.660 6.140 ;
  LAYER VI3 ;
  RECT 1539.060 6.340 1539.260 6.540 ;
  LAYER VI3 ;
  RECT 1539.060 5.940 1539.260 6.140 ;
  LAYER VI3 ;
  RECT 1538.660 6.340 1538.860 6.540 ;
  LAYER VI3 ;
  RECT 1538.660 5.940 1538.860 6.140 ;
  LAYER VI3 ;
  RECT 1538.260 6.340 1538.460 6.540 ;
  LAYER VI3 ;
  RECT 1538.260 5.940 1538.460 6.140 ;
  LAYER VI3 ;
  RECT 1537.860 6.340 1538.060 6.540 ;
  LAYER VI3 ;
  RECT 1537.860 5.940 1538.060 6.140 ;
  LAYER VI3 ;
  RECT 1537.460 6.340 1537.660 6.540 ;
  LAYER VI3 ;
  RECT 1537.460 5.940 1537.660 6.140 ;
  LAYER VI3 ;
  RECT 1537.060 6.340 1537.260 6.540 ;
  LAYER VI3 ;
  RECT 1537.060 5.940 1537.260 6.140 ;
  LAYER VI3 ;
  RECT 1536.660 6.340 1536.860 6.540 ;
  LAYER VI3 ;
  RECT 1536.660 5.940 1536.860 6.140 ;
  LAYER VI3 ;
  RECT 1536.260 6.340 1536.460 6.540 ;
  LAYER VI3 ;
  RECT 1536.260 5.940 1536.460 6.140 ;
  LAYER VI3 ;
  RECT 1535.860 6.340 1536.060 6.540 ;
  LAYER VI3 ;
  RECT 1535.860 5.940 1536.060 6.140 ;
  LAYER VI3 ;
  RECT 1535.460 6.340 1535.660 6.540 ;
  LAYER VI3 ;
  RECT 1535.460 5.940 1535.660 6.140 ;
  LAYER VI3 ;
  RECT 1535.060 6.340 1535.260 6.540 ;
  LAYER VI3 ;
  RECT 1535.060 5.940 1535.260 6.140 ;
  LAYER VI3 ;
  RECT 1534.660 6.340 1534.860 6.540 ;
  LAYER VI3 ;
  RECT 1534.660 5.940 1534.860 6.140 ;
  LAYER VI3 ;
  RECT 1534.260 6.340 1534.460 6.540 ;
  LAYER VI3 ;
  RECT 1534.260 5.940 1534.460 6.140 ;
  LAYER VI3 ;
  RECT 1533.860 6.340 1534.060 6.540 ;
  LAYER VI3 ;
  RECT 1533.860 5.940 1534.060 6.140 ;
  LAYER VI3 ;
  RECT 1553.700 5.880 1561.700 6.740 ;
  LAYER VI3 ;
  RECT 1561.300 6.340 1561.500 6.540 ;
  LAYER VI3 ;
  RECT 1561.300 5.940 1561.500 6.140 ;
  LAYER VI3 ;
  RECT 1560.900 6.340 1561.100 6.540 ;
  LAYER VI3 ;
  RECT 1560.900 5.940 1561.100 6.140 ;
  LAYER VI3 ;
  RECT 1560.500 6.340 1560.700 6.540 ;
  LAYER VI3 ;
  RECT 1560.500 5.940 1560.700 6.140 ;
  LAYER VI3 ;
  RECT 1560.100 6.340 1560.300 6.540 ;
  LAYER VI3 ;
  RECT 1560.100 5.940 1560.300 6.140 ;
  LAYER VI3 ;
  RECT 1559.700 6.340 1559.900 6.540 ;
  LAYER VI3 ;
  RECT 1559.700 5.940 1559.900 6.140 ;
  LAYER VI3 ;
  RECT 1559.300 6.340 1559.500 6.540 ;
  LAYER VI3 ;
  RECT 1559.300 5.940 1559.500 6.140 ;
  LAYER VI3 ;
  RECT 1558.900 6.340 1559.100 6.540 ;
  LAYER VI3 ;
  RECT 1558.900 5.940 1559.100 6.140 ;
  LAYER VI3 ;
  RECT 1558.500 6.340 1558.700 6.540 ;
  LAYER VI3 ;
  RECT 1558.500 5.940 1558.700 6.140 ;
  LAYER VI3 ;
  RECT 1558.100 6.340 1558.300 6.540 ;
  LAYER VI3 ;
  RECT 1558.100 5.940 1558.300 6.140 ;
  LAYER VI3 ;
  RECT 1557.700 6.340 1557.900 6.540 ;
  LAYER VI3 ;
  RECT 1557.700 5.940 1557.900 6.140 ;
  LAYER VI3 ;
  RECT 1557.300 6.340 1557.500 6.540 ;
  LAYER VI3 ;
  RECT 1557.300 5.940 1557.500 6.140 ;
  LAYER VI3 ;
  RECT 1556.900 6.340 1557.100 6.540 ;
  LAYER VI3 ;
  RECT 1556.900 5.940 1557.100 6.140 ;
  LAYER VI3 ;
  RECT 1556.500 6.340 1556.700 6.540 ;
  LAYER VI3 ;
  RECT 1556.500 5.940 1556.700 6.140 ;
  LAYER VI3 ;
  RECT 1556.100 6.340 1556.300 6.540 ;
  LAYER VI3 ;
  RECT 1556.100 5.940 1556.300 6.140 ;
  LAYER VI3 ;
  RECT 1555.700 6.340 1555.900 6.540 ;
  LAYER VI3 ;
  RECT 1555.700 5.940 1555.900 6.140 ;
  LAYER VI3 ;
  RECT 1555.300 6.340 1555.500 6.540 ;
  LAYER VI3 ;
  RECT 1555.300 5.940 1555.500 6.140 ;
  LAYER VI3 ;
  RECT 1554.900 6.340 1555.100 6.540 ;
  LAYER VI3 ;
  RECT 1554.900 5.940 1555.100 6.140 ;
  LAYER VI3 ;
  RECT 1554.500 6.340 1554.700 6.540 ;
  LAYER VI3 ;
  RECT 1554.500 5.940 1554.700 6.140 ;
  LAYER VI3 ;
  RECT 1554.100 6.340 1554.300 6.540 ;
  LAYER VI3 ;
  RECT 1554.100 5.940 1554.300 6.140 ;
  LAYER VI3 ;
  RECT 1553.700 6.340 1553.900 6.540 ;
  LAYER VI3 ;
  RECT 1553.700 5.940 1553.900 6.140 ;
  LAYER VI3 ;
  RECT 1574.780 5.880 1582.780 6.740 ;
  LAYER VI3 ;
  RECT 1582.380 6.340 1582.580 6.540 ;
  LAYER VI3 ;
  RECT 1582.380 5.940 1582.580 6.140 ;
  LAYER VI3 ;
  RECT 1581.980 6.340 1582.180 6.540 ;
  LAYER VI3 ;
  RECT 1581.980 5.940 1582.180 6.140 ;
  LAYER VI3 ;
  RECT 1581.580 6.340 1581.780 6.540 ;
  LAYER VI3 ;
  RECT 1581.580 5.940 1581.780 6.140 ;
  LAYER VI3 ;
  RECT 1581.180 6.340 1581.380 6.540 ;
  LAYER VI3 ;
  RECT 1581.180 5.940 1581.380 6.140 ;
  LAYER VI3 ;
  RECT 1580.780 6.340 1580.980 6.540 ;
  LAYER VI3 ;
  RECT 1580.780 5.940 1580.980 6.140 ;
  LAYER VI3 ;
  RECT 1580.380 6.340 1580.580 6.540 ;
  LAYER VI3 ;
  RECT 1580.380 5.940 1580.580 6.140 ;
  LAYER VI3 ;
  RECT 1579.980 6.340 1580.180 6.540 ;
  LAYER VI3 ;
  RECT 1579.980 5.940 1580.180 6.140 ;
  LAYER VI3 ;
  RECT 1579.580 6.340 1579.780 6.540 ;
  LAYER VI3 ;
  RECT 1579.580 5.940 1579.780 6.140 ;
  LAYER VI3 ;
  RECT 1579.180 6.340 1579.380 6.540 ;
  LAYER VI3 ;
  RECT 1579.180 5.940 1579.380 6.140 ;
  LAYER VI3 ;
  RECT 1578.780 6.340 1578.980 6.540 ;
  LAYER VI3 ;
  RECT 1578.780 5.940 1578.980 6.140 ;
  LAYER VI3 ;
  RECT 1578.380 6.340 1578.580 6.540 ;
  LAYER VI3 ;
  RECT 1578.380 5.940 1578.580 6.140 ;
  LAYER VI3 ;
  RECT 1577.980 6.340 1578.180 6.540 ;
  LAYER VI3 ;
  RECT 1577.980 5.940 1578.180 6.140 ;
  LAYER VI3 ;
  RECT 1577.580 6.340 1577.780 6.540 ;
  LAYER VI3 ;
  RECT 1577.580 5.940 1577.780 6.140 ;
  LAYER VI3 ;
  RECT 1577.180 6.340 1577.380 6.540 ;
  LAYER VI3 ;
  RECT 1577.180 5.940 1577.380 6.140 ;
  LAYER VI3 ;
  RECT 1576.780 6.340 1576.980 6.540 ;
  LAYER VI3 ;
  RECT 1576.780 5.940 1576.980 6.140 ;
  LAYER VI3 ;
  RECT 1576.380 6.340 1576.580 6.540 ;
  LAYER VI3 ;
  RECT 1576.380 5.940 1576.580 6.140 ;
  LAYER VI3 ;
  RECT 1575.980 6.340 1576.180 6.540 ;
  LAYER VI3 ;
  RECT 1575.980 5.940 1576.180 6.140 ;
  LAYER VI3 ;
  RECT 1575.580 6.340 1575.780 6.540 ;
  LAYER VI3 ;
  RECT 1575.580 5.940 1575.780 6.140 ;
  LAYER VI3 ;
  RECT 1575.180 6.340 1575.380 6.540 ;
  LAYER VI3 ;
  RECT 1575.180 5.940 1575.380 6.140 ;
  LAYER VI3 ;
  RECT 1574.780 6.340 1574.980 6.540 ;
  LAYER VI3 ;
  RECT 1574.780 5.940 1574.980 6.140 ;
  LAYER VI3 ;
  RECT 1594.620 5.880 1602.620 6.740 ;
  LAYER VI3 ;
  RECT 1602.220 6.340 1602.420 6.540 ;
  LAYER VI3 ;
  RECT 1602.220 5.940 1602.420 6.140 ;
  LAYER VI3 ;
  RECT 1601.820 6.340 1602.020 6.540 ;
  LAYER VI3 ;
  RECT 1601.820 5.940 1602.020 6.140 ;
  LAYER VI3 ;
  RECT 1601.420 6.340 1601.620 6.540 ;
  LAYER VI3 ;
  RECT 1601.420 5.940 1601.620 6.140 ;
  LAYER VI3 ;
  RECT 1601.020 6.340 1601.220 6.540 ;
  LAYER VI3 ;
  RECT 1601.020 5.940 1601.220 6.140 ;
  LAYER VI3 ;
  RECT 1600.620 6.340 1600.820 6.540 ;
  LAYER VI3 ;
  RECT 1600.620 5.940 1600.820 6.140 ;
  LAYER VI3 ;
  RECT 1600.220 6.340 1600.420 6.540 ;
  LAYER VI3 ;
  RECT 1600.220 5.940 1600.420 6.140 ;
  LAYER VI3 ;
  RECT 1599.820 6.340 1600.020 6.540 ;
  LAYER VI3 ;
  RECT 1599.820 5.940 1600.020 6.140 ;
  LAYER VI3 ;
  RECT 1599.420 6.340 1599.620 6.540 ;
  LAYER VI3 ;
  RECT 1599.420 5.940 1599.620 6.140 ;
  LAYER VI3 ;
  RECT 1599.020 6.340 1599.220 6.540 ;
  LAYER VI3 ;
  RECT 1599.020 5.940 1599.220 6.140 ;
  LAYER VI3 ;
  RECT 1598.620 6.340 1598.820 6.540 ;
  LAYER VI3 ;
  RECT 1598.620 5.940 1598.820 6.140 ;
  LAYER VI3 ;
  RECT 1598.220 6.340 1598.420 6.540 ;
  LAYER VI3 ;
  RECT 1598.220 5.940 1598.420 6.140 ;
  LAYER VI3 ;
  RECT 1597.820 6.340 1598.020 6.540 ;
  LAYER VI3 ;
  RECT 1597.820 5.940 1598.020 6.140 ;
  LAYER VI3 ;
  RECT 1597.420 6.340 1597.620 6.540 ;
  LAYER VI3 ;
  RECT 1597.420 5.940 1597.620 6.140 ;
  LAYER VI3 ;
  RECT 1597.020 6.340 1597.220 6.540 ;
  LAYER VI3 ;
  RECT 1597.020 5.940 1597.220 6.140 ;
  LAYER VI3 ;
  RECT 1596.620 6.340 1596.820 6.540 ;
  LAYER VI3 ;
  RECT 1596.620 5.940 1596.820 6.140 ;
  LAYER VI3 ;
  RECT 1596.220 6.340 1596.420 6.540 ;
  LAYER VI3 ;
  RECT 1596.220 5.940 1596.420 6.140 ;
  LAYER VI3 ;
  RECT 1595.820 6.340 1596.020 6.540 ;
  LAYER VI3 ;
  RECT 1595.820 5.940 1596.020 6.140 ;
  LAYER VI3 ;
  RECT 1595.420 6.340 1595.620 6.540 ;
  LAYER VI3 ;
  RECT 1595.420 5.940 1595.620 6.140 ;
  LAYER VI3 ;
  RECT 1595.020 6.340 1595.220 6.540 ;
  LAYER VI3 ;
  RECT 1595.020 5.940 1595.220 6.140 ;
  LAYER VI3 ;
  RECT 1594.620 6.340 1594.820 6.540 ;
  LAYER VI3 ;
  RECT 1594.620 5.940 1594.820 6.140 ;
  LAYER VI3 ;
  RECT 1615.700 5.880 1623.700 6.740 ;
  LAYER VI3 ;
  RECT 1623.300 6.340 1623.500 6.540 ;
  LAYER VI3 ;
  RECT 1623.300 5.940 1623.500 6.140 ;
  LAYER VI3 ;
  RECT 1622.900 6.340 1623.100 6.540 ;
  LAYER VI3 ;
  RECT 1622.900 5.940 1623.100 6.140 ;
  LAYER VI3 ;
  RECT 1622.500 6.340 1622.700 6.540 ;
  LAYER VI3 ;
  RECT 1622.500 5.940 1622.700 6.140 ;
  LAYER VI3 ;
  RECT 1622.100 6.340 1622.300 6.540 ;
  LAYER VI3 ;
  RECT 1622.100 5.940 1622.300 6.140 ;
  LAYER VI3 ;
  RECT 1621.700 6.340 1621.900 6.540 ;
  LAYER VI3 ;
  RECT 1621.700 5.940 1621.900 6.140 ;
  LAYER VI3 ;
  RECT 1621.300 6.340 1621.500 6.540 ;
  LAYER VI3 ;
  RECT 1621.300 5.940 1621.500 6.140 ;
  LAYER VI3 ;
  RECT 1620.900 6.340 1621.100 6.540 ;
  LAYER VI3 ;
  RECT 1620.900 5.940 1621.100 6.140 ;
  LAYER VI3 ;
  RECT 1620.500 6.340 1620.700 6.540 ;
  LAYER VI3 ;
  RECT 1620.500 5.940 1620.700 6.140 ;
  LAYER VI3 ;
  RECT 1620.100 6.340 1620.300 6.540 ;
  LAYER VI3 ;
  RECT 1620.100 5.940 1620.300 6.140 ;
  LAYER VI3 ;
  RECT 1619.700 6.340 1619.900 6.540 ;
  LAYER VI3 ;
  RECT 1619.700 5.940 1619.900 6.140 ;
  LAYER VI3 ;
  RECT 1619.300 6.340 1619.500 6.540 ;
  LAYER VI3 ;
  RECT 1619.300 5.940 1619.500 6.140 ;
  LAYER VI3 ;
  RECT 1618.900 6.340 1619.100 6.540 ;
  LAYER VI3 ;
  RECT 1618.900 5.940 1619.100 6.140 ;
  LAYER VI3 ;
  RECT 1618.500 6.340 1618.700 6.540 ;
  LAYER VI3 ;
  RECT 1618.500 5.940 1618.700 6.140 ;
  LAYER VI3 ;
  RECT 1618.100 6.340 1618.300 6.540 ;
  LAYER VI3 ;
  RECT 1618.100 5.940 1618.300 6.140 ;
  LAYER VI3 ;
  RECT 1617.700 6.340 1617.900 6.540 ;
  LAYER VI3 ;
  RECT 1617.700 5.940 1617.900 6.140 ;
  LAYER VI3 ;
  RECT 1617.300 6.340 1617.500 6.540 ;
  LAYER VI3 ;
  RECT 1617.300 5.940 1617.500 6.140 ;
  LAYER VI3 ;
  RECT 1616.900 6.340 1617.100 6.540 ;
  LAYER VI3 ;
  RECT 1616.900 5.940 1617.100 6.140 ;
  LAYER VI3 ;
  RECT 1616.500 6.340 1616.700 6.540 ;
  LAYER VI3 ;
  RECT 1616.500 5.940 1616.700 6.140 ;
  LAYER VI3 ;
  RECT 1616.100 6.340 1616.300 6.540 ;
  LAYER VI3 ;
  RECT 1616.100 5.940 1616.300 6.140 ;
  LAYER VI3 ;
  RECT 1615.700 6.340 1615.900 6.540 ;
  LAYER VI3 ;
  RECT 1615.700 5.940 1615.900 6.140 ;
  LAYER VI3 ;
  RECT 1635.540 5.880 1643.540 6.740 ;
  LAYER VI3 ;
  RECT 1643.140 6.340 1643.340 6.540 ;
  LAYER VI3 ;
  RECT 1643.140 5.940 1643.340 6.140 ;
  LAYER VI3 ;
  RECT 1642.740 6.340 1642.940 6.540 ;
  LAYER VI3 ;
  RECT 1642.740 5.940 1642.940 6.140 ;
  LAYER VI3 ;
  RECT 1642.340 6.340 1642.540 6.540 ;
  LAYER VI3 ;
  RECT 1642.340 5.940 1642.540 6.140 ;
  LAYER VI3 ;
  RECT 1641.940 6.340 1642.140 6.540 ;
  LAYER VI3 ;
  RECT 1641.940 5.940 1642.140 6.140 ;
  LAYER VI3 ;
  RECT 1641.540 6.340 1641.740 6.540 ;
  LAYER VI3 ;
  RECT 1641.540 5.940 1641.740 6.140 ;
  LAYER VI3 ;
  RECT 1641.140 6.340 1641.340 6.540 ;
  LAYER VI3 ;
  RECT 1641.140 5.940 1641.340 6.140 ;
  LAYER VI3 ;
  RECT 1640.740 6.340 1640.940 6.540 ;
  LAYER VI3 ;
  RECT 1640.740 5.940 1640.940 6.140 ;
  LAYER VI3 ;
  RECT 1640.340 6.340 1640.540 6.540 ;
  LAYER VI3 ;
  RECT 1640.340 5.940 1640.540 6.140 ;
  LAYER VI3 ;
  RECT 1639.940 6.340 1640.140 6.540 ;
  LAYER VI3 ;
  RECT 1639.940 5.940 1640.140 6.140 ;
  LAYER VI3 ;
  RECT 1639.540 6.340 1639.740 6.540 ;
  LAYER VI3 ;
  RECT 1639.540 5.940 1639.740 6.140 ;
  LAYER VI3 ;
  RECT 1639.140 6.340 1639.340 6.540 ;
  LAYER VI3 ;
  RECT 1639.140 5.940 1639.340 6.140 ;
  LAYER VI3 ;
  RECT 1638.740 6.340 1638.940 6.540 ;
  LAYER VI3 ;
  RECT 1638.740 5.940 1638.940 6.140 ;
  LAYER VI3 ;
  RECT 1638.340 6.340 1638.540 6.540 ;
  LAYER VI3 ;
  RECT 1638.340 5.940 1638.540 6.140 ;
  LAYER VI3 ;
  RECT 1637.940 6.340 1638.140 6.540 ;
  LAYER VI3 ;
  RECT 1637.940 5.940 1638.140 6.140 ;
  LAYER VI3 ;
  RECT 1637.540 6.340 1637.740 6.540 ;
  LAYER VI3 ;
  RECT 1637.540 5.940 1637.740 6.140 ;
  LAYER VI3 ;
  RECT 1637.140 6.340 1637.340 6.540 ;
  LAYER VI3 ;
  RECT 1637.140 5.940 1637.340 6.140 ;
  LAYER VI3 ;
  RECT 1636.740 6.340 1636.940 6.540 ;
  LAYER VI3 ;
  RECT 1636.740 5.940 1636.940 6.140 ;
  LAYER VI3 ;
  RECT 1636.340 6.340 1636.540 6.540 ;
  LAYER VI3 ;
  RECT 1636.340 5.940 1636.540 6.140 ;
  LAYER VI3 ;
  RECT 1635.940 6.340 1636.140 6.540 ;
  LAYER VI3 ;
  RECT 1635.940 5.940 1636.140 6.140 ;
  LAYER VI3 ;
  RECT 1635.540 6.340 1635.740 6.540 ;
  LAYER VI3 ;
  RECT 1635.540 5.940 1635.740 6.140 ;
  LAYER VI3 ;
  RECT 1656.620 5.880 1664.620 6.740 ;
  LAYER VI3 ;
  RECT 1664.220 6.340 1664.420 6.540 ;
  LAYER VI3 ;
  RECT 1664.220 5.940 1664.420 6.140 ;
  LAYER VI3 ;
  RECT 1663.820 6.340 1664.020 6.540 ;
  LAYER VI3 ;
  RECT 1663.820 5.940 1664.020 6.140 ;
  LAYER VI3 ;
  RECT 1663.420 6.340 1663.620 6.540 ;
  LAYER VI3 ;
  RECT 1663.420 5.940 1663.620 6.140 ;
  LAYER VI3 ;
  RECT 1663.020 6.340 1663.220 6.540 ;
  LAYER VI3 ;
  RECT 1663.020 5.940 1663.220 6.140 ;
  LAYER VI3 ;
  RECT 1662.620 6.340 1662.820 6.540 ;
  LAYER VI3 ;
  RECT 1662.620 5.940 1662.820 6.140 ;
  LAYER VI3 ;
  RECT 1662.220 6.340 1662.420 6.540 ;
  LAYER VI3 ;
  RECT 1662.220 5.940 1662.420 6.140 ;
  LAYER VI3 ;
  RECT 1661.820 6.340 1662.020 6.540 ;
  LAYER VI3 ;
  RECT 1661.820 5.940 1662.020 6.140 ;
  LAYER VI3 ;
  RECT 1661.420 6.340 1661.620 6.540 ;
  LAYER VI3 ;
  RECT 1661.420 5.940 1661.620 6.140 ;
  LAYER VI3 ;
  RECT 1661.020 6.340 1661.220 6.540 ;
  LAYER VI3 ;
  RECT 1661.020 5.940 1661.220 6.140 ;
  LAYER VI3 ;
  RECT 1660.620 6.340 1660.820 6.540 ;
  LAYER VI3 ;
  RECT 1660.620 5.940 1660.820 6.140 ;
  LAYER VI3 ;
  RECT 1660.220 6.340 1660.420 6.540 ;
  LAYER VI3 ;
  RECT 1660.220 5.940 1660.420 6.140 ;
  LAYER VI3 ;
  RECT 1659.820 6.340 1660.020 6.540 ;
  LAYER VI3 ;
  RECT 1659.820 5.940 1660.020 6.140 ;
  LAYER VI3 ;
  RECT 1659.420 6.340 1659.620 6.540 ;
  LAYER VI3 ;
  RECT 1659.420 5.940 1659.620 6.140 ;
  LAYER VI3 ;
  RECT 1659.020 6.340 1659.220 6.540 ;
  LAYER VI3 ;
  RECT 1659.020 5.940 1659.220 6.140 ;
  LAYER VI3 ;
  RECT 1658.620 6.340 1658.820 6.540 ;
  LAYER VI3 ;
  RECT 1658.620 5.940 1658.820 6.140 ;
  LAYER VI3 ;
  RECT 1658.220 6.340 1658.420 6.540 ;
  LAYER VI3 ;
  RECT 1658.220 5.940 1658.420 6.140 ;
  LAYER VI3 ;
  RECT 1657.820 6.340 1658.020 6.540 ;
  LAYER VI3 ;
  RECT 1657.820 5.940 1658.020 6.140 ;
  LAYER VI3 ;
  RECT 1657.420 6.340 1657.620 6.540 ;
  LAYER VI3 ;
  RECT 1657.420 5.940 1657.620 6.140 ;
  LAYER VI3 ;
  RECT 1657.020 6.340 1657.220 6.540 ;
  LAYER VI3 ;
  RECT 1657.020 5.940 1657.220 6.140 ;
  LAYER VI3 ;
  RECT 1656.620 6.340 1656.820 6.540 ;
  LAYER VI3 ;
  RECT 1656.620 5.940 1656.820 6.140 ;
  LAYER VI3 ;
  RECT 1676.460 5.880 1684.460 6.740 ;
  LAYER VI3 ;
  RECT 1684.060 6.340 1684.260 6.540 ;
  LAYER VI3 ;
  RECT 1684.060 5.940 1684.260 6.140 ;
  LAYER VI3 ;
  RECT 1683.660 6.340 1683.860 6.540 ;
  LAYER VI3 ;
  RECT 1683.660 5.940 1683.860 6.140 ;
  LAYER VI3 ;
  RECT 1683.260 6.340 1683.460 6.540 ;
  LAYER VI3 ;
  RECT 1683.260 5.940 1683.460 6.140 ;
  LAYER VI3 ;
  RECT 1682.860 6.340 1683.060 6.540 ;
  LAYER VI3 ;
  RECT 1682.860 5.940 1683.060 6.140 ;
  LAYER VI3 ;
  RECT 1682.460 6.340 1682.660 6.540 ;
  LAYER VI3 ;
  RECT 1682.460 5.940 1682.660 6.140 ;
  LAYER VI3 ;
  RECT 1682.060 6.340 1682.260 6.540 ;
  LAYER VI3 ;
  RECT 1682.060 5.940 1682.260 6.140 ;
  LAYER VI3 ;
  RECT 1681.660 6.340 1681.860 6.540 ;
  LAYER VI3 ;
  RECT 1681.660 5.940 1681.860 6.140 ;
  LAYER VI3 ;
  RECT 1681.260 6.340 1681.460 6.540 ;
  LAYER VI3 ;
  RECT 1681.260 5.940 1681.460 6.140 ;
  LAYER VI3 ;
  RECT 1680.860 6.340 1681.060 6.540 ;
  LAYER VI3 ;
  RECT 1680.860 5.940 1681.060 6.140 ;
  LAYER VI3 ;
  RECT 1680.460 6.340 1680.660 6.540 ;
  LAYER VI3 ;
  RECT 1680.460 5.940 1680.660 6.140 ;
  LAYER VI3 ;
  RECT 1680.060 6.340 1680.260 6.540 ;
  LAYER VI3 ;
  RECT 1680.060 5.940 1680.260 6.140 ;
  LAYER VI3 ;
  RECT 1679.660 6.340 1679.860 6.540 ;
  LAYER VI3 ;
  RECT 1679.660 5.940 1679.860 6.140 ;
  LAYER VI3 ;
  RECT 1679.260 6.340 1679.460 6.540 ;
  LAYER VI3 ;
  RECT 1679.260 5.940 1679.460 6.140 ;
  LAYER VI3 ;
  RECT 1678.860 6.340 1679.060 6.540 ;
  LAYER VI3 ;
  RECT 1678.860 5.940 1679.060 6.140 ;
  LAYER VI3 ;
  RECT 1678.460 6.340 1678.660 6.540 ;
  LAYER VI3 ;
  RECT 1678.460 5.940 1678.660 6.140 ;
  LAYER VI3 ;
  RECT 1678.060 6.340 1678.260 6.540 ;
  LAYER VI3 ;
  RECT 1678.060 5.940 1678.260 6.140 ;
  LAYER VI3 ;
  RECT 1677.660 6.340 1677.860 6.540 ;
  LAYER VI3 ;
  RECT 1677.660 5.940 1677.860 6.140 ;
  LAYER VI3 ;
  RECT 1677.260 6.340 1677.460 6.540 ;
  LAYER VI3 ;
  RECT 1677.260 5.940 1677.460 6.140 ;
  LAYER VI3 ;
  RECT 1676.860 6.340 1677.060 6.540 ;
  LAYER VI3 ;
  RECT 1676.860 5.940 1677.060 6.140 ;
  LAYER VI3 ;
  RECT 1676.460 6.340 1676.660 6.540 ;
  LAYER VI3 ;
  RECT 1676.460 5.940 1676.660 6.140 ;
  LAYER VI3 ;
  RECT 1697.540 5.880 1705.540 6.740 ;
  LAYER VI3 ;
  RECT 1705.140 6.340 1705.340 6.540 ;
  LAYER VI3 ;
  RECT 1705.140 5.940 1705.340 6.140 ;
  LAYER VI3 ;
  RECT 1704.740 6.340 1704.940 6.540 ;
  LAYER VI3 ;
  RECT 1704.740 5.940 1704.940 6.140 ;
  LAYER VI3 ;
  RECT 1704.340 6.340 1704.540 6.540 ;
  LAYER VI3 ;
  RECT 1704.340 5.940 1704.540 6.140 ;
  LAYER VI3 ;
  RECT 1703.940 6.340 1704.140 6.540 ;
  LAYER VI3 ;
  RECT 1703.940 5.940 1704.140 6.140 ;
  LAYER VI3 ;
  RECT 1703.540 6.340 1703.740 6.540 ;
  LAYER VI3 ;
  RECT 1703.540 5.940 1703.740 6.140 ;
  LAYER VI3 ;
  RECT 1703.140 6.340 1703.340 6.540 ;
  LAYER VI3 ;
  RECT 1703.140 5.940 1703.340 6.140 ;
  LAYER VI3 ;
  RECT 1702.740 6.340 1702.940 6.540 ;
  LAYER VI3 ;
  RECT 1702.740 5.940 1702.940 6.140 ;
  LAYER VI3 ;
  RECT 1702.340 6.340 1702.540 6.540 ;
  LAYER VI3 ;
  RECT 1702.340 5.940 1702.540 6.140 ;
  LAYER VI3 ;
  RECT 1701.940 6.340 1702.140 6.540 ;
  LAYER VI3 ;
  RECT 1701.940 5.940 1702.140 6.140 ;
  LAYER VI3 ;
  RECT 1701.540 6.340 1701.740 6.540 ;
  LAYER VI3 ;
  RECT 1701.540 5.940 1701.740 6.140 ;
  LAYER VI3 ;
  RECT 1701.140 6.340 1701.340 6.540 ;
  LAYER VI3 ;
  RECT 1701.140 5.940 1701.340 6.140 ;
  LAYER VI3 ;
  RECT 1700.740 6.340 1700.940 6.540 ;
  LAYER VI3 ;
  RECT 1700.740 5.940 1700.940 6.140 ;
  LAYER VI3 ;
  RECT 1700.340 6.340 1700.540 6.540 ;
  LAYER VI3 ;
  RECT 1700.340 5.940 1700.540 6.140 ;
  LAYER VI3 ;
  RECT 1699.940 6.340 1700.140 6.540 ;
  LAYER VI3 ;
  RECT 1699.940 5.940 1700.140 6.140 ;
  LAYER VI3 ;
  RECT 1699.540 6.340 1699.740 6.540 ;
  LAYER VI3 ;
  RECT 1699.540 5.940 1699.740 6.140 ;
  LAYER VI3 ;
  RECT 1699.140 6.340 1699.340 6.540 ;
  LAYER VI3 ;
  RECT 1699.140 5.940 1699.340 6.140 ;
  LAYER VI3 ;
  RECT 1698.740 6.340 1698.940 6.540 ;
  LAYER VI3 ;
  RECT 1698.740 5.940 1698.940 6.140 ;
  LAYER VI3 ;
  RECT 1698.340 6.340 1698.540 6.540 ;
  LAYER VI3 ;
  RECT 1698.340 5.940 1698.540 6.140 ;
  LAYER VI3 ;
  RECT 1697.940 6.340 1698.140 6.540 ;
  LAYER VI3 ;
  RECT 1697.940 5.940 1698.140 6.140 ;
  LAYER VI3 ;
  RECT 1697.540 6.340 1697.740 6.540 ;
  LAYER VI3 ;
  RECT 1697.540 5.940 1697.740 6.140 ;
  LAYER VI3 ;
  RECT 1717.380 5.880 1725.380 6.740 ;
  LAYER VI3 ;
  RECT 1724.980 6.340 1725.180 6.540 ;
  LAYER VI3 ;
  RECT 1724.980 5.940 1725.180 6.140 ;
  LAYER VI3 ;
  RECT 1724.580 6.340 1724.780 6.540 ;
  LAYER VI3 ;
  RECT 1724.580 5.940 1724.780 6.140 ;
  LAYER VI3 ;
  RECT 1724.180 6.340 1724.380 6.540 ;
  LAYER VI3 ;
  RECT 1724.180 5.940 1724.380 6.140 ;
  LAYER VI3 ;
  RECT 1723.780 6.340 1723.980 6.540 ;
  LAYER VI3 ;
  RECT 1723.780 5.940 1723.980 6.140 ;
  LAYER VI3 ;
  RECT 1723.380 6.340 1723.580 6.540 ;
  LAYER VI3 ;
  RECT 1723.380 5.940 1723.580 6.140 ;
  LAYER VI3 ;
  RECT 1722.980 6.340 1723.180 6.540 ;
  LAYER VI3 ;
  RECT 1722.980 5.940 1723.180 6.140 ;
  LAYER VI3 ;
  RECT 1722.580 6.340 1722.780 6.540 ;
  LAYER VI3 ;
  RECT 1722.580 5.940 1722.780 6.140 ;
  LAYER VI3 ;
  RECT 1722.180 6.340 1722.380 6.540 ;
  LAYER VI3 ;
  RECT 1722.180 5.940 1722.380 6.140 ;
  LAYER VI3 ;
  RECT 1721.780 6.340 1721.980 6.540 ;
  LAYER VI3 ;
  RECT 1721.780 5.940 1721.980 6.140 ;
  LAYER VI3 ;
  RECT 1721.380 6.340 1721.580 6.540 ;
  LAYER VI3 ;
  RECT 1721.380 5.940 1721.580 6.140 ;
  LAYER VI3 ;
  RECT 1720.980 6.340 1721.180 6.540 ;
  LAYER VI3 ;
  RECT 1720.980 5.940 1721.180 6.140 ;
  LAYER VI3 ;
  RECT 1720.580 6.340 1720.780 6.540 ;
  LAYER VI3 ;
  RECT 1720.580 5.940 1720.780 6.140 ;
  LAYER VI3 ;
  RECT 1720.180 6.340 1720.380 6.540 ;
  LAYER VI3 ;
  RECT 1720.180 5.940 1720.380 6.140 ;
  LAYER VI3 ;
  RECT 1719.780 6.340 1719.980 6.540 ;
  LAYER VI3 ;
  RECT 1719.780 5.940 1719.980 6.140 ;
  LAYER VI3 ;
  RECT 1719.380 6.340 1719.580 6.540 ;
  LAYER VI3 ;
  RECT 1719.380 5.940 1719.580 6.140 ;
  LAYER VI3 ;
  RECT 1718.980 6.340 1719.180 6.540 ;
  LAYER VI3 ;
  RECT 1718.980 5.940 1719.180 6.140 ;
  LAYER VI3 ;
  RECT 1718.580 6.340 1718.780 6.540 ;
  LAYER VI3 ;
  RECT 1718.580 5.940 1718.780 6.140 ;
  LAYER VI3 ;
  RECT 1718.180 6.340 1718.380 6.540 ;
  LAYER VI3 ;
  RECT 1718.180 5.940 1718.380 6.140 ;
  LAYER VI3 ;
  RECT 1717.780 6.340 1717.980 6.540 ;
  LAYER VI3 ;
  RECT 1717.780 5.940 1717.980 6.140 ;
  LAYER VI3 ;
  RECT 1717.380 6.340 1717.580 6.540 ;
  LAYER VI3 ;
  RECT 1717.380 5.940 1717.580 6.140 ;
  LAYER VI3 ;
  RECT 1738.460 5.880 1746.460 6.740 ;
  LAYER VI3 ;
  RECT 1746.060 6.340 1746.260 6.540 ;
  LAYER VI3 ;
  RECT 1746.060 5.940 1746.260 6.140 ;
  LAYER VI3 ;
  RECT 1745.660 6.340 1745.860 6.540 ;
  LAYER VI3 ;
  RECT 1745.660 5.940 1745.860 6.140 ;
  LAYER VI3 ;
  RECT 1745.260 6.340 1745.460 6.540 ;
  LAYER VI3 ;
  RECT 1745.260 5.940 1745.460 6.140 ;
  LAYER VI3 ;
  RECT 1744.860 6.340 1745.060 6.540 ;
  LAYER VI3 ;
  RECT 1744.860 5.940 1745.060 6.140 ;
  LAYER VI3 ;
  RECT 1744.460 6.340 1744.660 6.540 ;
  LAYER VI3 ;
  RECT 1744.460 5.940 1744.660 6.140 ;
  LAYER VI3 ;
  RECT 1744.060 6.340 1744.260 6.540 ;
  LAYER VI3 ;
  RECT 1744.060 5.940 1744.260 6.140 ;
  LAYER VI3 ;
  RECT 1743.660 6.340 1743.860 6.540 ;
  LAYER VI3 ;
  RECT 1743.660 5.940 1743.860 6.140 ;
  LAYER VI3 ;
  RECT 1743.260 6.340 1743.460 6.540 ;
  LAYER VI3 ;
  RECT 1743.260 5.940 1743.460 6.140 ;
  LAYER VI3 ;
  RECT 1742.860 6.340 1743.060 6.540 ;
  LAYER VI3 ;
  RECT 1742.860 5.940 1743.060 6.140 ;
  LAYER VI3 ;
  RECT 1742.460 6.340 1742.660 6.540 ;
  LAYER VI3 ;
  RECT 1742.460 5.940 1742.660 6.140 ;
  LAYER VI3 ;
  RECT 1742.060 6.340 1742.260 6.540 ;
  LAYER VI3 ;
  RECT 1742.060 5.940 1742.260 6.140 ;
  LAYER VI3 ;
  RECT 1741.660 6.340 1741.860 6.540 ;
  LAYER VI3 ;
  RECT 1741.660 5.940 1741.860 6.140 ;
  LAYER VI3 ;
  RECT 1741.260 6.340 1741.460 6.540 ;
  LAYER VI3 ;
  RECT 1741.260 5.940 1741.460 6.140 ;
  LAYER VI3 ;
  RECT 1740.860 6.340 1741.060 6.540 ;
  LAYER VI3 ;
  RECT 1740.860 5.940 1741.060 6.140 ;
  LAYER VI3 ;
  RECT 1740.460 6.340 1740.660 6.540 ;
  LAYER VI3 ;
  RECT 1740.460 5.940 1740.660 6.140 ;
  LAYER VI3 ;
  RECT 1740.060 6.340 1740.260 6.540 ;
  LAYER VI3 ;
  RECT 1740.060 5.940 1740.260 6.140 ;
  LAYER VI3 ;
  RECT 1739.660 6.340 1739.860 6.540 ;
  LAYER VI3 ;
  RECT 1739.660 5.940 1739.860 6.140 ;
  LAYER VI3 ;
  RECT 1739.260 6.340 1739.460 6.540 ;
  LAYER VI3 ;
  RECT 1739.260 5.940 1739.460 6.140 ;
  LAYER VI3 ;
  RECT 1738.860 6.340 1739.060 6.540 ;
  LAYER VI3 ;
  RECT 1738.860 5.940 1739.060 6.140 ;
  LAYER VI3 ;
  RECT 1738.460 6.340 1738.660 6.540 ;
  LAYER VI3 ;
  RECT 1738.460 5.940 1738.660 6.140 ;
  LAYER VI3 ;
  RECT 1758.300 5.880 1766.300 6.740 ;
  LAYER VI3 ;
  RECT 1765.900 6.340 1766.100 6.540 ;
  LAYER VI3 ;
  RECT 1765.900 5.940 1766.100 6.140 ;
  LAYER VI3 ;
  RECT 1765.500 6.340 1765.700 6.540 ;
  LAYER VI3 ;
  RECT 1765.500 5.940 1765.700 6.140 ;
  LAYER VI3 ;
  RECT 1765.100 6.340 1765.300 6.540 ;
  LAYER VI3 ;
  RECT 1765.100 5.940 1765.300 6.140 ;
  LAYER VI3 ;
  RECT 1764.700 6.340 1764.900 6.540 ;
  LAYER VI3 ;
  RECT 1764.700 5.940 1764.900 6.140 ;
  LAYER VI3 ;
  RECT 1764.300 6.340 1764.500 6.540 ;
  LAYER VI3 ;
  RECT 1764.300 5.940 1764.500 6.140 ;
  LAYER VI3 ;
  RECT 1763.900 6.340 1764.100 6.540 ;
  LAYER VI3 ;
  RECT 1763.900 5.940 1764.100 6.140 ;
  LAYER VI3 ;
  RECT 1763.500 6.340 1763.700 6.540 ;
  LAYER VI3 ;
  RECT 1763.500 5.940 1763.700 6.140 ;
  LAYER VI3 ;
  RECT 1763.100 6.340 1763.300 6.540 ;
  LAYER VI3 ;
  RECT 1763.100 5.940 1763.300 6.140 ;
  LAYER VI3 ;
  RECT 1762.700 6.340 1762.900 6.540 ;
  LAYER VI3 ;
  RECT 1762.700 5.940 1762.900 6.140 ;
  LAYER VI3 ;
  RECT 1762.300 6.340 1762.500 6.540 ;
  LAYER VI3 ;
  RECT 1762.300 5.940 1762.500 6.140 ;
  LAYER VI3 ;
  RECT 1761.900 6.340 1762.100 6.540 ;
  LAYER VI3 ;
  RECT 1761.900 5.940 1762.100 6.140 ;
  LAYER VI3 ;
  RECT 1761.500 6.340 1761.700 6.540 ;
  LAYER VI3 ;
  RECT 1761.500 5.940 1761.700 6.140 ;
  LAYER VI3 ;
  RECT 1761.100 6.340 1761.300 6.540 ;
  LAYER VI3 ;
  RECT 1761.100 5.940 1761.300 6.140 ;
  LAYER VI3 ;
  RECT 1760.700 6.340 1760.900 6.540 ;
  LAYER VI3 ;
  RECT 1760.700 5.940 1760.900 6.140 ;
  LAYER VI3 ;
  RECT 1760.300 6.340 1760.500 6.540 ;
  LAYER VI3 ;
  RECT 1760.300 5.940 1760.500 6.140 ;
  LAYER VI3 ;
  RECT 1759.900 6.340 1760.100 6.540 ;
  LAYER VI3 ;
  RECT 1759.900 5.940 1760.100 6.140 ;
  LAYER VI3 ;
  RECT 1759.500 6.340 1759.700 6.540 ;
  LAYER VI3 ;
  RECT 1759.500 5.940 1759.700 6.140 ;
  LAYER VI3 ;
  RECT 1759.100 6.340 1759.300 6.540 ;
  LAYER VI3 ;
  RECT 1759.100 5.940 1759.300 6.140 ;
  LAYER VI3 ;
  RECT 1758.700 6.340 1758.900 6.540 ;
  LAYER VI3 ;
  RECT 1758.700 5.940 1758.900 6.140 ;
  LAYER VI3 ;
  RECT 1758.300 6.340 1758.500 6.540 ;
  LAYER VI3 ;
  RECT 1758.300 5.940 1758.500 6.140 ;
  LAYER VI3 ;
  RECT 1779.380 5.880 1787.380 6.740 ;
  LAYER VI3 ;
  RECT 1786.980 6.340 1787.180 6.540 ;
  LAYER VI3 ;
  RECT 1786.980 5.940 1787.180 6.140 ;
  LAYER VI3 ;
  RECT 1786.580 6.340 1786.780 6.540 ;
  LAYER VI3 ;
  RECT 1786.580 5.940 1786.780 6.140 ;
  LAYER VI3 ;
  RECT 1786.180 6.340 1786.380 6.540 ;
  LAYER VI3 ;
  RECT 1786.180 5.940 1786.380 6.140 ;
  LAYER VI3 ;
  RECT 1785.780 6.340 1785.980 6.540 ;
  LAYER VI3 ;
  RECT 1785.780 5.940 1785.980 6.140 ;
  LAYER VI3 ;
  RECT 1785.380 6.340 1785.580 6.540 ;
  LAYER VI3 ;
  RECT 1785.380 5.940 1785.580 6.140 ;
  LAYER VI3 ;
  RECT 1784.980 6.340 1785.180 6.540 ;
  LAYER VI3 ;
  RECT 1784.980 5.940 1785.180 6.140 ;
  LAYER VI3 ;
  RECT 1784.580 6.340 1784.780 6.540 ;
  LAYER VI3 ;
  RECT 1784.580 5.940 1784.780 6.140 ;
  LAYER VI3 ;
  RECT 1784.180 6.340 1784.380 6.540 ;
  LAYER VI3 ;
  RECT 1784.180 5.940 1784.380 6.140 ;
  LAYER VI3 ;
  RECT 1783.780 6.340 1783.980 6.540 ;
  LAYER VI3 ;
  RECT 1783.780 5.940 1783.980 6.140 ;
  LAYER VI3 ;
  RECT 1783.380 6.340 1783.580 6.540 ;
  LAYER VI3 ;
  RECT 1783.380 5.940 1783.580 6.140 ;
  LAYER VI3 ;
  RECT 1782.980 6.340 1783.180 6.540 ;
  LAYER VI3 ;
  RECT 1782.980 5.940 1783.180 6.140 ;
  LAYER VI3 ;
  RECT 1782.580 6.340 1782.780 6.540 ;
  LAYER VI3 ;
  RECT 1782.580 5.940 1782.780 6.140 ;
  LAYER VI3 ;
  RECT 1782.180 6.340 1782.380 6.540 ;
  LAYER VI3 ;
  RECT 1782.180 5.940 1782.380 6.140 ;
  LAYER VI3 ;
  RECT 1781.780 6.340 1781.980 6.540 ;
  LAYER VI3 ;
  RECT 1781.780 5.940 1781.980 6.140 ;
  LAYER VI3 ;
  RECT 1781.380 6.340 1781.580 6.540 ;
  LAYER VI3 ;
  RECT 1781.380 5.940 1781.580 6.140 ;
  LAYER VI3 ;
  RECT 1780.980 6.340 1781.180 6.540 ;
  LAYER VI3 ;
  RECT 1780.980 5.940 1781.180 6.140 ;
  LAYER VI3 ;
  RECT 1780.580 6.340 1780.780 6.540 ;
  LAYER VI3 ;
  RECT 1780.580 5.940 1780.780 6.140 ;
  LAYER VI3 ;
  RECT 1780.180 6.340 1780.380 6.540 ;
  LAYER VI3 ;
  RECT 1780.180 5.940 1780.380 6.140 ;
  LAYER VI3 ;
  RECT 1779.780 6.340 1779.980 6.540 ;
  LAYER VI3 ;
  RECT 1779.780 5.940 1779.980 6.140 ;
  LAYER VI3 ;
  RECT 1779.380 6.340 1779.580 6.540 ;
  LAYER VI3 ;
  RECT 1779.380 5.940 1779.580 6.140 ;
  LAYER VI3 ;
  RECT 1799.220 5.880 1807.220 6.740 ;
  LAYER VI3 ;
  RECT 1806.820 6.340 1807.020 6.540 ;
  LAYER VI3 ;
  RECT 1806.820 5.940 1807.020 6.140 ;
  LAYER VI3 ;
  RECT 1806.420 6.340 1806.620 6.540 ;
  LAYER VI3 ;
  RECT 1806.420 5.940 1806.620 6.140 ;
  LAYER VI3 ;
  RECT 1806.020 6.340 1806.220 6.540 ;
  LAYER VI3 ;
  RECT 1806.020 5.940 1806.220 6.140 ;
  LAYER VI3 ;
  RECT 1805.620 6.340 1805.820 6.540 ;
  LAYER VI3 ;
  RECT 1805.620 5.940 1805.820 6.140 ;
  LAYER VI3 ;
  RECT 1805.220 6.340 1805.420 6.540 ;
  LAYER VI3 ;
  RECT 1805.220 5.940 1805.420 6.140 ;
  LAYER VI3 ;
  RECT 1804.820 6.340 1805.020 6.540 ;
  LAYER VI3 ;
  RECT 1804.820 5.940 1805.020 6.140 ;
  LAYER VI3 ;
  RECT 1804.420 6.340 1804.620 6.540 ;
  LAYER VI3 ;
  RECT 1804.420 5.940 1804.620 6.140 ;
  LAYER VI3 ;
  RECT 1804.020 6.340 1804.220 6.540 ;
  LAYER VI3 ;
  RECT 1804.020 5.940 1804.220 6.140 ;
  LAYER VI3 ;
  RECT 1803.620 6.340 1803.820 6.540 ;
  LAYER VI3 ;
  RECT 1803.620 5.940 1803.820 6.140 ;
  LAYER VI3 ;
  RECT 1803.220 6.340 1803.420 6.540 ;
  LAYER VI3 ;
  RECT 1803.220 5.940 1803.420 6.140 ;
  LAYER VI3 ;
  RECT 1802.820 6.340 1803.020 6.540 ;
  LAYER VI3 ;
  RECT 1802.820 5.940 1803.020 6.140 ;
  LAYER VI3 ;
  RECT 1802.420 6.340 1802.620 6.540 ;
  LAYER VI3 ;
  RECT 1802.420 5.940 1802.620 6.140 ;
  LAYER VI3 ;
  RECT 1802.020 6.340 1802.220 6.540 ;
  LAYER VI3 ;
  RECT 1802.020 5.940 1802.220 6.140 ;
  LAYER VI3 ;
  RECT 1801.620 6.340 1801.820 6.540 ;
  LAYER VI3 ;
  RECT 1801.620 5.940 1801.820 6.140 ;
  LAYER VI3 ;
  RECT 1801.220 6.340 1801.420 6.540 ;
  LAYER VI3 ;
  RECT 1801.220 5.940 1801.420 6.140 ;
  LAYER VI3 ;
  RECT 1800.820 6.340 1801.020 6.540 ;
  LAYER VI3 ;
  RECT 1800.820 5.940 1801.020 6.140 ;
  LAYER VI3 ;
  RECT 1800.420 6.340 1800.620 6.540 ;
  LAYER VI3 ;
  RECT 1800.420 5.940 1800.620 6.140 ;
  LAYER VI3 ;
  RECT 1800.020 6.340 1800.220 6.540 ;
  LAYER VI3 ;
  RECT 1800.020 5.940 1800.220 6.140 ;
  LAYER VI3 ;
  RECT 1799.620 6.340 1799.820 6.540 ;
  LAYER VI3 ;
  RECT 1799.620 5.940 1799.820 6.140 ;
  LAYER VI3 ;
  RECT 1799.220 6.340 1799.420 6.540 ;
  LAYER VI3 ;
  RECT 1799.220 5.940 1799.420 6.140 ;
  LAYER VI3 ;
  RECT 1820.300 5.880 1828.300 6.740 ;
  LAYER VI3 ;
  RECT 1827.900 6.340 1828.100 6.540 ;
  LAYER VI3 ;
  RECT 1827.900 5.940 1828.100 6.140 ;
  LAYER VI3 ;
  RECT 1827.500 6.340 1827.700 6.540 ;
  LAYER VI3 ;
  RECT 1827.500 5.940 1827.700 6.140 ;
  LAYER VI3 ;
  RECT 1827.100 6.340 1827.300 6.540 ;
  LAYER VI3 ;
  RECT 1827.100 5.940 1827.300 6.140 ;
  LAYER VI3 ;
  RECT 1826.700 6.340 1826.900 6.540 ;
  LAYER VI3 ;
  RECT 1826.700 5.940 1826.900 6.140 ;
  LAYER VI3 ;
  RECT 1826.300 6.340 1826.500 6.540 ;
  LAYER VI3 ;
  RECT 1826.300 5.940 1826.500 6.140 ;
  LAYER VI3 ;
  RECT 1825.900 6.340 1826.100 6.540 ;
  LAYER VI3 ;
  RECT 1825.900 5.940 1826.100 6.140 ;
  LAYER VI3 ;
  RECT 1825.500 6.340 1825.700 6.540 ;
  LAYER VI3 ;
  RECT 1825.500 5.940 1825.700 6.140 ;
  LAYER VI3 ;
  RECT 1825.100 6.340 1825.300 6.540 ;
  LAYER VI3 ;
  RECT 1825.100 5.940 1825.300 6.140 ;
  LAYER VI3 ;
  RECT 1824.700 6.340 1824.900 6.540 ;
  LAYER VI3 ;
  RECT 1824.700 5.940 1824.900 6.140 ;
  LAYER VI3 ;
  RECT 1824.300 6.340 1824.500 6.540 ;
  LAYER VI3 ;
  RECT 1824.300 5.940 1824.500 6.140 ;
  LAYER VI3 ;
  RECT 1823.900 6.340 1824.100 6.540 ;
  LAYER VI3 ;
  RECT 1823.900 5.940 1824.100 6.140 ;
  LAYER VI3 ;
  RECT 1823.500 6.340 1823.700 6.540 ;
  LAYER VI3 ;
  RECT 1823.500 5.940 1823.700 6.140 ;
  LAYER VI3 ;
  RECT 1823.100 6.340 1823.300 6.540 ;
  LAYER VI3 ;
  RECT 1823.100 5.940 1823.300 6.140 ;
  LAYER VI3 ;
  RECT 1822.700 6.340 1822.900 6.540 ;
  LAYER VI3 ;
  RECT 1822.700 5.940 1822.900 6.140 ;
  LAYER VI3 ;
  RECT 1822.300 6.340 1822.500 6.540 ;
  LAYER VI3 ;
  RECT 1822.300 5.940 1822.500 6.140 ;
  LAYER VI3 ;
  RECT 1821.900 6.340 1822.100 6.540 ;
  LAYER VI3 ;
  RECT 1821.900 5.940 1822.100 6.140 ;
  LAYER VI3 ;
  RECT 1821.500 6.340 1821.700 6.540 ;
  LAYER VI3 ;
  RECT 1821.500 5.940 1821.700 6.140 ;
  LAYER VI3 ;
  RECT 1821.100 6.340 1821.300 6.540 ;
  LAYER VI3 ;
  RECT 1821.100 5.940 1821.300 6.140 ;
  LAYER VI3 ;
  RECT 1820.700 6.340 1820.900 6.540 ;
  LAYER VI3 ;
  RECT 1820.700 5.940 1820.900 6.140 ;
  LAYER VI3 ;
  RECT 1820.300 6.340 1820.500 6.540 ;
  LAYER VI3 ;
  RECT 1820.300 5.940 1820.500 6.140 ;
  LAYER VI3 ;
  RECT 1840.140 5.880 1848.140 6.740 ;
  LAYER VI3 ;
  RECT 1847.740 6.340 1847.940 6.540 ;
  LAYER VI3 ;
  RECT 1847.740 5.940 1847.940 6.140 ;
  LAYER VI3 ;
  RECT 1847.340 6.340 1847.540 6.540 ;
  LAYER VI3 ;
  RECT 1847.340 5.940 1847.540 6.140 ;
  LAYER VI3 ;
  RECT 1846.940 6.340 1847.140 6.540 ;
  LAYER VI3 ;
  RECT 1846.940 5.940 1847.140 6.140 ;
  LAYER VI3 ;
  RECT 1846.540 6.340 1846.740 6.540 ;
  LAYER VI3 ;
  RECT 1846.540 5.940 1846.740 6.140 ;
  LAYER VI3 ;
  RECT 1846.140 6.340 1846.340 6.540 ;
  LAYER VI3 ;
  RECT 1846.140 5.940 1846.340 6.140 ;
  LAYER VI3 ;
  RECT 1845.740 6.340 1845.940 6.540 ;
  LAYER VI3 ;
  RECT 1845.740 5.940 1845.940 6.140 ;
  LAYER VI3 ;
  RECT 1845.340 6.340 1845.540 6.540 ;
  LAYER VI3 ;
  RECT 1845.340 5.940 1845.540 6.140 ;
  LAYER VI3 ;
  RECT 1844.940 6.340 1845.140 6.540 ;
  LAYER VI3 ;
  RECT 1844.940 5.940 1845.140 6.140 ;
  LAYER VI3 ;
  RECT 1844.540 6.340 1844.740 6.540 ;
  LAYER VI3 ;
  RECT 1844.540 5.940 1844.740 6.140 ;
  LAYER VI3 ;
  RECT 1844.140 6.340 1844.340 6.540 ;
  LAYER VI3 ;
  RECT 1844.140 5.940 1844.340 6.140 ;
  LAYER VI3 ;
  RECT 1843.740 6.340 1843.940 6.540 ;
  LAYER VI3 ;
  RECT 1843.740 5.940 1843.940 6.140 ;
  LAYER VI3 ;
  RECT 1843.340 6.340 1843.540 6.540 ;
  LAYER VI3 ;
  RECT 1843.340 5.940 1843.540 6.140 ;
  LAYER VI3 ;
  RECT 1842.940 6.340 1843.140 6.540 ;
  LAYER VI3 ;
  RECT 1842.940 5.940 1843.140 6.140 ;
  LAYER VI3 ;
  RECT 1842.540 6.340 1842.740 6.540 ;
  LAYER VI3 ;
  RECT 1842.540 5.940 1842.740 6.140 ;
  LAYER VI3 ;
  RECT 1842.140 6.340 1842.340 6.540 ;
  LAYER VI3 ;
  RECT 1842.140 5.940 1842.340 6.140 ;
  LAYER VI3 ;
  RECT 1841.740 6.340 1841.940 6.540 ;
  LAYER VI3 ;
  RECT 1841.740 5.940 1841.940 6.140 ;
  LAYER VI3 ;
  RECT 1841.340 6.340 1841.540 6.540 ;
  LAYER VI3 ;
  RECT 1841.340 5.940 1841.540 6.140 ;
  LAYER VI3 ;
  RECT 1840.940 6.340 1841.140 6.540 ;
  LAYER VI3 ;
  RECT 1840.940 5.940 1841.140 6.140 ;
  LAYER VI3 ;
  RECT 1840.540 6.340 1840.740 6.540 ;
  LAYER VI3 ;
  RECT 1840.540 5.940 1840.740 6.140 ;
  LAYER VI3 ;
  RECT 1840.140 6.340 1840.340 6.540 ;
  LAYER VI3 ;
  RECT 1840.140 5.940 1840.340 6.140 ;
  LAYER VI3 ;
  RECT 1861.220 5.880 1869.220 6.740 ;
  LAYER VI3 ;
  RECT 1868.820 6.340 1869.020 6.540 ;
  LAYER VI3 ;
  RECT 1868.820 5.940 1869.020 6.140 ;
  LAYER VI3 ;
  RECT 1868.420 6.340 1868.620 6.540 ;
  LAYER VI3 ;
  RECT 1868.420 5.940 1868.620 6.140 ;
  LAYER VI3 ;
  RECT 1868.020 6.340 1868.220 6.540 ;
  LAYER VI3 ;
  RECT 1868.020 5.940 1868.220 6.140 ;
  LAYER VI3 ;
  RECT 1867.620 6.340 1867.820 6.540 ;
  LAYER VI3 ;
  RECT 1867.620 5.940 1867.820 6.140 ;
  LAYER VI3 ;
  RECT 1867.220 6.340 1867.420 6.540 ;
  LAYER VI3 ;
  RECT 1867.220 5.940 1867.420 6.140 ;
  LAYER VI3 ;
  RECT 1866.820 6.340 1867.020 6.540 ;
  LAYER VI3 ;
  RECT 1866.820 5.940 1867.020 6.140 ;
  LAYER VI3 ;
  RECT 1866.420 6.340 1866.620 6.540 ;
  LAYER VI3 ;
  RECT 1866.420 5.940 1866.620 6.140 ;
  LAYER VI3 ;
  RECT 1866.020 6.340 1866.220 6.540 ;
  LAYER VI3 ;
  RECT 1866.020 5.940 1866.220 6.140 ;
  LAYER VI3 ;
  RECT 1865.620 6.340 1865.820 6.540 ;
  LAYER VI3 ;
  RECT 1865.620 5.940 1865.820 6.140 ;
  LAYER VI3 ;
  RECT 1865.220 6.340 1865.420 6.540 ;
  LAYER VI3 ;
  RECT 1865.220 5.940 1865.420 6.140 ;
  LAYER VI3 ;
  RECT 1864.820 6.340 1865.020 6.540 ;
  LAYER VI3 ;
  RECT 1864.820 5.940 1865.020 6.140 ;
  LAYER VI3 ;
  RECT 1864.420 6.340 1864.620 6.540 ;
  LAYER VI3 ;
  RECT 1864.420 5.940 1864.620 6.140 ;
  LAYER VI3 ;
  RECT 1864.020 6.340 1864.220 6.540 ;
  LAYER VI3 ;
  RECT 1864.020 5.940 1864.220 6.140 ;
  LAYER VI3 ;
  RECT 1863.620 6.340 1863.820 6.540 ;
  LAYER VI3 ;
  RECT 1863.620 5.940 1863.820 6.140 ;
  LAYER VI3 ;
  RECT 1863.220 6.340 1863.420 6.540 ;
  LAYER VI3 ;
  RECT 1863.220 5.940 1863.420 6.140 ;
  LAYER VI3 ;
  RECT 1862.820 6.340 1863.020 6.540 ;
  LAYER VI3 ;
  RECT 1862.820 5.940 1863.020 6.140 ;
  LAYER VI3 ;
  RECT 1862.420 6.340 1862.620 6.540 ;
  LAYER VI3 ;
  RECT 1862.420 5.940 1862.620 6.140 ;
  LAYER VI3 ;
  RECT 1862.020 6.340 1862.220 6.540 ;
  LAYER VI3 ;
  RECT 1862.020 5.940 1862.220 6.140 ;
  LAYER VI3 ;
  RECT 1861.620 6.340 1861.820 6.540 ;
  LAYER VI3 ;
  RECT 1861.620 5.940 1861.820 6.140 ;
  LAYER VI3 ;
  RECT 1861.220 6.340 1861.420 6.540 ;
  LAYER VI3 ;
  RECT 1861.220 5.940 1861.420 6.140 ;
  LAYER VI3 ;
  RECT 1881.060 5.880 1889.060 6.740 ;
  LAYER VI3 ;
  RECT 1888.660 6.340 1888.860 6.540 ;
  LAYER VI3 ;
  RECT 1888.660 5.940 1888.860 6.140 ;
  LAYER VI3 ;
  RECT 1888.260 6.340 1888.460 6.540 ;
  LAYER VI3 ;
  RECT 1888.260 5.940 1888.460 6.140 ;
  LAYER VI3 ;
  RECT 1887.860 6.340 1888.060 6.540 ;
  LAYER VI3 ;
  RECT 1887.860 5.940 1888.060 6.140 ;
  LAYER VI3 ;
  RECT 1887.460 6.340 1887.660 6.540 ;
  LAYER VI3 ;
  RECT 1887.460 5.940 1887.660 6.140 ;
  LAYER VI3 ;
  RECT 1887.060 6.340 1887.260 6.540 ;
  LAYER VI3 ;
  RECT 1887.060 5.940 1887.260 6.140 ;
  LAYER VI3 ;
  RECT 1886.660 6.340 1886.860 6.540 ;
  LAYER VI3 ;
  RECT 1886.660 5.940 1886.860 6.140 ;
  LAYER VI3 ;
  RECT 1886.260 6.340 1886.460 6.540 ;
  LAYER VI3 ;
  RECT 1886.260 5.940 1886.460 6.140 ;
  LAYER VI3 ;
  RECT 1885.860 6.340 1886.060 6.540 ;
  LAYER VI3 ;
  RECT 1885.860 5.940 1886.060 6.140 ;
  LAYER VI3 ;
  RECT 1885.460 6.340 1885.660 6.540 ;
  LAYER VI3 ;
  RECT 1885.460 5.940 1885.660 6.140 ;
  LAYER VI3 ;
  RECT 1885.060 6.340 1885.260 6.540 ;
  LAYER VI3 ;
  RECT 1885.060 5.940 1885.260 6.140 ;
  LAYER VI3 ;
  RECT 1884.660 6.340 1884.860 6.540 ;
  LAYER VI3 ;
  RECT 1884.660 5.940 1884.860 6.140 ;
  LAYER VI3 ;
  RECT 1884.260 6.340 1884.460 6.540 ;
  LAYER VI3 ;
  RECT 1884.260 5.940 1884.460 6.140 ;
  LAYER VI3 ;
  RECT 1883.860 6.340 1884.060 6.540 ;
  LAYER VI3 ;
  RECT 1883.860 5.940 1884.060 6.140 ;
  LAYER VI3 ;
  RECT 1883.460 6.340 1883.660 6.540 ;
  LAYER VI3 ;
  RECT 1883.460 5.940 1883.660 6.140 ;
  LAYER VI3 ;
  RECT 1883.060 6.340 1883.260 6.540 ;
  LAYER VI3 ;
  RECT 1883.060 5.940 1883.260 6.140 ;
  LAYER VI3 ;
  RECT 1882.660 6.340 1882.860 6.540 ;
  LAYER VI3 ;
  RECT 1882.660 5.940 1882.860 6.140 ;
  LAYER VI3 ;
  RECT 1882.260 6.340 1882.460 6.540 ;
  LAYER VI3 ;
  RECT 1882.260 5.940 1882.460 6.140 ;
  LAYER VI3 ;
  RECT 1881.860 6.340 1882.060 6.540 ;
  LAYER VI3 ;
  RECT 1881.860 5.940 1882.060 6.140 ;
  LAYER VI3 ;
  RECT 1881.460 6.340 1881.660 6.540 ;
  LAYER VI3 ;
  RECT 1881.460 5.940 1881.660 6.140 ;
  LAYER VI3 ;
  RECT 1881.060 6.340 1881.260 6.540 ;
  LAYER VI3 ;
  RECT 1881.060 5.940 1881.260 6.140 ;
  LAYER VI3 ;
  RECT 1902.140 5.880 1910.140 6.740 ;
  LAYER VI3 ;
  RECT 1909.740 6.340 1909.940 6.540 ;
  LAYER VI3 ;
  RECT 1909.740 5.940 1909.940 6.140 ;
  LAYER VI3 ;
  RECT 1909.340 6.340 1909.540 6.540 ;
  LAYER VI3 ;
  RECT 1909.340 5.940 1909.540 6.140 ;
  LAYER VI3 ;
  RECT 1908.940 6.340 1909.140 6.540 ;
  LAYER VI3 ;
  RECT 1908.940 5.940 1909.140 6.140 ;
  LAYER VI3 ;
  RECT 1908.540 6.340 1908.740 6.540 ;
  LAYER VI3 ;
  RECT 1908.540 5.940 1908.740 6.140 ;
  LAYER VI3 ;
  RECT 1908.140 6.340 1908.340 6.540 ;
  LAYER VI3 ;
  RECT 1908.140 5.940 1908.340 6.140 ;
  LAYER VI3 ;
  RECT 1907.740 6.340 1907.940 6.540 ;
  LAYER VI3 ;
  RECT 1907.740 5.940 1907.940 6.140 ;
  LAYER VI3 ;
  RECT 1907.340 6.340 1907.540 6.540 ;
  LAYER VI3 ;
  RECT 1907.340 5.940 1907.540 6.140 ;
  LAYER VI3 ;
  RECT 1906.940 6.340 1907.140 6.540 ;
  LAYER VI3 ;
  RECT 1906.940 5.940 1907.140 6.140 ;
  LAYER VI3 ;
  RECT 1906.540 6.340 1906.740 6.540 ;
  LAYER VI3 ;
  RECT 1906.540 5.940 1906.740 6.140 ;
  LAYER VI3 ;
  RECT 1906.140 6.340 1906.340 6.540 ;
  LAYER VI3 ;
  RECT 1906.140 5.940 1906.340 6.140 ;
  LAYER VI3 ;
  RECT 1905.740 6.340 1905.940 6.540 ;
  LAYER VI3 ;
  RECT 1905.740 5.940 1905.940 6.140 ;
  LAYER VI3 ;
  RECT 1905.340 6.340 1905.540 6.540 ;
  LAYER VI3 ;
  RECT 1905.340 5.940 1905.540 6.140 ;
  LAYER VI3 ;
  RECT 1904.940 6.340 1905.140 6.540 ;
  LAYER VI3 ;
  RECT 1904.940 5.940 1905.140 6.140 ;
  LAYER VI3 ;
  RECT 1904.540 6.340 1904.740 6.540 ;
  LAYER VI3 ;
  RECT 1904.540 5.940 1904.740 6.140 ;
  LAYER VI3 ;
  RECT 1904.140 6.340 1904.340 6.540 ;
  LAYER VI3 ;
  RECT 1904.140 5.940 1904.340 6.140 ;
  LAYER VI3 ;
  RECT 1903.740 6.340 1903.940 6.540 ;
  LAYER VI3 ;
  RECT 1903.740 5.940 1903.940 6.140 ;
  LAYER VI3 ;
  RECT 1903.340 6.340 1903.540 6.540 ;
  LAYER VI3 ;
  RECT 1903.340 5.940 1903.540 6.140 ;
  LAYER VI3 ;
  RECT 1902.940 6.340 1903.140 6.540 ;
  LAYER VI3 ;
  RECT 1902.940 5.940 1903.140 6.140 ;
  LAYER VI3 ;
  RECT 1902.540 6.340 1902.740 6.540 ;
  LAYER VI3 ;
  RECT 1902.540 5.940 1902.740 6.140 ;
  LAYER VI3 ;
  RECT 1902.140 6.340 1902.340 6.540 ;
  LAYER VI3 ;
  RECT 1902.140 5.940 1902.340 6.140 ;
  LAYER VI3 ;
  RECT 1921.980 5.880 1929.980 6.740 ;
  LAYER VI3 ;
  RECT 1929.580 6.340 1929.780 6.540 ;
  LAYER VI3 ;
  RECT 1929.580 5.940 1929.780 6.140 ;
  LAYER VI3 ;
  RECT 1929.180 6.340 1929.380 6.540 ;
  LAYER VI3 ;
  RECT 1929.180 5.940 1929.380 6.140 ;
  LAYER VI3 ;
  RECT 1928.780 6.340 1928.980 6.540 ;
  LAYER VI3 ;
  RECT 1928.780 5.940 1928.980 6.140 ;
  LAYER VI3 ;
  RECT 1928.380 6.340 1928.580 6.540 ;
  LAYER VI3 ;
  RECT 1928.380 5.940 1928.580 6.140 ;
  LAYER VI3 ;
  RECT 1927.980 6.340 1928.180 6.540 ;
  LAYER VI3 ;
  RECT 1927.980 5.940 1928.180 6.140 ;
  LAYER VI3 ;
  RECT 1927.580 6.340 1927.780 6.540 ;
  LAYER VI3 ;
  RECT 1927.580 5.940 1927.780 6.140 ;
  LAYER VI3 ;
  RECT 1927.180 6.340 1927.380 6.540 ;
  LAYER VI3 ;
  RECT 1927.180 5.940 1927.380 6.140 ;
  LAYER VI3 ;
  RECT 1926.780 6.340 1926.980 6.540 ;
  LAYER VI3 ;
  RECT 1926.780 5.940 1926.980 6.140 ;
  LAYER VI3 ;
  RECT 1926.380 6.340 1926.580 6.540 ;
  LAYER VI3 ;
  RECT 1926.380 5.940 1926.580 6.140 ;
  LAYER VI3 ;
  RECT 1925.980 6.340 1926.180 6.540 ;
  LAYER VI3 ;
  RECT 1925.980 5.940 1926.180 6.140 ;
  LAYER VI3 ;
  RECT 1925.580 6.340 1925.780 6.540 ;
  LAYER VI3 ;
  RECT 1925.580 5.940 1925.780 6.140 ;
  LAYER VI3 ;
  RECT 1925.180 6.340 1925.380 6.540 ;
  LAYER VI3 ;
  RECT 1925.180 5.940 1925.380 6.140 ;
  LAYER VI3 ;
  RECT 1924.780 6.340 1924.980 6.540 ;
  LAYER VI3 ;
  RECT 1924.780 5.940 1924.980 6.140 ;
  LAYER VI3 ;
  RECT 1924.380 6.340 1924.580 6.540 ;
  LAYER VI3 ;
  RECT 1924.380 5.940 1924.580 6.140 ;
  LAYER VI3 ;
  RECT 1923.980 6.340 1924.180 6.540 ;
  LAYER VI3 ;
  RECT 1923.980 5.940 1924.180 6.140 ;
  LAYER VI3 ;
  RECT 1923.580 6.340 1923.780 6.540 ;
  LAYER VI3 ;
  RECT 1923.580 5.940 1923.780 6.140 ;
  LAYER VI3 ;
  RECT 1923.180 6.340 1923.380 6.540 ;
  LAYER VI3 ;
  RECT 1923.180 5.940 1923.380 6.140 ;
  LAYER VI3 ;
  RECT 1922.780 6.340 1922.980 6.540 ;
  LAYER VI3 ;
  RECT 1922.780 5.940 1922.980 6.140 ;
  LAYER VI3 ;
  RECT 1922.380 6.340 1922.580 6.540 ;
  LAYER VI3 ;
  RECT 1922.380 5.940 1922.580 6.140 ;
  LAYER VI3 ;
  RECT 1921.980 6.340 1922.180 6.540 ;
  LAYER VI3 ;
  RECT 1921.980 5.940 1922.180 6.140 ;
  LAYER VI3 ;
  RECT 1943.060 5.880 1951.060 6.740 ;
  LAYER VI3 ;
  RECT 1950.660 6.340 1950.860 6.540 ;
  LAYER VI3 ;
  RECT 1950.660 5.940 1950.860 6.140 ;
  LAYER VI3 ;
  RECT 1950.260 6.340 1950.460 6.540 ;
  LAYER VI3 ;
  RECT 1950.260 5.940 1950.460 6.140 ;
  LAYER VI3 ;
  RECT 1949.860 6.340 1950.060 6.540 ;
  LAYER VI3 ;
  RECT 1949.860 5.940 1950.060 6.140 ;
  LAYER VI3 ;
  RECT 1949.460 6.340 1949.660 6.540 ;
  LAYER VI3 ;
  RECT 1949.460 5.940 1949.660 6.140 ;
  LAYER VI3 ;
  RECT 1949.060 6.340 1949.260 6.540 ;
  LAYER VI3 ;
  RECT 1949.060 5.940 1949.260 6.140 ;
  LAYER VI3 ;
  RECT 1948.660 6.340 1948.860 6.540 ;
  LAYER VI3 ;
  RECT 1948.660 5.940 1948.860 6.140 ;
  LAYER VI3 ;
  RECT 1948.260 6.340 1948.460 6.540 ;
  LAYER VI3 ;
  RECT 1948.260 5.940 1948.460 6.140 ;
  LAYER VI3 ;
  RECT 1947.860 6.340 1948.060 6.540 ;
  LAYER VI3 ;
  RECT 1947.860 5.940 1948.060 6.140 ;
  LAYER VI3 ;
  RECT 1947.460 6.340 1947.660 6.540 ;
  LAYER VI3 ;
  RECT 1947.460 5.940 1947.660 6.140 ;
  LAYER VI3 ;
  RECT 1947.060 6.340 1947.260 6.540 ;
  LAYER VI3 ;
  RECT 1947.060 5.940 1947.260 6.140 ;
  LAYER VI3 ;
  RECT 1946.660 6.340 1946.860 6.540 ;
  LAYER VI3 ;
  RECT 1946.660 5.940 1946.860 6.140 ;
  LAYER VI3 ;
  RECT 1946.260 6.340 1946.460 6.540 ;
  LAYER VI3 ;
  RECT 1946.260 5.940 1946.460 6.140 ;
  LAYER VI3 ;
  RECT 1945.860 6.340 1946.060 6.540 ;
  LAYER VI3 ;
  RECT 1945.860 5.940 1946.060 6.140 ;
  LAYER VI3 ;
  RECT 1945.460 6.340 1945.660 6.540 ;
  LAYER VI3 ;
  RECT 1945.460 5.940 1945.660 6.140 ;
  LAYER VI3 ;
  RECT 1945.060 6.340 1945.260 6.540 ;
  LAYER VI3 ;
  RECT 1945.060 5.940 1945.260 6.140 ;
  LAYER VI3 ;
  RECT 1944.660 6.340 1944.860 6.540 ;
  LAYER VI3 ;
  RECT 1944.660 5.940 1944.860 6.140 ;
  LAYER VI3 ;
  RECT 1944.260 6.340 1944.460 6.540 ;
  LAYER VI3 ;
  RECT 1944.260 5.940 1944.460 6.140 ;
  LAYER VI3 ;
  RECT 1943.860 6.340 1944.060 6.540 ;
  LAYER VI3 ;
  RECT 1943.860 5.940 1944.060 6.140 ;
  LAYER VI3 ;
  RECT 1943.460 6.340 1943.660 6.540 ;
  LAYER VI3 ;
  RECT 1943.460 5.940 1943.660 6.140 ;
  LAYER VI3 ;
  RECT 1943.060 6.340 1943.260 6.540 ;
  LAYER VI3 ;
  RECT 1943.060 5.940 1943.260 6.140 ;
  LAYER VI3 ;
  RECT 1962.900 5.880 1970.900 6.740 ;
  LAYER VI3 ;
  RECT 1970.500 6.340 1970.700 6.540 ;
  LAYER VI3 ;
  RECT 1970.500 5.940 1970.700 6.140 ;
  LAYER VI3 ;
  RECT 1970.100 6.340 1970.300 6.540 ;
  LAYER VI3 ;
  RECT 1970.100 5.940 1970.300 6.140 ;
  LAYER VI3 ;
  RECT 1969.700 6.340 1969.900 6.540 ;
  LAYER VI3 ;
  RECT 1969.700 5.940 1969.900 6.140 ;
  LAYER VI3 ;
  RECT 1969.300 6.340 1969.500 6.540 ;
  LAYER VI3 ;
  RECT 1969.300 5.940 1969.500 6.140 ;
  LAYER VI3 ;
  RECT 1968.900 6.340 1969.100 6.540 ;
  LAYER VI3 ;
  RECT 1968.900 5.940 1969.100 6.140 ;
  LAYER VI3 ;
  RECT 1968.500 6.340 1968.700 6.540 ;
  LAYER VI3 ;
  RECT 1968.500 5.940 1968.700 6.140 ;
  LAYER VI3 ;
  RECT 1968.100 6.340 1968.300 6.540 ;
  LAYER VI3 ;
  RECT 1968.100 5.940 1968.300 6.140 ;
  LAYER VI3 ;
  RECT 1967.700 6.340 1967.900 6.540 ;
  LAYER VI3 ;
  RECT 1967.700 5.940 1967.900 6.140 ;
  LAYER VI3 ;
  RECT 1967.300 6.340 1967.500 6.540 ;
  LAYER VI3 ;
  RECT 1967.300 5.940 1967.500 6.140 ;
  LAYER VI3 ;
  RECT 1966.900 6.340 1967.100 6.540 ;
  LAYER VI3 ;
  RECT 1966.900 5.940 1967.100 6.140 ;
  LAYER VI3 ;
  RECT 1966.500 6.340 1966.700 6.540 ;
  LAYER VI3 ;
  RECT 1966.500 5.940 1966.700 6.140 ;
  LAYER VI3 ;
  RECT 1966.100 6.340 1966.300 6.540 ;
  LAYER VI3 ;
  RECT 1966.100 5.940 1966.300 6.140 ;
  LAYER VI3 ;
  RECT 1965.700 6.340 1965.900 6.540 ;
  LAYER VI3 ;
  RECT 1965.700 5.940 1965.900 6.140 ;
  LAYER VI3 ;
  RECT 1965.300 6.340 1965.500 6.540 ;
  LAYER VI3 ;
  RECT 1965.300 5.940 1965.500 6.140 ;
  LAYER VI3 ;
  RECT 1964.900 6.340 1965.100 6.540 ;
  LAYER VI3 ;
  RECT 1964.900 5.940 1965.100 6.140 ;
  LAYER VI3 ;
  RECT 1964.500 6.340 1964.700 6.540 ;
  LAYER VI3 ;
  RECT 1964.500 5.940 1964.700 6.140 ;
  LAYER VI3 ;
  RECT 1964.100 6.340 1964.300 6.540 ;
  LAYER VI3 ;
  RECT 1964.100 5.940 1964.300 6.140 ;
  LAYER VI3 ;
  RECT 1963.700 6.340 1963.900 6.540 ;
  LAYER VI3 ;
  RECT 1963.700 5.940 1963.900 6.140 ;
  LAYER VI3 ;
  RECT 1963.300 6.340 1963.500 6.540 ;
  LAYER VI3 ;
  RECT 1963.300 5.940 1963.500 6.140 ;
  LAYER VI3 ;
  RECT 1962.900 6.340 1963.100 6.540 ;
  LAYER VI3 ;
  RECT 1962.900 5.940 1963.100 6.140 ;
  LAYER VI3 ;
  RECT 1983.980 5.880 1991.980 6.740 ;
  LAYER VI3 ;
  RECT 1991.580 6.340 1991.780 6.540 ;
  LAYER VI3 ;
  RECT 1991.580 5.940 1991.780 6.140 ;
  LAYER VI3 ;
  RECT 1991.180 6.340 1991.380 6.540 ;
  LAYER VI3 ;
  RECT 1991.180 5.940 1991.380 6.140 ;
  LAYER VI3 ;
  RECT 1990.780 6.340 1990.980 6.540 ;
  LAYER VI3 ;
  RECT 1990.780 5.940 1990.980 6.140 ;
  LAYER VI3 ;
  RECT 1990.380 6.340 1990.580 6.540 ;
  LAYER VI3 ;
  RECT 1990.380 5.940 1990.580 6.140 ;
  LAYER VI3 ;
  RECT 1989.980 6.340 1990.180 6.540 ;
  LAYER VI3 ;
  RECT 1989.980 5.940 1990.180 6.140 ;
  LAYER VI3 ;
  RECT 1989.580 6.340 1989.780 6.540 ;
  LAYER VI3 ;
  RECT 1989.580 5.940 1989.780 6.140 ;
  LAYER VI3 ;
  RECT 1989.180 6.340 1989.380 6.540 ;
  LAYER VI3 ;
  RECT 1989.180 5.940 1989.380 6.140 ;
  LAYER VI3 ;
  RECT 1988.780 6.340 1988.980 6.540 ;
  LAYER VI3 ;
  RECT 1988.780 5.940 1988.980 6.140 ;
  LAYER VI3 ;
  RECT 1988.380 6.340 1988.580 6.540 ;
  LAYER VI3 ;
  RECT 1988.380 5.940 1988.580 6.140 ;
  LAYER VI3 ;
  RECT 1987.980 6.340 1988.180 6.540 ;
  LAYER VI3 ;
  RECT 1987.980 5.940 1988.180 6.140 ;
  LAYER VI3 ;
  RECT 1987.580 6.340 1987.780 6.540 ;
  LAYER VI3 ;
  RECT 1987.580 5.940 1987.780 6.140 ;
  LAYER VI3 ;
  RECT 1987.180 6.340 1987.380 6.540 ;
  LAYER VI3 ;
  RECT 1987.180 5.940 1987.380 6.140 ;
  LAYER VI3 ;
  RECT 1986.780 6.340 1986.980 6.540 ;
  LAYER VI3 ;
  RECT 1986.780 5.940 1986.980 6.140 ;
  LAYER VI3 ;
  RECT 1986.380 6.340 1986.580 6.540 ;
  LAYER VI3 ;
  RECT 1986.380 5.940 1986.580 6.140 ;
  LAYER VI3 ;
  RECT 1985.980 6.340 1986.180 6.540 ;
  LAYER VI3 ;
  RECT 1985.980 5.940 1986.180 6.140 ;
  LAYER VI3 ;
  RECT 1985.580 6.340 1985.780 6.540 ;
  LAYER VI3 ;
  RECT 1985.580 5.940 1985.780 6.140 ;
  LAYER VI3 ;
  RECT 1985.180 6.340 1985.380 6.540 ;
  LAYER VI3 ;
  RECT 1985.180 5.940 1985.380 6.140 ;
  LAYER VI3 ;
  RECT 1984.780 6.340 1984.980 6.540 ;
  LAYER VI3 ;
  RECT 1984.780 5.940 1984.980 6.140 ;
  LAYER VI3 ;
  RECT 1984.380 6.340 1984.580 6.540 ;
  LAYER VI3 ;
  RECT 1984.380 5.940 1984.580 6.140 ;
  LAYER VI3 ;
  RECT 1983.980 6.340 1984.180 6.540 ;
  LAYER VI3 ;
  RECT 1983.980 5.940 1984.180 6.140 ;
  LAYER VI3 ;
  RECT 2003.820 5.880 2011.820 6.740 ;
  LAYER VI3 ;
  RECT 2011.420 6.340 2011.620 6.540 ;
  LAYER VI3 ;
  RECT 2011.420 5.940 2011.620 6.140 ;
  LAYER VI3 ;
  RECT 2011.020 6.340 2011.220 6.540 ;
  LAYER VI3 ;
  RECT 2011.020 5.940 2011.220 6.140 ;
  LAYER VI3 ;
  RECT 2010.620 6.340 2010.820 6.540 ;
  LAYER VI3 ;
  RECT 2010.620 5.940 2010.820 6.140 ;
  LAYER VI3 ;
  RECT 2010.220 6.340 2010.420 6.540 ;
  LAYER VI3 ;
  RECT 2010.220 5.940 2010.420 6.140 ;
  LAYER VI3 ;
  RECT 2009.820 6.340 2010.020 6.540 ;
  LAYER VI3 ;
  RECT 2009.820 5.940 2010.020 6.140 ;
  LAYER VI3 ;
  RECT 2009.420 6.340 2009.620 6.540 ;
  LAYER VI3 ;
  RECT 2009.420 5.940 2009.620 6.140 ;
  LAYER VI3 ;
  RECT 2009.020 6.340 2009.220 6.540 ;
  LAYER VI3 ;
  RECT 2009.020 5.940 2009.220 6.140 ;
  LAYER VI3 ;
  RECT 2008.620 6.340 2008.820 6.540 ;
  LAYER VI3 ;
  RECT 2008.620 5.940 2008.820 6.140 ;
  LAYER VI3 ;
  RECT 2008.220 6.340 2008.420 6.540 ;
  LAYER VI3 ;
  RECT 2008.220 5.940 2008.420 6.140 ;
  LAYER VI3 ;
  RECT 2007.820 6.340 2008.020 6.540 ;
  LAYER VI3 ;
  RECT 2007.820 5.940 2008.020 6.140 ;
  LAYER VI3 ;
  RECT 2007.420 6.340 2007.620 6.540 ;
  LAYER VI3 ;
  RECT 2007.420 5.940 2007.620 6.140 ;
  LAYER VI3 ;
  RECT 2007.020 6.340 2007.220 6.540 ;
  LAYER VI3 ;
  RECT 2007.020 5.940 2007.220 6.140 ;
  LAYER VI3 ;
  RECT 2006.620 6.340 2006.820 6.540 ;
  LAYER VI3 ;
  RECT 2006.620 5.940 2006.820 6.140 ;
  LAYER VI3 ;
  RECT 2006.220 6.340 2006.420 6.540 ;
  LAYER VI3 ;
  RECT 2006.220 5.940 2006.420 6.140 ;
  LAYER VI3 ;
  RECT 2005.820 6.340 2006.020 6.540 ;
  LAYER VI3 ;
  RECT 2005.820 5.940 2006.020 6.140 ;
  LAYER VI3 ;
  RECT 2005.420 6.340 2005.620 6.540 ;
  LAYER VI3 ;
  RECT 2005.420 5.940 2005.620 6.140 ;
  LAYER VI3 ;
  RECT 2005.020 6.340 2005.220 6.540 ;
  LAYER VI3 ;
  RECT 2005.020 5.940 2005.220 6.140 ;
  LAYER VI3 ;
  RECT 2004.620 6.340 2004.820 6.540 ;
  LAYER VI3 ;
  RECT 2004.620 5.940 2004.820 6.140 ;
  LAYER VI3 ;
  RECT 2004.220 6.340 2004.420 6.540 ;
  LAYER VI3 ;
  RECT 2004.220 5.940 2004.420 6.140 ;
  LAYER VI3 ;
  RECT 2003.820 6.340 2004.020 6.540 ;
  LAYER VI3 ;
  RECT 2003.820 5.940 2004.020 6.140 ;
  LAYER VI3 ;
  RECT 2024.900 5.880 2032.900 6.740 ;
  LAYER VI3 ;
  RECT 2032.500 6.340 2032.700 6.540 ;
  LAYER VI3 ;
  RECT 2032.500 5.940 2032.700 6.140 ;
  LAYER VI3 ;
  RECT 2032.100 6.340 2032.300 6.540 ;
  LAYER VI3 ;
  RECT 2032.100 5.940 2032.300 6.140 ;
  LAYER VI3 ;
  RECT 2031.700 6.340 2031.900 6.540 ;
  LAYER VI3 ;
  RECT 2031.700 5.940 2031.900 6.140 ;
  LAYER VI3 ;
  RECT 2031.300 6.340 2031.500 6.540 ;
  LAYER VI3 ;
  RECT 2031.300 5.940 2031.500 6.140 ;
  LAYER VI3 ;
  RECT 2030.900 6.340 2031.100 6.540 ;
  LAYER VI3 ;
  RECT 2030.900 5.940 2031.100 6.140 ;
  LAYER VI3 ;
  RECT 2030.500 6.340 2030.700 6.540 ;
  LAYER VI3 ;
  RECT 2030.500 5.940 2030.700 6.140 ;
  LAYER VI3 ;
  RECT 2030.100 6.340 2030.300 6.540 ;
  LAYER VI3 ;
  RECT 2030.100 5.940 2030.300 6.140 ;
  LAYER VI3 ;
  RECT 2029.700 6.340 2029.900 6.540 ;
  LAYER VI3 ;
  RECT 2029.700 5.940 2029.900 6.140 ;
  LAYER VI3 ;
  RECT 2029.300 6.340 2029.500 6.540 ;
  LAYER VI3 ;
  RECT 2029.300 5.940 2029.500 6.140 ;
  LAYER VI3 ;
  RECT 2028.900 6.340 2029.100 6.540 ;
  LAYER VI3 ;
  RECT 2028.900 5.940 2029.100 6.140 ;
  LAYER VI3 ;
  RECT 2028.500 6.340 2028.700 6.540 ;
  LAYER VI3 ;
  RECT 2028.500 5.940 2028.700 6.140 ;
  LAYER VI3 ;
  RECT 2028.100 6.340 2028.300 6.540 ;
  LAYER VI3 ;
  RECT 2028.100 5.940 2028.300 6.140 ;
  LAYER VI3 ;
  RECT 2027.700 6.340 2027.900 6.540 ;
  LAYER VI3 ;
  RECT 2027.700 5.940 2027.900 6.140 ;
  LAYER VI3 ;
  RECT 2027.300 6.340 2027.500 6.540 ;
  LAYER VI3 ;
  RECT 2027.300 5.940 2027.500 6.140 ;
  LAYER VI3 ;
  RECT 2026.900 6.340 2027.100 6.540 ;
  LAYER VI3 ;
  RECT 2026.900 5.940 2027.100 6.140 ;
  LAYER VI3 ;
  RECT 2026.500 6.340 2026.700 6.540 ;
  LAYER VI3 ;
  RECT 2026.500 5.940 2026.700 6.140 ;
  LAYER VI3 ;
  RECT 2026.100 6.340 2026.300 6.540 ;
  LAYER VI3 ;
  RECT 2026.100 5.940 2026.300 6.140 ;
  LAYER VI3 ;
  RECT 2025.700 6.340 2025.900 6.540 ;
  LAYER VI3 ;
  RECT 2025.700 5.940 2025.900 6.140 ;
  LAYER VI3 ;
  RECT 2025.300 6.340 2025.500 6.540 ;
  LAYER VI3 ;
  RECT 2025.300 5.940 2025.500 6.140 ;
  LAYER VI3 ;
  RECT 2024.900 6.340 2025.100 6.540 ;
  LAYER VI3 ;
  RECT 2024.900 5.940 2025.100 6.140 ;
  LAYER VI3 ;
  RECT 2044.740 5.880 2052.740 6.740 ;
  LAYER VI3 ;
  RECT 2052.340 6.340 2052.540 6.540 ;
  LAYER VI3 ;
  RECT 2052.340 5.940 2052.540 6.140 ;
  LAYER VI3 ;
  RECT 2051.940 6.340 2052.140 6.540 ;
  LAYER VI3 ;
  RECT 2051.940 5.940 2052.140 6.140 ;
  LAYER VI3 ;
  RECT 2051.540 6.340 2051.740 6.540 ;
  LAYER VI3 ;
  RECT 2051.540 5.940 2051.740 6.140 ;
  LAYER VI3 ;
  RECT 2051.140 6.340 2051.340 6.540 ;
  LAYER VI3 ;
  RECT 2051.140 5.940 2051.340 6.140 ;
  LAYER VI3 ;
  RECT 2050.740 6.340 2050.940 6.540 ;
  LAYER VI3 ;
  RECT 2050.740 5.940 2050.940 6.140 ;
  LAYER VI3 ;
  RECT 2050.340 6.340 2050.540 6.540 ;
  LAYER VI3 ;
  RECT 2050.340 5.940 2050.540 6.140 ;
  LAYER VI3 ;
  RECT 2049.940 6.340 2050.140 6.540 ;
  LAYER VI3 ;
  RECT 2049.940 5.940 2050.140 6.140 ;
  LAYER VI3 ;
  RECT 2049.540 6.340 2049.740 6.540 ;
  LAYER VI3 ;
  RECT 2049.540 5.940 2049.740 6.140 ;
  LAYER VI3 ;
  RECT 2049.140 6.340 2049.340 6.540 ;
  LAYER VI3 ;
  RECT 2049.140 5.940 2049.340 6.140 ;
  LAYER VI3 ;
  RECT 2048.740 6.340 2048.940 6.540 ;
  LAYER VI3 ;
  RECT 2048.740 5.940 2048.940 6.140 ;
  LAYER VI3 ;
  RECT 2048.340 6.340 2048.540 6.540 ;
  LAYER VI3 ;
  RECT 2048.340 5.940 2048.540 6.140 ;
  LAYER VI3 ;
  RECT 2047.940 6.340 2048.140 6.540 ;
  LAYER VI3 ;
  RECT 2047.940 5.940 2048.140 6.140 ;
  LAYER VI3 ;
  RECT 2047.540 6.340 2047.740 6.540 ;
  LAYER VI3 ;
  RECT 2047.540 5.940 2047.740 6.140 ;
  LAYER VI3 ;
  RECT 2047.140 6.340 2047.340 6.540 ;
  LAYER VI3 ;
  RECT 2047.140 5.940 2047.340 6.140 ;
  LAYER VI3 ;
  RECT 2046.740 6.340 2046.940 6.540 ;
  LAYER VI3 ;
  RECT 2046.740 5.940 2046.940 6.140 ;
  LAYER VI3 ;
  RECT 2046.340 6.340 2046.540 6.540 ;
  LAYER VI3 ;
  RECT 2046.340 5.940 2046.540 6.140 ;
  LAYER VI3 ;
  RECT 2045.940 6.340 2046.140 6.540 ;
  LAYER VI3 ;
  RECT 2045.940 5.940 2046.140 6.140 ;
  LAYER VI3 ;
  RECT 2045.540 6.340 2045.740 6.540 ;
  LAYER VI3 ;
  RECT 2045.540 5.940 2045.740 6.140 ;
  LAYER VI3 ;
  RECT 2045.140 6.340 2045.340 6.540 ;
  LAYER VI3 ;
  RECT 2045.140 5.940 2045.340 6.140 ;
  LAYER VI3 ;
  RECT 2044.740 6.340 2044.940 6.540 ;
  LAYER VI3 ;
  RECT 2044.740 5.940 2044.940 6.140 ;
  LAYER VI3 ;
  RECT 2065.820 5.880 2073.820 6.740 ;
  LAYER VI3 ;
  RECT 2073.420 6.340 2073.620 6.540 ;
  LAYER VI3 ;
  RECT 2073.420 5.940 2073.620 6.140 ;
  LAYER VI3 ;
  RECT 2073.020 6.340 2073.220 6.540 ;
  LAYER VI3 ;
  RECT 2073.020 5.940 2073.220 6.140 ;
  LAYER VI3 ;
  RECT 2072.620 6.340 2072.820 6.540 ;
  LAYER VI3 ;
  RECT 2072.620 5.940 2072.820 6.140 ;
  LAYER VI3 ;
  RECT 2072.220 6.340 2072.420 6.540 ;
  LAYER VI3 ;
  RECT 2072.220 5.940 2072.420 6.140 ;
  LAYER VI3 ;
  RECT 2071.820 6.340 2072.020 6.540 ;
  LAYER VI3 ;
  RECT 2071.820 5.940 2072.020 6.140 ;
  LAYER VI3 ;
  RECT 2071.420 6.340 2071.620 6.540 ;
  LAYER VI3 ;
  RECT 2071.420 5.940 2071.620 6.140 ;
  LAYER VI3 ;
  RECT 2071.020 6.340 2071.220 6.540 ;
  LAYER VI3 ;
  RECT 2071.020 5.940 2071.220 6.140 ;
  LAYER VI3 ;
  RECT 2070.620 6.340 2070.820 6.540 ;
  LAYER VI3 ;
  RECT 2070.620 5.940 2070.820 6.140 ;
  LAYER VI3 ;
  RECT 2070.220 6.340 2070.420 6.540 ;
  LAYER VI3 ;
  RECT 2070.220 5.940 2070.420 6.140 ;
  LAYER VI3 ;
  RECT 2069.820 6.340 2070.020 6.540 ;
  LAYER VI3 ;
  RECT 2069.820 5.940 2070.020 6.140 ;
  LAYER VI3 ;
  RECT 2069.420 6.340 2069.620 6.540 ;
  LAYER VI3 ;
  RECT 2069.420 5.940 2069.620 6.140 ;
  LAYER VI3 ;
  RECT 2069.020 6.340 2069.220 6.540 ;
  LAYER VI3 ;
  RECT 2069.020 5.940 2069.220 6.140 ;
  LAYER VI3 ;
  RECT 2068.620 6.340 2068.820 6.540 ;
  LAYER VI3 ;
  RECT 2068.620 5.940 2068.820 6.140 ;
  LAYER VI3 ;
  RECT 2068.220 6.340 2068.420 6.540 ;
  LAYER VI3 ;
  RECT 2068.220 5.940 2068.420 6.140 ;
  LAYER VI3 ;
  RECT 2067.820 6.340 2068.020 6.540 ;
  LAYER VI3 ;
  RECT 2067.820 5.940 2068.020 6.140 ;
  LAYER VI3 ;
  RECT 2067.420 6.340 2067.620 6.540 ;
  LAYER VI3 ;
  RECT 2067.420 5.940 2067.620 6.140 ;
  LAYER VI3 ;
  RECT 2067.020 6.340 2067.220 6.540 ;
  LAYER VI3 ;
  RECT 2067.020 5.940 2067.220 6.140 ;
  LAYER VI3 ;
  RECT 2066.620 6.340 2066.820 6.540 ;
  LAYER VI3 ;
  RECT 2066.620 5.940 2066.820 6.140 ;
  LAYER VI3 ;
  RECT 2066.220 6.340 2066.420 6.540 ;
  LAYER VI3 ;
  RECT 2066.220 5.940 2066.420 6.140 ;
  LAYER VI3 ;
  RECT 2065.820 6.340 2066.020 6.540 ;
  LAYER VI3 ;
  RECT 2065.820 5.940 2066.020 6.140 ;
  LAYER VI3 ;
  RECT 2085.660 5.880 2093.660 6.740 ;
  LAYER VI3 ;
  RECT 2093.260 6.340 2093.460 6.540 ;
  LAYER VI3 ;
  RECT 2093.260 5.940 2093.460 6.140 ;
  LAYER VI3 ;
  RECT 2092.860 6.340 2093.060 6.540 ;
  LAYER VI3 ;
  RECT 2092.860 5.940 2093.060 6.140 ;
  LAYER VI3 ;
  RECT 2092.460 6.340 2092.660 6.540 ;
  LAYER VI3 ;
  RECT 2092.460 5.940 2092.660 6.140 ;
  LAYER VI3 ;
  RECT 2092.060 6.340 2092.260 6.540 ;
  LAYER VI3 ;
  RECT 2092.060 5.940 2092.260 6.140 ;
  LAYER VI3 ;
  RECT 2091.660 6.340 2091.860 6.540 ;
  LAYER VI3 ;
  RECT 2091.660 5.940 2091.860 6.140 ;
  LAYER VI3 ;
  RECT 2091.260 6.340 2091.460 6.540 ;
  LAYER VI3 ;
  RECT 2091.260 5.940 2091.460 6.140 ;
  LAYER VI3 ;
  RECT 2090.860 6.340 2091.060 6.540 ;
  LAYER VI3 ;
  RECT 2090.860 5.940 2091.060 6.140 ;
  LAYER VI3 ;
  RECT 2090.460 6.340 2090.660 6.540 ;
  LAYER VI3 ;
  RECT 2090.460 5.940 2090.660 6.140 ;
  LAYER VI3 ;
  RECT 2090.060 6.340 2090.260 6.540 ;
  LAYER VI3 ;
  RECT 2090.060 5.940 2090.260 6.140 ;
  LAYER VI3 ;
  RECT 2089.660 6.340 2089.860 6.540 ;
  LAYER VI3 ;
  RECT 2089.660 5.940 2089.860 6.140 ;
  LAYER VI3 ;
  RECT 2089.260 6.340 2089.460 6.540 ;
  LAYER VI3 ;
  RECT 2089.260 5.940 2089.460 6.140 ;
  LAYER VI3 ;
  RECT 2088.860 6.340 2089.060 6.540 ;
  LAYER VI3 ;
  RECT 2088.860 5.940 2089.060 6.140 ;
  LAYER VI3 ;
  RECT 2088.460 6.340 2088.660 6.540 ;
  LAYER VI3 ;
  RECT 2088.460 5.940 2088.660 6.140 ;
  LAYER VI3 ;
  RECT 2088.060 6.340 2088.260 6.540 ;
  LAYER VI3 ;
  RECT 2088.060 5.940 2088.260 6.140 ;
  LAYER VI3 ;
  RECT 2087.660 6.340 2087.860 6.540 ;
  LAYER VI3 ;
  RECT 2087.660 5.940 2087.860 6.140 ;
  LAYER VI3 ;
  RECT 2087.260 6.340 2087.460 6.540 ;
  LAYER VI3 ;
  RECT 2087.260 5.940 2087.460 6.140 ;
  LAYER VI3 ;
  RECT 2086.860 6.340 2087.060 6.540 ;
  LAYER VI3 ;
  RECT 2086.860 5.940 2087.060 6.140 ;
  LAYER VI3 ;
  RECT 2086.460 6.340 2086.660 6.540 ;
  LAYER VI3 ;
  RECT 2086.460 5.940 2086.660 6.140 ;
  LAYER VI3 ;
  RECT 2086.060 6.340 2086.260 6.540 ;
  LAYER VI3 ;
  RECT 2086.060 5.940 2086.260 6.140 ;
  LAYER VI3 ;
  RECT 2085.660 6.340 2085.860 6.540 ;
  LAYER VI3 ;
  RECT 2085.660 5.940 2085.860 6.140 ;
  LAYER VI3 ;
  RECT 2106.740 5.880 2114.740 6.740 ;
  LAYER VI3 ;
  RECT 2114.340 6.340 2114.540 6.540 ;
  LAYER VI3 ;
  RECT 2114.340 5.940 2114.540 6.140 ;
  LAYER VI3 ;
  RECT 2113.940 6.340 2114.140 6.540 ;
  LAYER VI3 ;
  RECT 2113.940 5.940 2114.140 6.140 ;
  LAYER VI3 ;
  RECT 2113.540 6.340 2113.740 6.540 ;
  LAYER VI3 ;
  RECT 2113.540 5.940 2113.740 6.140 ;
  LAYER VI3 ;
  RECT 2113.140 6.340 2113.340 6.540 ;
  LAYER VI3 ;
  RECT 2113.140 5.940 2113.340 6.140 ;
  LAYER VI3 ;
  RECT 2112.740 6.340 2112.940 6.540 ;
  LAYER VI3 ;
  RECT 2112.740 5.940 2112.940 6.140 ;
  LAYER VI3 ;
  RECT 2112.340 6.340 2112.540 6.540 ;
  LAYER VI3 ;
  RECT 2112.340 5.940 2112.540 6.140 ;
  LAYER VI3 ;
  RECT 2111.940 6.340 2112.140 6.540 ;
  LAYER VI3 ;
  RECT 2111.940 5.940 2112.140 6.140 ;
  LAYER VI3 ;
  RECT 2111.540 6.340 2111.740 6.540 ;
  LAYER VI3 ;
  RECT 2111.540 5.940 2111.740 6.140 ;
  LAYER VI3 ;
  RECT 2111.140 6.340 2111.340 6.540 ;
  LAYER VI3 ;
  RECT 2111.140 5.940 2111.340 6.140 ;
  LAYER VI3 ;
  RECT 2110.740 6.340 2110.940 6.540 ;
  LAYER VI3 ;
  RECT 2110.740 5.940 2110.940 6.140 ;
  LAYER VI3 ;
  RECT 2110.340 6.340 2110.540 6.540 ;
  LAYER VI3 ;
  RECT 2110.340 5.940 2110.540 6.140 ;
  LAYER VI3 ;
  RECT 2109.940 6.340 2110.140 6.540 ;
  LAYER VI3 ;
  RECT 2109.940 5.940 2110.140 6.140 ;
  LAYER VI3 ;
  RECT 2109.540 6.340 2109.740 6.540 ;
  LAYER VI3 ;
  RECT 2109.540 5.940 2109.740 6.140 ;
  LAYER VI3 ;
  RECT 2109.140 6.340 2109.340 6.540 ;
  LAYER VI3 ;
  RECT 2109.140 5.940 2109.340 6.140 ;
  LAYER VI3 ;
  RECT 2108.740 6.340 2108.940 6.540 ;
  LAYER VI3 ;
  RECT 2108.740 5.940 2108.940 6.140 ;
  LAYER VI3 ;
  RECT 2108.340 6.340 2108.540 6.540 ;
  LAYER VI3 ;
  RECT 2108.340 5.940 2108.540 6.140 ;
  LAYER VI3 ;
  RECT 2107.940 6.340 2108.140 6.540 ;
  LAYER VI3 ;
  RECT 2107.940 5.940 2108.140 6.140 ;
  LAYER VI3 ;
  RECT 2107.540 6.340 2107.740 6.540 ;
  LAYER VI3 ;
  RECT 2107.540 5.940 2107.740 6.140 ;
  LAYER VI3 ;
  RECT 2107.140 6.340 2107.340 6.540 ;
  LAYER VI3 ;
  RECT 2107.140 5.940 2107.340 6.140 ;
  LAYER VI3 ;
  RECT 2106.740 6.340 2106.940 6.540 ;
  LAYER VI3 ;
  RECT 2106.740 5.940 2106.940 6.140 ;
  LAYER VI3 ;
  RECT 2126.580 5.880 2134.580 6.740 ;
  LAYER VI3 ;
  RECT 2134.180 6.340 2134.380 6.540 ;
  LAYER VI3 ;
  RECT 2134.180 5.940 2134.380 6.140 ;
  LAYER VI3 ;
  RECT 2133.780 6.340 2133.980 6.540 ;
  LAYER VI3 ;
  RECT 2133.780 5.940 2133.980 6.140 ;
  LAYER VI3 ;
  RECT 2133.380 6.340 2133.580 6.540 ;
  LAYER VI3 ;
  RECT 2133.380 5.940 2133.580 6.140 ;
  LAYER VI3 ;
  RECT 2132.980 6.340 2133.180 6.540 ;
  LAYER VI3 ;
  RECT 2132.980 5.940 2133.180 6.140 ;
  LAYER VI3 ;
  RECT 2132.580 6.340 2132.780 6.540 ;
  LAYER VI3 ;
  RECT 2132.580 5.940 2132.780 6.140 ;
  LAYER VI3 ;
  RECT 2132.180 6.340 2132.380 6.540 ;
  LAYER VI3 ;
  RECT 2132.180 5.940 2132.380 6.140 ;
  LAYER VI3 ;
  RECT 2131.780 6.340 2131.980 6.540 ;
  LAYER VI3 ;
  RECT 2131.780 5.940 2131.980 6.140 ;
  LAYER VI3 ;
  RECT 2131.380 6.340 2131.580 6.540 ;
  LAYER VI3 ;
  RECT 2131.380 5.940 2131.580 6.140 ;
  LAYER VI3 ;
  RECT 2130.980 6.340 2131.180 6.540 ;
  LAYER VI3 ;
  RECT 2130.980 5.940 2131.180 6.140 ;
  LAYER VI3 ;
  RECT 2130.580 6.340 2130.780 6.540 ;
  LAYER VI3 ;
  RECT 2130.580 5.940 2130.780 6.140 ;
  LAYER VI3 ;
  RECT 2130.180 6.340 2130.380 6.540 ;
  LAYER VI3 ;
  RECT 2130.180 5.940 2130.380 6.140 ;
  LAYER VI3 ;
  RECT 2129.780 6.340 2129.980 6.540 ;
  LAYER VI3 ;
  RECT 2129.780 5.940 2129.980 6.140 ;
  LAYER VI3 ;
  RECT 2129.380 6.340 2129.580 6.540 ;
  LAYER VI3 ;
  RECT 2129.380 5.940 2129.580 6.140 ;
  LAYER VI3 ;
  RECT 2128.980 6.340 2129.180 6.540 ;
  LAYER VI3 ;
  RECT 2128.980 5.940 2129.180 6.140 ;
  LAYER VI3 ;
  RECT 2128.580 6.340 2128.780 6.540 ;
  LAYER VI3 ;
  RECT 2128.580 5.940 2128.780 6.140 ;
  LAYER VI3 ;
  RECT 2128.180 6.340 2128.380 6.540 ;
  LAYER VI3 ;
  RECT 2128.180 5.940 2128.380 6.140 ;
  LAYER VI3 ;
  RECT 2127.780 6.340 2127.980 6.540 ;
  LAYER VI3 ;
  RECT 2127.780 5.940 2127.980 6.140 ;
  LAYER VI3 ;
  RECT 2127.380 6.340 2127.580 6.540 ;
  LAYER VI3 ;
  RECT 2127.380 5.940 2127.580 6.140 ;
  LAYER VI3 ;
  RECT 2126.980 6.340 2127.180 6.540 ;
  LAYER VI3 ;
  RECT 2126.980 5.940 2127.180 6.140 ;
  LAYER VI3 ;
  RECT 2126.580 6.340 2126.780 6.540 ;
  LAYER VI3 ;
  RECT 2126.580 5.940 2126.780 6.140 ;
  LAYER VI3 ;
  RECT 2147.660 5.880 2155.660 6.740 ;
  LAYER VI3 ;
  RECT 2155.260 6.340 2155.460 6.540 ;
  LAYER VI3 ;
  RECT 2155.260 5.940 2155.460 6.140 ;
  LAYER VI3 ;
  RECT 2154.860 6.340 2155.060 6.540 ;
  LAYER VI3 ;
  RECT 2154.860 5.940 2155.060 6.140 ;
  LAYER VI3 ;
  RECT 2154.460 6.340 2154.660 6.540 ;
  LAYER VI3 ;
  RECT 2154.460 5.940 2154.660 6.140 ;
  LAYER VI3 ;
  RECT 2154.060 6.340 2154.260 6.540 ;
  LAYER VI3 ;
  RECT 2154.060 5.940 2154.260 6.140 ;
  LAYER VI3 ;
  RECT 2153.660 6.340 2153.860 6.540 ;
  LAYER VI3 ;
  RECT 2153.660 5.940 2153.860 6.140 ;
  LAYER VI3 ;
  RECT 2153.260 6.340 2153.460 6.540 ;
  LAYER VI3 ;
  RECT 2153.260 5.940 2153.460 6.140 ;
  LAYER VI3 ;
  RECT 2152.860 6.340 2153.060 6.540 ;
  LAYER VI3 ;
  RECT 2152.860 5.940 2153.060 6.140 ;
  LAYER VI3 ;
  RECT 2152.460 6.340 2152.660 6.540 ;
  LAYER VI3 ;
  RECT 2152.460 5.940 2152.660 6.140 ;
  LAYER VI3 ;
  RECT 2152.060 6.340 2152.260 6.540 ;
  LAYER VI3 ;
  RECT 2152.060 5.940 2152.260 6.140 ;
  LAYER VI3 ;
  RECT 2151.660 6.340 2151.860 6.540 ;
  LAYER VI3 ;
  RECT 2151.660 5.940 2151.860 6.140 ;
  LAYER VI3 ;
  RECT 2151.260 6.340 2151.460 6.540 ;
  LAYER VI3 ;
  RECT 2151.260 5.940 2151.460 6.140 ;
  LAYER VI3 ;
  RECT 2150.860 6.340 2151.060 6.540 ;
  LAYER VI3 ;
  RECT 2150.860 5.940 2151.060 6.140 ;
  LAYER VI3 ;
  RECT 2150.460 6.340 2150.660 6.540 ;
  LAYER VI3 ;
  RECT 2150.460 5.940 2150.660 6.140 ;
  LAYER VI3 ;
  RECT 2150.060 6.340 2150.260 6.540 ;
  LAYER VI3 ;
  RECT 2150.060 5.940 2150.260 6.140 ;
  LAYER VI3 ;
  RECT 2149.660 6.340 2149.860 6.540 ;
  LAYER VI3 ;
  RECT 2149.660 5.940 2149.860 6.140 ;
  LAYER VI3 ;
  RECT 2149.260 6.340 2149.460 6.540 ;
  LAYER VI3 ;
  RECT 2149.260 5.940 2149.460 6.140 ;
  LAYER VI3 ;
  RECT 2148.860 6.340 2149.060 6.540 ;
  LAYER VI3 ;
  RECT 2148.860 5.940 2149.060 6.140 ;
  LAYER VI3 ;
  RECT 2148.460 6.340 2148.660 6.540 ;
  LAYER VI3 ;
  RECT 2148.460 5.940 2148.660 6.140 ;
  LAYER VI3 ;
  RECT 2148.060 6.340 2148.260 6.540 ;
  LAYER VI3 ;
  RECT 2148.060 5.940 2148.260 6.140 ;
  LAYER VI3 ;
  RECT 2147.660 6.340 2147.860 6.540 ;
  LAYER VI3 ;
  RECT 2147.660 5.940 2147.860 6.140 ;
  LAYER VI3 ;
  RECT 2167.500 5.880 2175.500 6.740 ;
  LAYER VI3 ;
  RECT 2175.100 6.340 2175.300 6.540 ;
  LAYER VI3 ;
  RECT 2175.100 5.940 2175.300 6.140 ;
  LAYER VI3 ;
  RECT 2174.700 6.340 2174.900 6.540 ;
  LAYER VI3 ;
  RECT 2174.700 5.940 2174.900 6.140 ;
  LAYER VI3 ;
  RECT 2174.300 6.340 2174.500 6.540 ;
  LAYER VI3 ;
  RECT 2174.300 5.940 2174.500 6.140 ;
  LAYER VI3 ;
  RECT 2173.900 6.340 2174.100 6.540 ;
  LAYER VI3 ;
  RECT 2173.900 5.940 2174.100 6.140 ;
  LAYER VI3 ;
  RECT 2173.500 6.340 2173.700 6.540 ;
  LAYER VI3 ;
  RECT 2173.500 5.940 2173.700 6.140 ;
  LAYER VI3 ;
  RECT 2173.100 6.340 2173.300 6.540 ;
  LAYER VI3 ;
  RECT 2173.100 5.940 2173.300 6.140 ;
  LAYER VI3 ;
  RECT 2172.700 6.340 2172.900 6.540 ;
  LAYER VI3 ;
  RECT 2172.700 5.940 2172.900 6.140 ;
  LAYER VI3 ;
  RECT 2172.300 6.340 2172.500 6.540 ;
  LAYER VI3 ;
  RECT 2172.300 5.940 2172.500 6.140 ;
  LAYER VI3 ;
  RECT 2171.900 6.340 2172.100 6.540 ;
  LAYER VI3 ;
  RECT 2171.900 5.940 2172.100 6.140 ;
  LAYER VI3 ;
  RECT 2171.500 6.340 2171.700 6.540 ;
  LAYER VI3 ;
  RECT 2171.500 5.940 2171.700 6.140 ;
  LAYER VI3 ;
  RECT 2171.100 6.340 2171.300 6.540 ;
  LAYER VI3 ;
  RECT 2171.100 5.940 2171.300 6.140 ;
  LAYER VI3 ;
  RECT 2170.700 6.340 2170.900 6.540 ;
  LAYER VI3 ;
  RECT 2170.700 5.940 2170.900 6.140 ;
  LAYER VI3 ;
  RECT 2170.300 6.340 2170.500 6.540 ;
  LAYER VI3 ;
  RECT 2170.300 5.940 2170.500 6.140 ;
  LAYER VI3 ;
  RECT 2169.900 6.340 2170.100 6.540 ;
  LAYER VI3 ;
  RECT 2169.900 5.940 2170.100 6.140 ;
  LAYER VI3 ;
  RECT 2169.500 6.340 2169.700 6.540 ;
  LAYER VI3 ;
  RECT 2169.500 5.940 2169.700 6.140 ;
  LAYER VI3 ;
  RECT 2169.100 6.340 2169.300 6.540 ;
  LAYER VI3 ;
  RECT 2169.100 5.940 2169.300 6.140 ;
  LAYER VI3 ;
  RECT 2168.700 6.340 2168.900 6.540 ;
  LAYER VI3 ;
  RECT 2168.700 5.940 2168.900 6.140 ;
  LAYER VI3 ;
  RECT 2168.300 6.340 2168.500 6.540 ;
  LAYER VI3 ;
  RECT 2168.300 5.940 2168.500 6.140 ;
  LAYER VI3 ;
  RECT 2167.900 6.340 2168.100 6.540 ;
  LAYER VI3 ;
  RECT 2167.900 5.940 2168.100 6.140 ;
  LAYER VI3 ;
  RECT 2167.500 6.340 2167.700 6.540 ;
  LAYER VI3 ;
  RECT 2167.500 5.940 2167.700 6.140 ;
  LAYER VI3 ;
  RECT 2188.580 5.880 2196.580 6.740 ;
  LAYER VI3 ;
  RECT 2196.180 6.340 2196.380 6.540 ;
  LAYER VI3 ;
  RECT 2196.180 5.940 2196.380 6.140 ;
  LAYER VI3 ;
  RECT 2195.780 6.340 2195.980 6.540 ;
  LAYER VI3 ;
  RECT 2195.780 5.940 2195.980 6.140 ;
  LAYER VI3 ;
  RECT 2195.380 6.340 2195.580 6.540 ;
  LAYER VI3 ;
  RECT 2195.380 5.940 2195.580 6.140 ;
  LAYER VI3 ;
  RECT 2194.980 6.340 2195.180 6.540 ;
  LAYER VI3 ;
  RECT 2194.980 5.940 2195.180 6.140 ;
  LAYER VI3 ;
  RECT 2194.580 6.340 2194.780 6.540 ;
  LAYER VI3 ;
  RECT 2194.580 5.940 2194.780 6.140 ;
  LAYER VI3 ;
  RECT 2194.180 6.340 2194.380 6.540 ;
  LAYER VI3 ;
  RECT 2194.180 5.940 2194.380 6.140 ;
  LAYER VI3 ;
  RECT 2193.780 6.340 2193.980 6.540 ;
  LAYER VI3 ;
  RECT 2193.780 5.940 2193.980 6.140 ;
  LAYER VI3 ;
  RECT 2193.380 6.340 2193.580 6.540 ;
  LAYER VI3 ;
  RECT 2193.380 5.940 2193.580 6.140 ;
  LAYER VI3 ;
  RECT 2192.980 6.340 2193.180 6.540 ;
  LAYER VI3 ;
  RECT 2192.980 5.940 2193.180 6.140 ;
  LAYER VI3 ;
  RECT 2192.580 6.340 2192.780 6.540 ;
  LAYER VI3 ;
  RECT 2192.580 5.940 2192.780 6.140 ;
  LAYER VI3 ;
  RECT 2192.180 6.340 2192.380 6.540 ;
  LAYER VI3 ;
  RECT 2192.180 5.940 2192.380 6.140 ;
  LAYER VI3 ;
  RECT 2191.780 6.340 2191.980 6.540 ;
  LAYER VI3 ;
  RECT 2191.780 5.940 2191.980 6.140 ;
  LAYER VI3 ;
  RECT 2191.380 6.340 2191.580 6.540 ;
  LAYER VI3 ;
  RECT 2191.380 5.940 2191.580 6.140 ;
  LAYER VI3 ;
  RECT 2190.980 6.340 2191.180 6.540 ;
  LAYER VI3 ;
  RECT 2190.980 5.940 2191.180 6.140 ;
  LAYER VI3 ;
  RECT 2190.580 6.340 2190.780 6.540 ;
  LAYER VI3 ;
  RECT 2190.580 5.940 2190.780 6.140 ;
  LAYER VI3 ;
  RECT 2190.180 6.340 2190.380 6.540 ;
  LAYER VI3 ;
  RECT 2190.180 5.940 2190.380 6.140 ;
  LAYER VI3 ;
  RECT 2189.780 6.340 2189.980 6.540 ;
  LAYER VI3 ;
  RECT 2189.780 5.940 2189.980 6.140 ;
  LAYER VI3 ;
  RECT 2189.380 6.340 2189.580 6.540 ;
  LAYER VI3 ;
  RECT 2189.380 5.940 2189.580 6.140 ;
  LAYER VI3 ;
  RECT 2188.980 6.340 2189.180 6.540 ;
  LAYER VI3 ;
  RECT 2188.980 5.940 2189.180 6.140 ;
  LAYER VI3 ;
  RECT 2188.580 6.340 2188.780 6.540 ;
  LAYER VI3 ;
  RECT 2188.580 5.940 2188.780 6.140 ;
  LAYER VI3 ;
  RECT 2208.420 5.880 2216.420 6.740 ;
  LAYER VI3 ;
  RECT 2216.020 6.340 2216.220 6.540 ;
  LAYER VI3 ;
  RECT 2216.020 5.940 2216.220 6.140 ;
  LAYER VI3 ;
  RECT 2215.620 6.340 2215.820 6.540 ;
  LAYER VI3 ;
  RECT 2215.620 5.940 2215.820 6.140 ;
  LAYER VI3 ;
  RECT 2215.220 6.340 2215.420 6.540 ;
  LAYER VI3 ;
  RECT 2215.220 5.940 2215.420 6.140 ;
  LAYER VI3 ;
  RECT 2214.820 6.340 2215.020 6.540 ;
  LAYER VI3 ;
  RECT 2214.820 5.940 2215.020 6.140 ;
  LAYER VI3 ;
  RECT 2214.420 6.340 2214.620 6.540 ;
  LAYER VI3 ;
  RECT 2214.420 5.940 2214.620 6.140 ;
  LAYER VI3 ;
  RECT 2214.020 6.340 2214.220 6.540 ;
  LAYER VI3 ;
  RECT 2214.020 5.940 2214.220 6.140 ;
  LAYER VI3 ;
  RECT 2213.620 6.340 2213.820 6.540 ;
  LAYER VI3 ;
  RECT 2213.620 5.940 2213.820 6.140 ;
  LAYER VI3 ;
  RECT 2213.220 6.340 2213.420 6.540 ;
  LAYER VI3 ;
  RECT 2213.220 5.940 2213.420 6.140 ;
  LAYER VI3 ;
  RECT 2212.820 6.340 2213.020 6.540 ;
  LAYER VI3 ;
  RECT 2212.820 5.940 2213.020 6.140 ;
  LAYER VI3 ;
  RECT 2212.420 6.340 2212.620 6.540 ;
  LAYER VI3 ;
  RECT 2212.420 5.940 2212.620 6.140 ;
  LAYER VI3 ;
  RECT 2212.020 6.340 2212.220 6.540 ;
  LAYER VI3 ;
  RECT 2212.020 5.940 2212.220 6.140 ;
  LAYER VI3 ;
  RECT 2211.620 6.340 2211.820 6.540 ;
  LAYER VI3 ;
  RECT 2211.620 5.940 2211.820 6.140 ;
  LAYER VI3 ;
  RECT 2211.220 6.340 2211.420 6.540 ;
  LAYER VI3 ;
  RECT 2211.220 5.940 2211.420 6.140 ;
  LAYER VI3 ;
  RECT 2210.820 6.340 2211.020 6.540 ;
  LAYER VI3 ;
  RECT 2210.820 5.940 2211.020 6.140 ;
  LAYER VI3 ;
  RECT 2210.420 6.340 2210.620 6.540 ;
  LAYER VI3 ;
  RECT 2210.420 5.940 2210.620 6.140 ;
  LAYER VI3 ;
  RECT 2210.020 6.340 2210.220 6.540 ;
  LAYER VI3 ;
  RECT 2210.020 5.940 2210.220 6.140 ;
  LAYER VI3 ;
  RECT 2209.620 6.340 2209.820 6.540 ;
  LAYER VI3 ;
  RECT 2209.620 5.940 2209.820 6.140 ;
  LAYER VI3 ;
  RECT 2209.220 6.340 2209.420 6.540 ;
  LAYER VI3 ;
  RECT 2209.220 5.940 2209.420 6.140 ;
  LAYER VI3 ;
  RECT 2208.820 6.340 2209.020 6.540 ;
  LAYER VI3 ;
  RECT 2208.820 5.940 2209.020 6.140 ;
  LAYER VI3 ;
  RECT 2208.420 6.340 2208.620 6.540 ;
  LAYER VI3 ;
  RECT 2208.420 5.940 2208.620 6.140 ;
  LAYER VI3 ;
  RECT 2229.500 5.880 2237.500 6.740 ;
  LAYER VI3 ;
  RECT 2237.100 6.340 2237.300 6.540 ;
  LAYER VI3 ;
  RECT 2237.100 5.940 2237.300 6.140 ;
  LAYER VI3 ;
  RECT 2236.700 6.340 2236.900 6.540 ;
  LAYER VI3 ;
  RECT 2236.700 5.940 2236.900 6.140 ;
  LAYER VI3 ;
  RECT 2236.300 6.340 2236.500 6.540 ;
  LAYER VI3 ;
  RECT 2236.300 5.940 2236.500 6.140 ;
  LAYER VI3 ;
  RECT 2235.900 6.340 2236.100 6.540 ;
  LAYER VI3 ;
  RECT 2235.900 5.940 2236.100 6.140 ;
  LAYER VI3 ;
  RECT 2235.500 6.340 2235.700 6.540 ;
  LAYER VI3 ;
  RECT 2235.500 5.940 2235.700 6.140 ;
  LAYER VI3 ;
  RECT 2235.100 6.340 2235.300 6.540 ;
  LAYER VI3 ;
  RECT 2235.100 5.940 2235.300 6.140 ;
  LAYER VI3 ;
  RECT 2234.700 6.340 2234.900 6.540 ;
  LAYER VI3 ;
  RECT 2234.700 5.940 2234.900 6.140 ;
  LAYER VI3 ;
  RECT 2234.300 6.340 2234.500 6.540 ;
  LAYER VI3 ;
  RECT 2234.300 5.940 2234.500 6.140 ;
  LAYER VI3 ;
  RECT 2233.900 6.340 2234.100 6.540 ;
  LAYER VI3 ;
  RECT 2233.900 5.940 2234.100 6.140 ;
  LAYER VI3 ;
  RECT 2233.500 6.340 2233.700 6.540 ;
  LAYER VI3 ;
  RECT 2233.500 5.940 2233.700 6.140 ;
  LAYER VI3 ;
  RECT 2233.100 6.340 2233.300 6.540 ;
  LAYER VI3 ;
  RECT 2233.100 5.940 2233.300 6.140 ;
  LAYER VI3 ;
  RECT 2232.700 6.340 2232.900 6.540 ;
  LAYER VI3 ;
  RECT 2232.700 5.940 2232.900 6.140 ;
  LAYER VI3 ;
  RECT 2232.300 6.340 2232.500 6.540 ;
  LAYER VI3 ;
  RECT 2232.300 5.940 2232.500 6.140 ;
  LAYER VI3 ;
  RECT 2231.900 6.340 2232.100 6.540 ;
  LAYER VI3 ;
  RECT 2231.900 5.940 2232.100 6.140 ;
  LAYER VI3 ;
  RECT 2231.500 6.340 2231.700 6.540 ;
  LAYER VI3 ;
  RECT 2231.500 5.940 2231.700 6.140 ;
  LAYER VI3 ;
  RECT 2231.100 6.340 2231.300 6.540 ;
  LAYER VI3 ;
  RECT 2231.100 5.940 2231.300 6.140 ;
  LAYER VI3 ;
  RECT 2230.700 6.340 2230.900 6.540 ;
  LAYER VI3 ;
  RECT 2230.700 5.940 2230.900 6.140 ;
  LAYER VI3 ;
  RECT 2230.300 6.340 2230.500 6.540 ;
  LAYER VI3 ;
  RECT 2230.300 5.940 2230.500 6.140 ;
  LAYER VI3 ;
  RECT 2229.900 6.340 2230.100 6.540 ;
  LAYER VI3 ;
  RECT 2229.900 5.940 2230.100 6.140 ;
  LAYER VI3 ;
  RECT 2229.500 6.340 2229.700 6.540 ;
  LAYER VI3 ;
  RECT 2229.500 5.940 2229.700 6.140 ;
  LAYER VI3 ;
  RECT 2249.340 5.880 2257.340 6.740 ;
  LAYER VI3 ;
  RECT 2256.940 6.340 2257.140 6.540 ;
  LAYER VI3 ;
  RECT 2256.940 5.940 2257.140 6.140 ;
  LAYER VI3 ;
  RECT 2256.540 6.340 2256.740 6.540 ;
  LAYER VI3 ;
  RECT 2256.540 5.940 2256.740 6.140 ;
  LAYER VI3 ;
  RECT 2256.140 6.340 2256.340 6.540 ;
  LAYER VI3 ;
  RECT 2256.140 5.940 2256.340 6.140 ;
  LAYER VI3 ;
  RECT 2255.740 6.340 2255.940 6.540 ;
  LAYER VI3 ;
  RECT 2255.740 5.940 2255.940 6.140 ;
  LAYER VI3 ;
  RECT 2255.340 6.340 2255.540 6.540 ;
  LAYER VI3 ;
  RECT 2255.340 5.940 2255.540 6.140 ;
  LAYER VI3 ;
  RECT 2254.940 6.340 2255.140 6.540 ;
  LAYER VI3 ;
  RECT 2254.940 5.940 2255.140 6.140 ;
  LAYER VI3 ;
  RECT 2254.540 6.340 2254.740 6.540 ;
  LAYER VI3 ;
  RECT 2254.540 5.940 2254.740 6.140 ;
  LAYER VI3 ;
  RECT 2254.140 6.340 2254.340 6.540 ;
  LAYER VI3 ;
  RECT 2254.140 5.940 2254.340 6.140 ;
  LAYER VI3 ;
  RECT 2253.740 6.340 2253.940 6.540 ;
  LAYER VI3 ;
  RECT 2253.740 5.940 2253.940 6.140 ;
  LAYER VI3 ;
  RECT 2253.340 6.340 2253.540 6.540 ;
  LAYER VI3 ;
  RECT 2253.340 5.940 2253.540 6.140 ;
  LAYER VI3 ;
  RECT 2252.940 6.340 2253.140 6.540 ;
  LAYER VI3 ;
  RECT 2252.940 5.940 2253.140 6.140 ;
  LAYER VI3 ;
  RECT 2252.540 6.340 2252.740 6.540 ;
  LAYER VI3 ;
  RECT 2252.540 5.940 2252.740 6.140 ;
  LAYER VI3 ;
  RECT 2252.140 6.340 2252.340 6.540 ;
  LAYER VI3 ;
  RECT 2252.140 5.940 2252.340 6.140 ;
  LAYER VI3 ;
  RECT 2251.740 6.340 2251.940 6.540 ;
  LAYER VI3 ;
  RECT 2251.740 5.940 2251.940 6.140 ;
  LAYER VI3 ;
  RECT 2251.340 6.340 2251.540 6.540 ;
  LAYER VI3 ;
  RECT 2251.340 5.940 2251.540 6.140 ;
  LAYER VI3 ;
  RECT 2250.940 6.340 2251.140 6.540 ;
  LAYER VI3 ;
  RECT 2250.940 5.940 2251.140 6.140 ;
  LAYER VI3 ;
  RECT 2250.540 6.340 2250.740 6.540 ;
  LAYER VI3 ;
  RECT 2250.540 5.940 2250.740 6.140 ;
  LAYER VI3 ;
  RECT 2250.140 6.340 2250.340 6.540 ;
  LAYER VI3 ;
  RECT 2250.140 5.940 2250.340 6.140 ;
  LAYER VI3 ;
  RECT 2249.740 6.340 2249.940 6.540 ;
  LAYER VI3 ;
  RECT 2249.740 5.940 2249.940 6.140 ;
  LAYER VI3 ;
  RECT 2249.340 6.340 2249.540 6.540 ;
  LAYER VI3 ;
  RECT 2249.340 5.940 2249.540 6.140 ;
  LAYER VI3 ;
  RECT 2270.420 5.880 2278.420 6.740 ;
  LAYER VI3 ;
  RECT 2278.020 6.340 2278.220 6.540 ;
  LAYER VI3 ;
  RECT 2278.020 5.940 2278.220 6.140 ;
  LAYER VI3 ;
  RECT 2277.620 6.340 2277.820 6.540 ;
  LAYER VI3 ;
  RECT 2277.620 5.940 2277.820 6.140 ;
  LAYER VI3 ;
  RECT 2277.220 6.340 2277.420 6.540 ;
  LAYER VI3 ;
  RECT 2277.220 5.940 2277.420 6.140 ;
  LAYER VI3 ;
  RECT 2276.820 6.340 2277.020 6.540 ;
  LAYER VI3 ;
  RECT 2276.820 5.940 2277.020 6.140 ;
  LAYER VI3 ;
  RECT 2276.420 6.340 2276.620 6.540 ;
  LAYER VI3 ;
  RECT 2276.420 5.940 2276.620 6.140 ;
  LAYER VI3 ;
  RECT 2276.020 6.340 2276.220 6.540 ;
  LAYER VI3 ;
  RECT 2276.020 5.940 2276.220 6.140 ;
  LAYER VI3 ;
  RECT 2275.620 6.340 2275.820 6.540 ;
  LAYER VI3 ;
  RECT 2275.620 5.940 2275.820 6.140 ;
  LAYER VI3 ;
  RECT 2275.220 6.340 2275.420 6.540 ;
  LAYER VI3 ;
  RECT 2275.220 5.940 2275.420 6.140 ;
  LAYER VI3 ;
  RECT 2274.820 6.340 2275.020 6.540 ;
  LAYER VI3 ;
  RECT 2274.820 5.940 2275.020 6.140 ;
  LAYER VI3 ;
  RECT 2274.420 6.340 2274.620 6.540 ;
  LAYER VI3 ;
  RECT 2274.420 5.940 2274.620 6.140 ;
  LAYER VI3 ;
  RECT 2274.020 6.340 2274.220 6.540 ;
  LAYER VI3 ;
  RECT 2274.020 5.940 2274.220 6.140 ;
  LAYER VI3 ;
  RECT 2273.620 6.340 2273.820 6.540 ;
  LAYER VI3 ;
  RECT 2273.620 5.940 2273.820 6.140 ;
  LAYER VI3 ;
  RECT 2273.220 6.340 2273.420 6.540 ;
  LAYER VI3 ;
  RECT 2273.220 5.940 2273.420 6.140 ;
  LAYER VI3 ;
  RECT 2272.820 6.340 2273.020 6.540 ;
  LAYER VI3 ;
  RECT 2272.820 5.940 2273.020 6.140 ;
  LAYER VI3 ;
  RECT 2272.420 6.340 2272.620 6.540 ;
  LAYER VI3 ;
  RECT 2272.420 5.940 2272.620 6.140 ;
  LAYER VI3 ;
  RECT 2272.020 6.340 2272.220 6.540 ;
  LAYER VI3 ;
  RECT 2272.020 5.940 2272.220 6.140 ;
  LAYER VI3 ;
  RECT 2271.620 6.340 2271.820 6.540 ;
  LAYER VI3 ;
  RECT 2271.620 5.940 2271.820 6.140 ;
  LAYER VI3 ;
  RECT 2271.220 6.340 2271.420 6.540 ;
  LAYER VI3 ;
  RECT 2271.220 5.940 2271.420 6.140 ;
  LAYER VI3 ;
  RECT 2270.820 6.340 2271.020 6.540 ;
  LAYER VI3 ;
  RECT 2270.820 5.940 2271.020 6.140 ;
  LAYER VI3 ;
  RECT 2270.420 6.340 2270.620 6.540 ;
  LAYER VI3 ;
  RECT 2270.420 5.940 2270.620 6.140 ;
  LAYER VI3 ;
  RECT 2290.260 5.880 2298.260 6.740 ;
  LAYER VI3 ;
  RECT 2297.860 6.340 2298.060 6.540 ;
  LAYER VI3 ;
  RECT 2297.860 5.940 2298.060 6.140 ;
  LAYER VI3 ;
  RECT 2297.460 6.340 2297.660 6.540 ;
  LAYER VI3 ;
  RECT 2297.460 5.940 2297.660 6.140 ;
  LAYER VI3 ;
  RECT 2297.060 6.340 2297.260 6.540 ;
  LAYER VI3 ;
  RECT 2297.060 5.940 2297.260 6.140 ;
  LAYER VI3 ;
  RECT 2296.660 6.340 2296.860 6.540 ;
  LAYER VI3 ;
  RECT 2296.660 5.940 2296.860 6.140 ;
  LAYER VI3 ;
  RECT 2296.260 6.340 2296.460 6.540 ;
  LAYER VI3 ;
  RECT 2296.260 5.940 2296.460 6.140 ;
  LAYER VI3 ;
  RECT 2295.860 6.340 2296.060 6.540 ;
  LAYER VI3 ;
  RECT 2295.860 5.940 2296.060 6.140 ;
  LAYER VI3 ;
  RECT 2295.460 6.340 2295.660 6.540 ;
  LAYER VI3 ;
  RECT 2295.460 5.940 2295.660 6.140 ;
  LAYER VI3 ;
  RECT 2295.060 6.340 2295.260 6.540 ;
  LAYER VI3 ;
  RECT 2295.060 5.940 2295.260 6.140 ;
  LAYER VI3 ;
  RECT 2294.660 6.340 2294.860 6.540 ;
  LAYER VI3 ;
  RECT 2294.660 5.940 2294.860 6.140 ;
  LAYER VI3 ;
  RECT 2294.260 6.340 2294.460 6.540 ;
  LAYER VI3 ;
  RECT 2294.260 5.940 2294.460 6.140 ;
  LAYER VI3 ;
  RECT 2293.860 6.340 2294.060 6.540 ;
  LAYER VI3 ;
  RECT 2293.860 5.940 2294.060 6.140 ;
  LAYER VI3 ;
  RECT 2293.460 6.340 2293.660 6.540 ;
  LAYER VI3 ;
  RECT 2293.460 5.940 2293.660 6.140 ;
  LAYER VI3 ;
  RECT 2293.060 6.340 2293.260 6.540 ;
  LAYER VI3 ;
  RECT 2293.060 5.940 2293.260 6.140 ;
  LAYER VI3 ;
  RECT 2292.660 6.340 2292.860 6.540 ;
  LAYER VI3 ;
  RECT 2292.660 5.940 2292.860 6.140 ;
  LAYER VI3 ;
  RECT 2292.260 6.340 2292.460 6.540 ;
  LAYER VI3 ;
  RECT 2292.260 5.940 2292.460 6.140 ;
  LAYER VI3 ;
  RECT 2291.860 6.340 2292.060 6.540 ;
  LAYER VI3 ;
  RECT 2291.860 5.940 2292.060 6.140 ;
  LAYER VI3 ;
  RECT 2291.460 6.340 2291.660 6.540 ;
  LAYER VI3 ;
  RECT 2291.460 5.940 2291.660 6.140 ;
  LAYER VI3 ;
  RECT 2291.060 6.340 2291.260 6.540 ;
  LAYER VI3 ;
  RECT 2291.060 5.940 2291.260 6.140 ;
  LAYER VI3 ;
  RECT 2290.660 6.340 2290.860 6.540 ;
  LAYER VI3 ;
  RECT 2290.660 5.940 2290.860 6.140 ;
  LAYER VI3 ;
  RECT 2290.260 6.340 2290.460 6.540 ;
  LAYER VI3 ;
  RECT 2290.260 5.940 2290.460 6.140 ;
  LAYER VI3 ;
  RECT 2311.340 5.880 2319.340 6.740 ;
  LAYER VI3 ;
  RECT 2318.940 6.340 2319.140 6.540 ;
  LAYER VI3 ;
  RECT 2318.940 5.940 2319.140 6.140 ;
  LAYER VI3 ;
  RECT 2318.540 6.340 2318.740 6.540 ;
  LAYER VI3 ;
  RECT 2318.540 5.940 2318.740 6.140 ;
  LAYER VI3 ;
  RECT 2318.140 6.340 2318.340 6.540 ;
  LAYER VI3 ;
  RECT 2318.140 5.940 2318.340 6.140 ;
  LAYER VI3 ;
  RECT 2317.740 6.340 2317.940 6.540 ;
  LAYER VI3 ;
  RECT 2317.740 5.940 2317.940 6.140 ;
  LAYER VI3 ;
  RECT 2317.340 6.340 2317.540 6.540 ;
  LAYER VI3 ;
  RECT 2317.340 5.940 2317.540 6.140 ;
  LAYER VI3 ;
  RECT 2316.940 6.340 2317.140 6.540 ;
  LAYER VI3 ;
  RECT 2316.940 5.940 2317.140 6.140 ;
  LAYER VI3 ;
  RECT 2316.540 6.340 2316.740 6.540 ;
  LAYER VI3 ;
  RECT 2316.540 5.940 2316.740 6.140 ;
  LAYER VI3 ;
  RECT 2316.140 6.340 2316.340 6.540 ;
  LAYER VI3 ;
  RECT 2316.140 5.940 2316.340 6.140 ;
  LAYER VI3 ;
  RECT 2315.740 6.340 2315.940 6.540 ;
  LAYER VI3 ;
  RECT 2315.740 5.940 2315.940 6.140 ;
  LAYER VI3 ;
  RECT 2315.340 6.340 2315.540 6.540 ;
  LAYER VI3 ;
  RECT 2315.340 5.940 2315.540 6.140 ;
  LAYER VI3 ;
  RECT 2314.940 6.340 2315.140 6.540 ;
  LAYER VI3 ;
  RECT 2314.940 5.940 2315.140 6.140 ;
  LAYER VI3 ;
  RECT 2314.540 6.340 2314.740 6.540 ;
  LAYER VI3 ;
  RECT 2314.540 5.940 2314.740 6.140 ;
  LAYER VI3 ;
  RECT 2314.140 6.340 2314.340 6.540 ;
  LAYER VI3 ;
  RECT 2314.140 5.940 2314.340 6.140 ;
  LAYER VI3 ;
  RECT 2313.740 6.340 2313.940 6.540 ;
  LAYER VI3 ;
  RECT 2313.740 5.940 2313.940 6.140 ;
  LAYER VI3 ;
  RECT 2313.340 6.340 2313.540 6.540 ;
  LAYER VI3 ;
  RECT 2313.340 5.940 2313.540 6.140 ;
  LAYER VI3 ;
  RECT 2312.940 6.340 2313.140 6.540 ;
  LAYER VI3 ;
  RECT 2312.940 5.940 2313.140 6.140 ;
  LAYER VI3 ;
  RECT 2312.540 6.340 2312.740 6.540 ;
  LAYER VI3 ;
  RECT 2312.540 5.940 2312.740 6.140 ;
  LAYER VI3 ;
  RECT 2312.140 6.340 2312.340 6.540 ;
  LAYER VI3 ;
  RECT 2312.140 5.940 2312.340 6.140 ;
  LAYER VI3 ;
  RECT 2311.740 6.340 2311.940 6.540 ;
  LAYER VI3 ;
  RECT 2311.740 5.940 2311.940 6.140 ;
  LAYER VI3 ;
  RECT 2311.340 6.340 2311.540 6.540 ;
  LAYER VI3 ;
  RECT 2311.340 5.940 2311.540 6.140 ;
  LAYER VI3 ;
  RECT 2331.180 5.880 2339.180 6.740 ;
  LAYER VI3 ;
  RECT 2338.780 6.340 2338.980 6.540 ;
  LAYER VI3 ;
  RECT 2338.780 5.940 2338.980 6.140 ;
  LAYER VI3 ;
  RECT 2338.380 6.340 2338.580 6.540 ;
  LAYER VI3 ;
  RECT 2338.380 5.940 2338.580 6.140 ;
  LAYER VI3 ;
  RECT 2337.980 6.340 2338.180 6.540 ;
  LAYER VI3 ;
  RECT 2337.980 5.940 2338.180 6.140 ;
  LAYER VI3 ;
  RECT 2337.580 6.340 2337.780 6.540 ;
  LAYER VI3 ;
  RECT 2337.580 5.940 2337.780 6.140 ;
  LAYER VI3 ;
  RECT 2337.180 6.340 2337.380 6.540 ;
  LAYER VI3 ;
  RECT 2337.180 5.940 2337.380 6.140 ;
  LAYER VI3 ;
  RECT 2336.780 6.340 2336.980 6.540 ;
  LAYER VI3 ;
  RECT 2336.780 5.940 2336.980 6.140 ;
  LAYER VI3 ;
  RECT 2336.380 6.340 2336.580 6.540 ;
  LAYER VI3 ;
  RECT 2336.380 5.940 2336.580 6.140 ;
  LAYER VI3 ;
  RECT 2335.980 6.340 2336.180 6.540 ;
  LAYER VI3 ;
  RECT 2335.980 5.940 2336.180 6.140 ;
  LAYER VI3 ;
  RECT 2335.580 6.340 2335.780 6.540 ;
  LAYER VI3 ;
  RECT 2335.580 5.940 2335.780 6.140 ;
  LAYER VI3 ;
  RECT 2335.180 6.340 2335.380 6.540 ;
  LAYER VI3 ;
  RECT 2335.180 5.940 2335.380 6.140 ;
  LAYER VI3 ;
  RECT 2334.780 6.340 2334.980 6.540 ;
  LAYER VI3 ;
  RECT 2334.780 5.940 2334.980 6.140 ;
  LAYER VI3 ;
  RECT 2334.380 6.340 2334.580 6.540 ;
  LAYER VI3 ;
  RECT 2334.380 5.940 2334.580 6.140 ;
  LAYER VI3 ;
  RECT 2333.980 6.340 2334.180 6.540 ;
  LAYER VI3 ;
  RECT 2333.980 5.940 2334.180 6.140 ;
  LAYER VI3 ;
  RECT 2333.580 6.340 2333.780 6.540 ;
  LAYER VI3 ;
  RECT 2333.580 5.940 2333.780 6.140 ;
  LAYER VI3 ;
  RECT 2333.180 6.340 2333.380 6.540 ;
  LAYER VI3 ;
  RECT 2333.180 5.940 2333.380 6.140 ;
  LAYER VI3 ;
  RECT 2332.780 6.340 2332.980 6.540 ;
  LAYER VI3 ;
  RECT 2332.780 5.940 2332.980 6.140 ;
  LAYER VI3 ;
  RECT 2332.380 6.340 2332.580 6.540 ;
  LAYER VI3 ;
  RECT 2332.380 5.940 2332.580 6.140 ;
  LAYER VI3 ;
  RECT 2331.980 6.340 2332.180 6.540 ;
  LAYER VI3 ;
  RECT 2331.980 5.940 2332.180 6.140 ;
  LAYER VI3 ;
  RECT 2331.580 6.340 2331.780 6.540 ;
  LAYER VI3 ;
  RECT 2331.580 5.940 2331.780 6.140 ;
  LAYER VI3 ;
  RECT 2331.180 6.340 2331.380 6.540 ;
  LAYER VI3 ;
  RECT 2331.180 5.940 2331.380 6.140 ;
  LAYER VI3 ;
  RECT 2352.260 5.880 2360.260 6.740 ;
  LAYER VI3 ;
  RECT 2359.860 6.340 2360.060 6.540 ;
  LAYER VI3 ;
  RECT 2359.860 5.940 2360.060 6.140 ;
  LAYER VI3 ;
  RECT 2359.460 6.340 2359.660 6.540 ;
  LAYER VI3 ;
  RECT 2359.460 5.940 2359.660 6.140 ;
  LAYER VI3 ;
  RECT 2359.060 6.340 2359.260 6.540 ;
  LAYER VI3 ;
  RECT 2359.060 5.940 2359.260 6.140 ;
  LAYER VI3 ;
  RECT 2358.660 6.340 2358.860 6.540 ;
  LAYER VI3 ;
  RECT 2358.660 5.940 2358.860 6.140 ;
  LAYER VI3 ;
  RECT 2358.260 6.340 2358.460 6.540 ;
  LAYER VI3 ;
  RECT 2358.260 5.940 2358.460 6.140 ;
  LAYER VI3 ;
  RECT 2357.860 6.340 2358.060 6.540 ;
  LAYER VI3 ;
  RECT 2357.860 5.940 2358.060 6.140 ;
  LAYER VI3 ;
  RECT 2357.460 6.340 2357.660 6.540 ;
  LAYER VI3 ;
  RECT 2357.460 5.940 2357.660 6.140 ;
  LAYER VI3 ;
  RECT 2357.060 6.340 2357.260 6.540 ;
  LAYER VI3 ;
  RECT 2357.060 5.940 2357.260 6.140 ;
  LAYER VI3 ;
  RECT 2356.660 6.340 2356.860 6.540 ;
  LAYER VI3 ;
  RECT 2356.660 5.940 2356.860 6.140 ;
  LAYER VI3 ;
  RECT 2356.260 6.340 2356.460 6.540 ;
  LAYER VI3 ;
  RECT 2356.260 5.940 2356.460 6.140 ;
  LAYER VI3 ;
  RECT 2355.860 6.340 2356.060 6.540 ;
  LAYER VI3 ;
  RECT 2355.860 5.940 2356.060 6.140 ;
  LAYER VI3 ;
  RECT 2355.460 6.340 2355.660 6.540 ;
  LAYER VI3 ;
  RECT 2355.460 5.940 2355.660 6.140 ;
  LAYER VI3 ;
  RECT 2355.060 6.340 2355.260 6.540 ;
  LAYER VI3 ;
  RECT 2355.060 5.940 2355.260 6.140 ;
  LAYER VI3 ;
  RECT 2354.660 6.340 2354.860 6.540 ;
  LAYER VI3 ;
  RECT 2354.660 5.940 2354.860 6.140 ;
  LAYER VI3 ;
  RECT 2354.260 6.340 2354.460 6.540 ;
  LAYER VI3 ;
  RECT 2354.260 5.940 2354.460 6.140 ;
  LAYER VI3 ;
  RECT 2353.860 6.340 2354.060 6.540 ;
  LAYER VI3 ;
  RECT 2353.860 5.940 2354.060 6.140 ;
  LAYER VI3 ;
  RECT 2353.460 6.340 2353.660 6.540 ;
  LAYER VI3 ;
  RECT 2353.460 5.940 2353.660 6.140 ;
  LAYER VI3 ;
  RECT 2353.060 6.340 2353.260 6.540 ;
  LAYER VI3 ;
  RECT 2353.060 5.940 2353.260 6.140 ;
  LAYER VI3 ;
  RECT 2352.660 6.340 2352.860 6.540 ;
  LAYER VI3 ;
  RECT 2352.660 5.940 2352.860 6.140 ;
  LAYER VI3 ;
  RECT 2352.260 6.340 2352.460 6.540 ;
  LAYER VI3 ;
  RECT 2352.260 5.940 2352.460 6.140 ;
  LAYER VI3 ;
  RECT 2372.100 5.880 2380.100 6.740 ;
  LAYER VI3 ;
  RECT 2379.700 6.340 2379.900 6.540 ;
  LAYER VI3 ;
  RECT 2379.700 5.940 2379.900 6.140 ;
  LAYER VI3 ;
  RECT 2379.300 6.340 2379.500 6.540 ;
  LAYER VI3 ;
  RECT 2379.300 5.940 2379.500 6.140 ;
  LAYER VI3 ;
  RECT 2378.900 6.340 2379.100 6.540 ;
  LAYER VI3 ;
  RECT 2378.900 5.940 2379.100 6.140 ;
  LAYER VI3 ;
  RECT 2378.500 6.340 2378.700 6.540 ;
  LAYER VI3 ;
  RECT 2378.500 5.940 2378.700 6.140 ;
  LAYER VI3 ;
  RECT 2378.100 6.340 2378.300 6.540 ;
  LAYER VI3 ;
  RECT 2378.100 5.940 2378.300 6.140 ;
  LAYER VI3 ;
  RECT 2377.700 6.340 2377.900 6.540 ;
  LAYER VI3 ;
  RECT 2377.700 5.940 2377.900 6.140 ;
  LAYER VI3 ;
  RECT 2377.300 6.340 2377.500 6.540 ;
  LAYER VI3 ;
  RECT 2377.300 5.940 2377.500 6.140 ;
  LAYER VI3 ;
  RECT 2376.900 6.340 2377.100 6.540 ;
  LAYER VI3 ;
  RECT 2376.900 5.940 2377.100 6.140 ;
  LAYER VI3 ;
  RECT 2376.500 6.340 2376.700 6.540 ;
  LAYER VI3 ;
  RECT 2376.500 5.940 2376.700 6.140 ;
  LAYER VI3 ;
  RECT 2376.100 6.340 2376.300 6.540 ;
  LAYER VI3 ;
  RECT 2376.100 5.940 2376.300 6.140 ;
  LAYER VI3 ;
  RECT 2375.700 6.340 2375.900 6.540 ;
  LAYER VI3 ;
  RECT 2375.700 5.940 2375.900 6.140 ;
  LAYER VI3 ;
  RECT 2375.300 6.340 2375.500 6.540 ;
  LAYER VI3 ;
  RECT 2375.300 5.940 2375.500 6.140 ;
  LAYER VI3 ;
  RECT 2374.900 6.340 2375.100 6.540 ;
  LAYER VI3 ;
  RECT 2374.900 5.940 2375.100 6.140 ;
  LAYER VI3 ;
  RECT 2374.500 6.340 2374.700 6.540 ;
  LAYER VI3 ;
  RECT 2374.500 5.940 2374.700 6.140 ;
  LAYER VI3 ;
  RECT 2374.100 6.340 2374.300 6.540 ;
  LAYER VI3 ;
  RECT 2374.100 5.940 2374.300 6.140 ;
  LAYER VI3 ;
  RECT 2373.700 6.340 2373.900 6.540 ;
  LAYER VI3 ;
  RECT 2373.700 5.940 2373.900 6.140 ;
  LAYER VI3 ;
  RECT 2373.300 6.340 2373.500 6.540 ;
  LAYER VI3 ;
  RECT 2373.300 5.940 2373.500 6.140 ;
  LAYER VI3 ;
  RECT 2372.900 6.340 2373.100 6.540 ;
  LAYER VI3 ;
  RECT 2372.900 5.940 2373.100 6.140 ;
  LAYER VI3 ;
  RECT 2372.500 6.340 2372.700 6.540 ;
  LAYER VI3 ;
  RECT 2372.500 5.940 2372.700 6.140 ;
  LAYER VI3 ;
  RECT 2372.100 6.340 2372.300 6.540 ;
  LAYER VI3 ;
  RECT 2372.100 5.940 2372.300 6.140 ;
  LAYER VI3 ;
  RECT 2393.180 5.880 2401.180 6.740 ;
  LAYER VI3 ;
  RECT 2400.780 6.340 2400.980 6.540 ;
  LAYER VI3 ;
  RECT 2400.780 5.940 2400.980 6.140 ;
  LAYER VI3 ;
  RECT 2400.380 6.340 2400.580 6.540 ;
  LAYER VI3 ;
  RECT 2400.380 5.940 2400.580 6.140 ;
  LAYER VI3 ;
  RECT 2399.980 6.340 2400.180 6.540 ;
  LAYER VI3 ;
  RECT 2399.980 5.940 2400.180 6.140 ;
  LAYER VI3 ;
  RECT 2399.580 6.340 2399.780 6.540 ;
  LAYER VI3 ;
  RECT 2399.580 5.940 2399.780 6.140 ;
  LAYER VI3 ;
  RECT 2399.180 6.340 2399.380 6.540 ;
  LAYER VI3 ;
  RECT 2399.180 5.940 2399.380 6.140 ;
  LAYER VI3 ;
  RECT 2398.780 6.340 2398.980 6.540 ;
  LAYER VI3 ;
  RECT 2398.780 5.940 2398.980 6.140 ;
  LAYER VI3 ;
  RECT 2398.380 6.340 2398.580 6.540 ;
  LAYER VI3 ;
  RECT 2398.380 5.940 2398.580 6.140 ;
  LAYER VI3 ;
  RECT 2397.980 6.340 2398.180 6.540 ;
  LAYER VI3 ;
  RECT 2397.980 5.940 2398.180 6.140 ;
  LAYER VI3 ;
  RECT 2397.580 6.340 2397.780 6.540 ;
  LAYER VI3 ;
  RECT 2397.580 5.940 2397.780 6.140 ;
  LAYER VI3 ;
  RECT 2397.180 6.340 2397.380 6.540 ;
  LAYER VI3 ;
  RECT 2397.180 5.940 2397.380 6.140 ;
  LAYER VI3 ;
  RECT 2396.780 6.340 2396.980 6.540 ;
  LAYER VI3 ;
  RECT 2396.780 5.940 2396.980 6.140 ;
  LAYER VI3 ;
  RECT 2396.380 6.340 2396.580 6.540 ;
  LAYER VI3 ;
  RECT 2396.380 5.940 2396.580 6.140 ;
  LAYER VI3 ;
  RECT 2395.980 6.340 2396.180 6.540 ;
  LAYER VI3 ;
  RECT 2395.980 5.940 2396.180 6.140 ;
  LAYER VI3 ;
  RECT 2395.580 6.340 2395.780 6.540 ;
  LAYER VI3 ;
  RECT 2395.580 5.940 2395.780 6.140 ;
  LAYER VI3 ;
  RECT 2395.180 6.340 2395.380 6.540 ;
  LAYER VI3 ;
  RECT 2395.180 5.940 2395.380 6.140 ;
  LAYER VI3 ;
  RECT 2394.780 6.340 2394.980 6.540 ;
  LAYER VI3 ;
  RECT 2394.780 5.940 2394.980 6.140 ;
  LAYER VI3 ;
  RECT 2394.380 6.340 2394.580 6.540 ;
  LAYER VI3 ;
  RECT 2394.380 5.940 2394.580 6.140 ;
  LAYER VI3 ;
  RECT 2393.980 6.340 2394.180 6.540 ;
  LAYER VI3 ;
  RECT 2393.980 5.940 2394.180 6.140 ;
  LAYER VI3 ;
  RECT 2393.580 6.340 2393.780 6.540 ;
  LAYER VI3 ;
  RECT 2393.580 5.940 2393.780 6.140 ;
  LAYER VI3 ;
  RECT 2393.180 6.340 2393.380 6.540 ;
  LAYER VI3 ;
  RECT 2393.180 5.940 2393.380 6.140 ;
  LAYER VI3 ;
  RECT 2413.020 5.880 2421.020 6.740 ;
  LAYER VI3 ;
  RECT 2420.620 6.340 2420.820 6.540 ;
  LAYER VI3 ;
  RECT 2420.620 5.940 2420.820 6.140 ;
  LAYER VI3 ;
  RECT 2420.220 6.340 2420.420 6.540 ;
  LAYER VI3 ;
  RECT 2420.220 5.940 2420.420 6.140 ;
  LAYER VI3 ;
  RECT 2419.820 6.340 2420.020 6.540 ;
  LAYER VI3 ;
  RECT 2419.820 5.940 2420.020 6.140 ;
  LAYER VI3 ;
  RECT 2419.420 6.340 2419.620 6.540 ;
  LAYER VI3 ;
  RECT 2419.420 5.940 2419.620 6.140 ;
  LAYER VI3 ;
  RECT 2419.020 6.340 2419.220 6.540 ;
  LAYER VI3 ;
  RECT 2419.020 5.940 2419.220 6.140 ;
  LAYER VI3 ;
  RECT 2418.620 6.340 2418.820 6.540 ;
  LAYER VI3 ;
  RECT 2418.620 5.940 2418.820 6.140 ;
  LAYER VI3 ;
  RECT 2418.220 6.340 2418.420 6.540 ;
  LAYER VI3 ;
  RECT 2418.220 5.940 2418.420 6.140 ;
  LAYER VI3 ;
  RECT 2417.820 6.340 2418.020 6.540 ;
  LAYER VI3 ;
  RECT 2417.820 5.940 2418.020 6.140 ;
  LAYER VI3 ;
  RECT 2417.420 6.340 2417.620 6.540 ;
  LAYER VI3 ;
  RECT 2417.420 5.940 2417.620 6.140 ;
  LAYER VI3 ;
  RECT 2417.020 6.340 2417.220 6.540 ;
  LAYER VI3 ;
  RECT 2417.020 5.940 2417.220 6.140 ;
  LAYER VI3 ;
  RECT 2416.620 6.340 2416.820 6.540 ;
  LAYER VI3 ;
  RECT 2416.620 5.940 2416.820 6.140 ;
  LAYER VI3 ;
  RECT 2416.220 6.340 2416.420 6.540 ;
  LAYER VI3 ;
  RECT 2416.220 5.940 2416.420 6.140 ;
  LAYER VI3 ;
  RECT 2415.820 6.340 2416.020 6.540 ;
  LAYER VI3 ;
  RECT 2415.820 5.940 2416.020 6.140 ;
  LAYER VI3 ;
  RECT 2415.420 6.340 2415.620 6.540 ;
  LAYER VI3 ;
  RECT 2415.420 5.940 2415.620 6.140 ;
  LAYER VI3 ;
  RECT 2415.020 6.340 2415.220 6.540 ;
  LAYER VI3 ;
  RECT 2415.020 5.940 2415.220 6.140 ;
  LAYER VI3 ;
  RECT 2414.620 6.340 2414.820 6.540 ;
  LAYER VI3 ;
  RECT 2414.620 5.940 2414.820 6.140 ;
  LAYER VI3 ;
  RECT 2414.220 6.340 2414.420 6.540 ;
  LAYER VI3 ;
  RECT 2414.220 5.940 2414.420 6.140 ;
  LAYER VI3 ;
  RECT 2413.820 6.340 2414.020 6.540 ;
  LAYER VI3 ;
  RECT 2413.820 5.940 2414.020 6.140 ;
  LAYER VI3 ;
  RECT 2413.420 6.340 2413.620 6.540 ;
  LAYER VI3 ;
  RECT 2413.420 5.940 2413.620 6.140 ;
  LAYER VI3 ;
  RECT 2413.020 6.340 2413.220 6.540 ;
  LAYER VI3 ;
  RECT 2413.020 5.940 2413.220 6.140 ;
  LAYER VI3 ;
  RECT 2434.100 5.880 2442.100 6.740 ;
  LAYER VI3 ;
  RECT 2441.700 6.340 2441.900 6.540 ;
  LAYER VI3 ;
  RECT 2441.700 5.940 2441.900 6.140 ;
  LAYER VI3 ;
  RECT 2441.300 6.340 2441.500 6.540 ;
  LAYER VI3 ;
  RECT 2441.300 5.940 2441.500 6.140 ;
  LAYER VI3 ;
  RECT 2440.900 6.340 2441.100 6.540 ;
  LAYER VI3 ;
  RECT 2440.900 5.940 2441.100 6.140 ;
  LAYER VI3 ;
  RECT 2440.500 6.340 2440.700 6.540 ;
  LAYER VI3 ;
  RECT 2440.500 5.940 2440.700 6.140 ;
  LAYER VI3 ;
  RECT 2440.100 6.340 2440.300 6.540 ;
  LAYER VI3 ;
  RECT 2440.100 5.940 2440.300 6.140 ;
  LAYER VI3 ;
  RECT 2439.700 6.340 2439.900 6.540 ;
  LAYER VI3 ;
  RECT 2439.700 5.940 2439.900 6.140 ;
  LAYER VI3 ;
  RECT 2439.300 6.340 2439.500 6.540 ;
  LAYER VI3 ;
  RECT 2439.300 5.940 2439.500 6.140 ;
  LAYER VI3 ;
  RECT 2438.900 6.340 2439.100 6.540 ;
  LAYER VI3 ;
  RECT 2438.900 5.940 2439.100 6.140 ;
  LAYER VI3 ;
  RECT 2438.500 6.340 2438.700 6.540 ;
  LAYER VI3 ;
  RECT 2438.500 5.940 2438.700 6.140 ;
  LAYER VI3 ;
  RECT 2438.100 6.340 2438.300 6.540 ;
  LAYER VI3 ;
  RECT 2438.100 5.940 2438.300 6.140 ;
  LAYER VI3 ;
  RECT 2437.700 6.340 2437.900 6.540 ;
  LAYER VI3 ;
  RECT 2437.700 5.940 2437.900 6.140 ;
  LAYER VI3 ;
  RECT 2437.300 6.340 2437.500 6.540 ;
  LAYER VI3 ;
  RECT 2437.300 5.940 2437.500 6.140 ;
  LAYER VI3 ;
  RECT 2436.900 6.340 2437.100 6.540 ;
  LAYER VI3 ;
  RECT 2436.900 5.940 2437.100 6.140 ;
  LAYER VI3 ;
  RECT 2436.500 6.340 2436.700 6.540 ;
  LAYER VI3 ;
  RECT 2436.500 5.940 2436.700 6.140 ;
  LAYER VI3 ;
  RECT 2436.100 6.340 2436.300 6.540 ;
  LAYER VI3 ;
  RECT 2436.100 5.940 2436.300 6.140 ;
  LAYER VI3 ;
  RECT 2435.700 6.340 2435.900 6.540 ;
  LAYER VI3 ;
  RECT 2435.700 5.940 2435.900 6.140 ;
  LAYER VI3 ;
  RECT 2435.300 6.340 2435.500 6.540 ;
  LAYER VI3 ;
  RECT 2435.300 5.940 2435.500 6.140 ;
  LAYER VI3 ;
  RECT 2434.900 6.340 2435.100 6.540 ;
  LAYER VI3 ;
  RECT 2434.900 5.940 2435.100 6.140 ;
  LAYER VI3 ;
  RECT 2434.500 6.340 2434.700 6.540 ;
  LAYER VI3 ;
  RECT 2434.500 5.940 2434.700 6.140 ;
  LAYER VI3 ;
  RECT 2434.100 6.340 2434.300 6.540 ;
  LAYER VI3 ;
  RECT 2434.100 5.940 2434.300 6.140 ;
  LAYER VI3 ;
  RECT 2453.940 5.880 2461.940 6.740 ;
  LAYER VI3 ;
  RECT 2461.540 6.340 2461.740 6.540 ;
  LAYER VI3 ;
  RECT 2461.540 5.940 2461.740 6.140 ;
  LAYER VI3 ;
  RECT 2461.140 6.340 2461.340 6.540 ;
  LAYER VI3 ;
  RECT 2461.140 5.940 2461.340 6.140 ;
  LAYER VI3 ;
  RECT 2460.740 6.340 2460.940 6.540 ;
  LAYER VI3 ;
  RECT 2460.740 5.940 2460.940 6.140 ;
  LAYER VI3 ;
  RECT 2460.340 6.340 2460.540 6.540 ;
  LAYER VI3 ;
  RECT 2460.340 5.940 2460.540 6.140 ;
  LAYER VI3 ;
  RECT 2459.940 6.340 2460.140 6.540 ;
  LAYER VI3 ;
  RECT 2459.940 5.940 2460.140 6.140 ;
  LAYER VI3 ;
  RECT 2459.540 6.340 2459.740 6.540 ;
  LAYER VI3 ;
  RECT 2459.540 5.940 2459.740 6.140 ;
  LAYER VI3 ;
  RECT 2459.140 6.340 2459.340 6.540 ;
  LAYER VI3 ;
  RECT 2459.140 5.940 2459.340 6.140 ;
  LAYER VI3 ;
  RECT 2458.740 6.340 2458.940 6.540 ;
  LAYER VI3 ;
  RECT 2458.740 5.940 2458.940 6.140 ;
  LAYER VI3 ;
  RECT 2458.340 6.340 2458.540 6.540 ;
  LAYER VI3 ;
  RECT 2458.340 5.940 2458.540 6.140 ;
  LAYER VI3 ;
  RECT 2457.940 6.340 2458.140 6.540 ;
  LAYER VI3 ;
  RECT 2457.940 5.940 2458.140 6.140 ;
  LAYER VI3 ;
  RECT 2457.540 6.340 2457.740 6.540 ;
  LAYER VI3 ;
  RECT 2457.540 5.940 2457.740 6.140 ;
  LAYER VI3 ;
  RECT 2457.140 6.340 2457.340 6.540 ;
  LAYER VI3 ;
  RECT 2457.140 5.940 2457.340 6.140 ;
  LAYER VI3 ;
  RECT 2456.740 6.340 2456.940 6.540 ;
  LAYER VI3 ;
  RECT 2456.740 5.940 2456.940 6.140 ;
  LAYER VI3 ;
  RECT 2456.340 6.340 2456.540 6.540 ;
  LAYER VI3 ;
  RECT 2456.340 5.940 2456.540 6.140 ;
  LAYER VI3 ;
  RECT 2455.940 6.340 2456.140 6.540 ;
  LAYER VI3 ;
  RECT 2455.940 5.940 2456.140 6.140 ;
  LAYER VI3 ;
  RECT 2455.540 6.340 2455.740 6.540 ;
  LAYER VI3 ;
  RECT 2455.540 5.940 2455.740 6.140 ;
  LAYER VI3 ;
  RECT 2455.140 6.340 2455.340 6.540 ;
  LAYER VI3 ;
  RECT 2455.140 5.940 2455.340 6.140 ;
  LAYER VI3 ;
  RECT 2454.740 6.340 2454.940 6.540 ;
  LAYER VI3 ;
  RECT 2454.740 5.940 2454.940 6.140 ;
  LAYER VI3 ;
  RECT 2454.340 6.340 2454.540 6.540 ;
  LAYER VI3 ;
  RECT 2454.340 5.940 2454.540 6.140 ;
  LAYER VI3 ;
  RECT 2453.940 6.340 2454.140 6.540 ;
  LAYER VI3 ;
  RECT 2453.940 5.940 2454.140 6.140 ;
  LAYER VI3 ;
  RECT 2475.020 5.880 2483.020 6.740 ;
  LAYER VI3 ;
  RECT 2482.620 6.340 2482.820 6.540 ;
  LAYER VI3 ;
  RECT 2482.620 5.940 2482.820 6.140 ;
  LAYER VI3 ;
  RECT 2482.220 6.340 2482.420 6.540 ;
  LAYER VI3 ;
  RECT 2482.220 5.940 2482.420 6.140 ;
  LAYER VI3 ;
  RECT 2481.820 6.340 2482.020 6.540 ;
  LAYER VI3 ;
  RECT 2481.820 5.940 2482.020 6.140 ;
  LAYER VI3 ;
  RECT 2481.420 6.340 2481.620 6.540 ;
  LAYER VI3 ;
  RECT 2481.420 5.940 2481.620 6.140 ;
  LAYER VI3 ;
  RECT 2481.020 6.340 2481.220 6.540 ;
  LAYER VI3 ;
  RECT 2481.020 5.940 2481.220 6.140 ;
  LAYER VI3 ;
  RECT 2480.620 6.340 2480.820 6.540 ;
  LAYER VI3 ;
  RECT 2480.620 5.940 2480.820 6.140 ;
  LAYER VI3 ;
  RECT 2480.220 6.340 2480.420 6.540 ;
  LAYER VI3 ;
  RECT 2480.220 5.940 2480.420 6.140 ;
  LAYER VI3 ;
  RECT 2479.820 6.340 2480.020 6.540 ;
  LAYER VI3 ;
  RECT 2479.820 5.940 2480.020 6.140 ;
  LAYER VI3 ;
  RECT 2479.420 6.340 2479.620 6.540 ;
  LAYER VI3 ;
  RECT 2479.420 5.940 2479.620 6.140 ;
  LAYER VI3 ;
  RECT 2479.020 6.340 2479.220 6.540 ;
  LAYER VI3 ;
  RECT 2479.020 5.940 2479.220 6.140 ;
  LAYER VI3 ;
  RECT 2478.620 6.340 2478.820 6.540 ;
  LAYER VI3 ;
  RECT 2478.620 5.940 2478.820 6.140 ;
  LAYER VI3 ;
  RECT 2478.220 6.340 2478.420 6.540 ;
  LAYER VI3 ;
  RECT 2478.220 5.940 2478.420 6.140 ;
  LAYER VI3 ;
  RECT 2477.820 6.340 2478.020 6.540 ;
  LAYER VI3 ;
  RECT 2477.820 5.940 2478.020 6.140 ;
  LAYER VI3 ;
  RECT 2477.420 6.340 2477.620 6.540 ;
  LAYER VI3 ;
  RECT 2477.420 5.940 2477.620 6.140 ;
  LAYER VI3 ;
  RECT 2477.020 6.340 2477.220 6.540 ;
  LAYER VI3 ;
  RECT 2477.020 5.940 2477.220 6.140 ;
  LAYER VI3 ;
  RECT 2476.620 6.340 2476.820 6.540 ;
  LAYER VI3 ;
  RECT 2476.620 5.940 2476.820 6.140 ;
  LAYER VI3 ;
  RECT 2476.220 6.340 2476.420 6.540 ;
  LAYER VI3 ;
  RECT 2476.220 5.940 2476.420 6.140 ;
  LAYER VI3 ;
  RECT 2475.820 6.340 2476.020 6.540 ;
  LAYER VI3 ;
  RECT 2475.820 5.940 2476.020 6.140 ;
  LAYER VI3 ;
  RECT 2475.420 6.340 2475.620 6.540 ;
  LAYER VI3 ;
  RECT 2475.420 5.940 2475.620 6.140 ;
  LAYER VI3 ;
  RECT 2475.020 6.340 2475.220 6.540 ;
  LAYER VI3 ;
  RECT 2475.020 5.940 2475.220 6.140 ;
  LAYER VI3 ;
  RECT 2494.860 5.880 2502.860 6.740 ;
  LAYER VI3 ;
  RECT 2502.460 6.340 2502.660 6.540 ;
  LAYER VI3 ;
  RECT 2502.460 5.940 2502.660 6.140 ;
  LAYER VI3 ;
  RECT 2502.060 6.340 2502.260 6.540 ;
  LAYER VI3 ;
  RECT 2502.060 5.940 2502.260 6.140 ;
  LAYER VI3 ;
  RECT 2501.660 6.340 2501.860 6.540 ;
  LAYER VI3 ;
  RECT 2501.660 5.940 2501.860 6.140 ;
  LAYER VI3 ;
  RECT 2501.260 6.340 2501.460 6.540 ;
  LAYER VI3 ;
  RECT 2501.260 5.940 2501.460 6.140 ;
  LAYER VI3 ;
  RECT 2500.860 6.340 2501.060 6.540 ;
  LAYER VI3 ;
  RECT 2500.860 5.940 2501.060 6.140 ;
  LAYER VI3 ;
  RECT 2500.460 6.340 2500.660 6.540 ;
  LAYER VI3 ;
  RECT 2500.460 5.940 2500.660 6.140 ;
  LAYER VI3 ;
  RECT 2500.060 6.340 2500.260 6.540 ;
  LAYER VI3 ;
  RECT 2500.060 5.940 2500.260 6.140 ;
  LAYER VI3 ;
  RECT 2499.660 6.340 2499.860 6.540 ;
  LAYER VI3 ;
  RECT 2499.660 5.940 2499.860 6.140 ;
  LAYER VI3 ;
  RECT 2499.260 6.340 2499.460 6.540 ;
  LAYER VI3 ;
  RECT 2499.260 5.940 2499.460 6.140 ;
  LAYER VI3 ;
  RECT 2498.860 6.340 2499.060 6.540 ;
  LAYER VI3 ;
  RECT 2498.860 5.940 2499.060 6.140 ;
  LAYER VI3 ;
  RECT 2498.460 6.340 2498.660 6.540 ;
  LAYER VI3 ;
  RECT 2498.460 5.940 2498.660 6.140 ;
  LAYER VI3 ;
  RECT 2498.060 6.340 2498.260 6.540 ;
  LAYER VI3 ;
  RECT 2498.060 5.940 2498.260 6.140 ;
  LAYER VI3 ;
  RECT 2497.660 6.340 2497.860 6.540 ;
  LAYER VI3 ;
  RECT 2497.660 5.940 2497.860 6.140 ;
  LAYER VI3 ;
  RECT 2497.260 6.340 2497.460 6.540 ;
  LAYER VI3 ;
  RECT 2497.260 5.940 2497.460 6.140 ;
  LAYER VI3 ;
  RECT 2496.860 6.340 2497.060 6.540 ;
  LAYER VI3 ;
  RECT 2496.860 5.940 2497.060 6.140 ;
  LAYER VI3 ;
  RECT 2496.460 6.340 2496.660 6.540 ;
  LAYER VI3 ;
  RECT 2496.460 5.940 2496.660 6.140 ;
  LAYER VI3 ;
  RECT 2496.060 6.340 2496.260 6.540 ;
  LAYER VI3 ;
  RECT 2496.060 5.940 2496.260 6.140 ;
  LAYER VI3 ;
  RECT 2495.660 6.340 2495.860 6.540 ;
  LAYER VI3 ;
  RECT 2495.660 5.940 2495.860 6.140 ;
  LAYER VI3 ;
  RECT 2495.260 6.340 2495.460 6.540 ;
  LAYER VI3 ;
  RECT 2495.260 5.940 2495.460 6.140 ;
  LAYER VI3 ;
  RECT 2494.860 6.340 2495.060 6.540 ;
  LAYER VI3 ;
  RECT 2494.860 5.940 2495.060 6.140 ;
  LAYER VI3 ;
  RECT 2515.940 5.880 2523.940 6.740 ;
  LAYER VI3 ;
  RECT 2523.540 6.340 2523.740 6.540 ;
  LAYER VI3 ;
  RECT 2523.540 5.940 2523.740 6.140 ;
  LAYER VI3 ;
  RECT 2523.140 6.340 2523.340 6.540 ;
  LAYER VI3 ;
  RECT 2523.140 5.940 2523.340 6.140 ;
  LAYER VI3 ;
  RECT 2522.740 6.340 2522.940 6.540 ;
  LAYER VI3 ;
  RECT 2522.740 5.940 2522.940 6.140 ;
  LAYER VI3 ;
  RECT 2522.340 6.340 2522.540 6.540 ;
  LAYER VI3 ;
  RECT 2522.340 5.940 2522.540 6.140 ;
  LAYER VI3 ;
  RECT 2521.940 6.340 2522.140 6.540 ;
  LAYER VI3 ;
  RECT 2521.940 5.940 2522.140 6.140 ;
  LAYER VI3 ;
  RECT 2521.540 6.340 2521.740 6.540 ;
  LAYER VI3 ;
  RECT 2521.540 5.940 2521.740 6.140 ;
  LAYER VI3 ;
  RECT 2521.140 6.340 2521.340 6.540 ;
  LAYER VI3 ;
  RECT 2521.140 5.940 2521.340 6.140 ;
  LAYER VI3 ;
  RECT 2520.740 6.340 2520.940 6.540 ;
  LAYER VI3 ;
  RECT 2520.740 5.940 2520.940 6.140 ;
  LAYER VI3 ;
  RECT 2520.340 6.340 2520.540 6.540 ;
  LAYER VI3 ;
  RECT 2520.340 5.940 2520.540 6.140 ;
  LAYER VI3 ;
  RECT 2519.940 6.340 2520.140 6.540 ;
  LAYER VI3 ;
  RECT 2519.940 5.940 2520.140 6.140 ;
  LAYER VI3 ;
  RECT 2519.540 6.340 2519.740 6.540 ;
  LAYER VI3 ;
  RECT 2519.540 5.940 2519.740 6.140 ;
  LAYER VI3 ;
  RECT 2519.140 6.340 2519.340 6.540 ;
  LAYER VI3 ;
  RECT 2519.140 5.940 2519.340 6.140 ;
  LAYER VI3 ;
  RECT 2518.740 6.340 2518.940 6.540 ;
  LAYER VI3 ;
  RECT 2518.740 5.940 2518.940 6.140 ;
  LAYER VI3 ;
  RECT 2518.340 6.340 2518.540 6.540 ;
  LAYER VI3 ;
  RECT 2518.340 5.940 2518.540 6.140 ;
  LAYER VI3 ;
  RECT 2517.940 6.340 2518.140 6.540 ;
  LAYER VI3 ;
  RECT 2517.940 5.940 2518.140 6.140 ;
  LAYER VI3 ;
  RECT 2517.540 6.340 2517.740 6.540 ;
  LAYER VI3 ;
  RECT 2517.540 5.940 2517.740 6.140 ;
  LAYER VI3 ;
  RECT 2517.140 6.340 2517.340 6.540 ;
  LAYER VI3 ;
  RECT 2517.140 5.940 2517.340 6.140 ;
  LAYER VI3 ;
  RECT 2516.740 6.340 2516.940 6.540 ;
  LAYER VI3 ;
  RECT 2516.740 5.940 2516.940 6.140 ;
  LAYER VI3 ;
  RECT 2516.340 6.340 2516.540 6.540 ;
  LAYER VI3 ;
  RECT 2516.340 5.940 2516.540 6.140 ;
  LAYER VI3 ;
  RECT 2515.940 6.340 2516.140 6.540 ;
  LAYER VI3 ;
  RECT 2515.940 5.940 2516.140 6.140 ;
  LAYER VI3 ;
  RECT 2535.780 5.880 2543.780 6.740 ;
  LAYER VI3 ;
  RECT 2543.380 6.340 2543.580 6.540 ;
  LAYER VI3 ;
  RECT 2543.380 5.940 2543.580 6.140 ;
  LAYER VI3 ;
  RECT 2542.980 6.340 2543.180 6.540 ;
  LAYER VI3 ;
  RECT 2542.980 5.940 2543.180 6.140 ;
  LAYER VI3 ;
  RECT 2542.580 6.340 2542.780 6.540 ;
  LAYER VI3 ;
  RECT 2542.580 5.940 2542.780 6.140 ;
  LAYER VI3 ;
  RECT 2542.180 6.340 2542.380 6.540 ;
  LAYER VI3 ;
  RECT 2542.180 5.940 2542.380 6.140 ;
  LAYER VI3 ;
  RECT 2541.780 6.340 2541.980 6.540 ;
  LAYER VI3 ;
  RECT 2541.780 5.940 2541.980 6.140 ;
  LAYER VI3 ;
  RECT 2541.380 6.340 2541.580 6.540 ;
  LAYER VI3 ;
  RECT 2541.380 5.940 2541.580 6.140 ;
  LAYER VI3 ;
  RECT 2540.980 6.340 2541.180 6.540 ;
  LAYER VI3 ;
  RECT 2540.980 5.940 2541.180 6.140 ;
  LAYER VI3 ;
  RECT 2540.580 6.340 2540.780 6.540 ;
  LAYER VI3 ;
  RECT 2540.580 5.940 2540.780 6.140 ;
  LAYER VI3 ;
  RECT 2540.180 6.340 2540.380 6.540 ;
  LAYER VI3 ;
  RECT 2540.180 5.940 2540.380 6.140 ;
  LAYER VI3 ;
  RECT 2539.780 6.340 2539.980 6.540 ;
  LAYER VI3 ;
  RECT 2539.780 5.940 2539.980 6.140 ;
  LAYER VI3 ;
  RECT 2539.380 6.340 2539.580 6.540 ;
  LAYER VI3 ;
  RECT 2539.380 5.940 2539.580 6.140 ;
  LAYER VI3 ;
  RECT 2538.980 6.340 2539.180 6.540 ;
  LAYER VI3 ;
  RECT 2538.980 5.940 2539.180 6.140 ;
  LAYER VI3 ;
  RECT 2538.580 6.340 2538.780 6.540 ;
  LAYER VI3 ;
  RECT 2538.580 5.940 2538.780 6.140 ;
  LAYER VI3 ;
  RECT 2538.180 6.340 2538.380 6.540 ;
  LAYER VI3 ;
  RECT 2538.180 5.940 2538.380 6.140 ;
  LAYER VI3 ;
  RECT 2537.780 6.340 2537.980 6.540 ;
  LAYER VI3 ;
  RECT 2537.780 5.940 2537.980 6.140 ;
  LAYER VI3 ;
  RECT 2537.380 6.340 2537.580 6.540 ;
  LAYER VI3 ;
  RECT 2537.380 5.940 2537.580 6.140 ;
  LAYER VI3 ;
  RECT 2536.980 6.340 2537.180 6.540 ;
  LAYER VI3 ;
  RECT 2536.980 5.940 2537.180 6.140 ;
  LAYER VI3 ;
  RECT 2536.580 6.340 2536.780 6.540 ;
  LAYER VI3 ;
  RECT 2536.580 5.940 2536.780 6.140 ;
  LAYER VI3 ;
  RECT 2536.180 6.340 2536.380 6.540 ;
  LAYER VI3 ;
  RECT 2536.180 5.940 2536.380 6.140 ;
  LAYER VI3 ;
  RECT 2535.780 6.340 2535.980 6.540 ;
  LAYER VI3 ;
  RECT 2535.780 5.940 2535.980 6.140 ;
  LAYER VI3 ;
  RECT 2556.860 5.880 2564.860 6.740 ;
  LAYER VI3 ;
  RECT 2564.460 6.340 2564.660 6.540 ;
  LAYER VI3 ;
  RECT 2564.460 5.940 2564.660 6.140 ;
  LAYER VI3 ;
  RECT 2564.060 6.340 2564.260 6.540 ;
  LAYER VI3 ;
  RECT 2564.060 5.940 2564.260 6.140 ;
  LAYER VI3 ;
  RECT 2563.660 6.340 2563.860 6.540 ;
  LAYER VI3 ;
  RECT 2563.660 5.940 2563.860 6.140 ;
  LAYER VI3 ;
  RECT 2563.260 6.340 2563.460 6.540 ;
  LAYER VI3 ;
  RECT 2563.260 5.940 2563.460 6.140 ;
  LAYER VI3 ;
  RECT 2562.860 6.340 2563.060 6.540 ;
  LAYER VI3 ;
  RECT 2562.860 5.940 2563.060 6.140 ;
  LAYER VI3 ;
  RECT 2562.460 6.340 2562.660 6.540 ;
  LAYER VI3 ;
  RECT 2562.460 5.940 2562.660 6.140 ;
  LAYER VI3 ;
  RECT 2562.060 6.340 2562.260 6.540 ;
  LAYER VI3 ;
  RECT 2562.060 5.940 2562.260 6.140 ;
  LAYER VI3 ;
  RECT 2561.660 6.340 2561.860 6.540 ;
  LAYER VI3 ;
  RECT 2561.660 5.940 2561.860 6.140 ;
  LAYER VI3 ;
  RECT 2561.260 6.340 2561.460 6.540 ;
  LAYER VI3 ;
  RECT 2561.260 5.940 2561.460 6.140 ;
  LAYER VI3 ;
  RECT 2560.860 6.340 2561.060 6.540 ;
  LAYER VI3 ;
  RECT 2560.860 5.940 2561.060 6.140 ;
  LAYER VI3 ;
  RECT 2560.460 6.340 2560.660 6.540 ;
  LAYER VI3 ;
  RECT 2560.460 5.940 2560.660 6.140 ;
  LAYER VI3 ;
  RECT 2560.060 6.340 2560.260 6.540 ;
  LAYER VI3 ;
  RECT 2560.060 5.940 2560.260 6.140 ;
  LAYER VI3 ;
  RECT 2559.660 6.340 2559.860 6.540 ;
  LAYER VI3 ;
  RECT 2559.660 5.940 2559.860 6.140 ;
  LAYER VI3 ;
  RECT 2559.260 6.340 2559.460 6.540 ;
  LAYER VI3 ;
  RECT 2559.260 5.940 2559.460 6.140 ;
  LAYER VI3 ;
  RECT 2558.860 6.340 2559.060 6.540 ;
  LAYER VI3 ;
  RECT 2558.860 5.940 2559.060 6.140 ;
  LAYER VI3 ;
  RECT 2558.460 6.340 2558.660 6.540 ;
  LAYER VI3 ;
  RECT 2558.460 5.940 2558.660 6.140 ;
  LAYER VI3 ;
  RECT 2558.060 6.340 2558.260 6.540 ;
  LAYER VI3 ;
  RECT 2558.060 5.940 2558.260 6.140 ;
  LAYER VI3 ;
  RECT 2557.660 6.340 2557.860 6.540 ;
  LAYER VI3 ;
  RECT 2557.660 5.940 2557.860 6.140 ;
  LAYER VI3 ;
  RECT 2557.260 6.340 2557.460 6.540 ;
  LAYER VI3 ;
  RECT 2557.260 5.940 2557.460 6.140 ;
  LAYER VI3 ;
  RECT 2556.860 6.340 2557.060 6.540 ;
  LAYER VI3 ;
  RECT 2556.860 5.940 2557.060 6.140 ;
  LAYER VI3 ;
  RECT 2576.700 5.880 2584.700 6.740 ;
  LAYER VI3 ;
  RECT 2584.300 6.340 2584.500 6.540 ;
  LAYER VI3 ;
  RECT 2584.300 5.940 2584.500 6.140 ;
  LAYER VI3 ;
  RECT 2583.900 6.340 2584.100 6.540 ;
  LAYER VI3 ;
  RECT 2583.900 5.940 2584.100 6.140 ;
  LAYER VI3 ;
  RECT 2583.500 6.340 2583.700 6.540 ;
  LAYER VI3 ;
  RECT 2583.500 5.940 2583.700 6.140 ;
  LAYER VI3 ;
  RECT 2583.100 6.340 2583.300 6.540 ;
  LAYER VI3 ;
  RECT 2583.100 5.940 2583.300 6.140 ;
  LAYER VI3 ;
  RECT 2582.700 6.340 2582.900 6.540 ;
  LAYER VI3 ;
  RECT 2582.700 5.940 2582.900 6.140 ;
  LAYER VI3 ;
  RECT 2582.300 6.340 2582.500 6.540 ;
  LAYER VI3 ;
  RECT 2582.300 5.940 2582.500 6.140 ;
  LAYER VI3 ;
  RECT 2581.900 6.340 2582.100 6.540 ;
  LAYER VI3 ;
  RECT 2581.900 5.940 2582.100 6.140 ;
  LAYER VI3 ;
  RECT 2581.500 6.340 2581.700 6.540 ;
  LAYER VI3 ;
  RECT 2581.500 5.940 2581.700 6.140 ;
  LAYER VI3 ;
  RECT 2581.100 6.340 2581.300 6.540 ;
  LAYER VI3 ;
  RECT 2581.100 5.940 2581.300 6.140 ;
  LAYER VI3 ;
  RECT 2580.700 6.340 2580.900 6.540 ;
  LAYER VI3 ;
  RECT 2580.700 5.940 2580.900 6.140 ;
  LAYER VI3 ;
  RECT 2580.300 6.340 2580.500 6.540 ;
  LAYER VI3 ;
  RECT 2580.300 5.940 2580.500 6.140 ;
  LAYER VI3 ;
  RECT 2579.900 6.340 2580.100 6.540 ;
  LAYER VI3 ;
  RECT 2579.900 5.940 2580.100 6.140 ;
  LAYER VI3 ;
  RECT 2579.500 6.340 2579.700 6.540 ;
  LAYER VI3 ;
  RECT 2579.500 5.940 2579.700 6.140 ;
  LAYER VI3 ;
  RECT 2579.100 6.340 2579.300 6.540 ;
  LAYER VI3 ;
  RECT 2579.100 5.940 2579.300 6.140 ;
  LAYER VI3 ;
  RECT 2578.700 6.340 2578.900 6.540 ;
  LAYER VI3 ;
  RECT 2578.700 5.940 2578.900 6.140 ;
  LAYER VI3 ;
  RECT 2578.300 6.340 2578.500 6.540 ;
  LAYER VI3 ;
  RECT 2578.300 5.940 2578.500 6.140 ;
  LAYER VI3 ;
  RECT 2577.900 6.340 2578.100 6.540 ;
  LAYER VI3 ;
  RECT 2577.900 5.940 2578.100 6.140 ;
  LAYER VI3 ;
  RECT 2577.500 6.340 2577.700 6.540 ;
  LAYER VI3 ;
  RECT 2577.500 5.940 2577.700 6.140 ;
  LAYER VI3 ;
  RECT 2577.100 6.340 2577.300 6.540 ;
  LAYER VI3 ;
  RECT 2577.100 5.940 2577.300 6.140 ;
  LAYER VI3 ;
  RECT 2576.700 6.340 2576.900 6.540 ;
  LAYER VI3 ;
  RECT 2576.700 5.940 2576.900 6.140 ;
  LAYER VI3 ;
  RECT 2597.780 5.880 2605.780 6.740 ;
  LAYER VI3 ;
  RECT 2605.380 6.340 2605.580 6.540 ;
  LAYER VI3 ;
  RECT 2605.380 5.940 2605.580 6.140 ;
  LAYER VI3 ;
  RECT 2604.980 6.340 2605.180 6.540 ;
  LAYER VI3 ;
  RECT 2604.980 5.940 2605.180 6.140 ;
  LAYER VI3 ;
  RECT 2604.580 6.340 2604.780 6.540 ;
  LAYER VI3 ;
  RECT 2604.580 5.940 2604.780 6.140 ;
  LAYER VI3 ;
  RECT 2604.180 6.340 2604.380 6.540 ;
  LAYER VI3 ;
  RECT 2604.180 5.940 2604.380 6.140 ;
  LAYER VI3 ;
  RECT 2603.780 6.340 2603.980 6.540 ;
  LAYER VI3 ;
  RECT 2603.780 5.940 2603.980 6.140 ;
  LAYER VI3 ;
  RECT 2603.380 6.340 2603.580 6.540 ;
  LAYER VI3 ;
  RECT 2603.380 5.940 2603.580 6.140 ;
  LAYER VI3 ;
  RECT 2602.980 6.340 2603.180 6.540 ;
  LAYER VI3 ;
  RECT 2602.980 5.940 2603.180 6.140 ;
  LAYER VI3 ;
  RECT 2602.580 6.340 2602.780 6.540 ;
  LAYER VI3 ;
  RECT 2602.580 5.940 2602.780 6.140 ;
  LAYER VI3 ;
  RECT 2602.180 6.340 2602.380 6.540 ;
  LAYER VI3 ;
  RECT 2602.180 5.940 2602.380 6.140 ;
  LAYER VI3 ;
  RECT 2601.780 6.340 2601.980 6.540 ;
  LAYER VI3 ;
  RECT 2601.780 5.940 2601.980 6.140 ;
  LAYER VI3 ;
  RECT 2601.380 6.340 2601.580 6.540 ;
  LAYER VI3 ;
  RECT 2601.380 5.940 2601.580 6.140 ;
  LAYER VI3 ;
  RECT 2600.980 6.340 2601.180 6.540 ;
  LAYER VI3 ;
  RECT 2600.980 5.940 2601.180 6.140 ;
  LAYER VI3 ;
  RECT 2600.580 6.340 2600.780 6.540 ;
  LAYER VI3 ;
  RECT 2600.580 5.940 2600.780 6.140 ;
  LAYER VI3 ;
  RECT 2600.180 6.340 2600.380 6.540 ;
  LAYER VI3 ;
  RECT 2600.180 5.940 2600.380 6.140 ;
  LAYER VI3 ;
  RECT 2599.780 6.340 2599.980 6.540 ;
  LAYER VI3 ;
  RECT 2599.780 5.940 2599.980 6.140 ;
  LAYER VI3 ;
  RECT 2599.380 6.340 2599.580 6.540 ;
  LAYER VI3 ;
  RECT 2599.380 5.940 2599.580 6.140 ;
  LAYER VI3 ;
  RECT 2598.980 6.340 2599.180 6.540 ;
  LAYER VI3 ;
  RECT 2598.980 5.940 2599.180 6.140 ;
  LAYER VI3 ;
  RECT 2598.580 6.340 2598.780 6.540 ;
  LAYER VI3 ;
  RECT 2598.580 5.940 2598.780 6.140 ;
  LAYER VI3 ;
  RECT 2598.180 6.340 2598.380 6.540 ;
  LAYER VI3 ;
  RECT 2598.180 5.940 2598.380 6.140 ;
  LAYER VI3 ;
  RECT 2597.780 6.340 2597.980 6.540 ;
  LAYER VI3 ;
  RECT 2597.780 5.940 2597.980 6.140 ;
  LAYER VI3 ;
  RECT 2617.620 5.880 2625.620 6.740 ;
  LAYER VI3 ;
  RECT 2625.220 6.340 2625.420 6.540 ;
  LAYER VI3 ;
  RECT 2625.220 5.940 2625.420 6.140 ;
  LAYER VI3 ;
  RECT 2624.820 6.340 2625.020 6.540 ;
  LAYER VI3 ;
  RECT 2624.820 5.940 2625.020 6.140 ;
  LAYER VI3 ;
  RECT 2624.420 6.340 2624.620 6.540 ;
  LAYER VI3 ;
  RECT 2624.420 5.940 2624.620 6.140 ;
  LAYER VI3 ;
  RECT 2624.020 6.340 2624.220 6.540 ;
  LAYER VI3 ;
  RECT 2624.020 5.940 2624.220 6.140 ;
  LAYER VI3 ;
  RECT 2623.620 6.340 2623.820 6.540 ;
  LAYER VI3 ;
  RECT 2623.620 5.940 2623.820 6.140 ;
  LAYER VI3 ;
  RECT 2623.220 6.340 2623.420 6.540 ;
  LAYER VI3 ;
  RECT 2623.220 5.940 2623.420 6.140 ;
  LAYER VI3 ;
  RECT 2622.820 6.340 2623.020 6.540 ;
  LAYER VI3 ;
  RECT 2622.820 5.940 2623.020 6.140 ;
  LAYER VI3 ;
  RECT 2622.420 6.340 2622.620 6.540 ;
  LAYER VI3 ;
  RECT 2622.420 5.940 2622.620 6.140 ;
  LAYER VI3 ;
  RECT 2622.020 6.340 2622.220 6.540 ;
  LAYER VI3 ;
  RECT 2622.020 5.940 2622.220 6.140 ;
  LAYER VI3 ;
  RECT 2621.620 6.340 2621.820 6.540 ;
  LAYER VI3 ;
  RECT 2621.620 5.940 2621.820 6.140 ;
  LAYER VI3 ;
  RECT 2621.220 6.340 2621.420 6.540 ;
  LAYER VI3 ;
  RECT 2621.220 5.940 2621.420 6.140 ;
  LAYER VI3 ;
  RECT 2620.820 6.340 2621.020 6.540 ;
  LAYER VI3 ;
  RECT 2620.820 5.940 2621.020 6.140 ;
  LAYER VI3 ;
  RECT 2620.420 6.340 2620.620 6.540 ;
  LAYER VI3 ;
  RECT 2620.420 5.940 2620.620 6.140 ;
  LAYER VI3 ;
  RECT 2620.020 6.340 2620.220 6.540 ;
  LAYER VI3 ;
  RECT 2620.020 5.940 2620.220 6.140 ;
  LAYER VI3 ;
  RECT 2619.620 6.340 2619.820 6.540 ;
  LAYER VI3 ;
  RECT 2619.620 5.940 2619.820 6.140 ;
  LAYER VI3 ;
  RECT 2619.220 6.340 2619.420 6.540 ;
  LAYER VI3 ;
  RECT 2619.220 5.940 2619.420 6.140 ;
  LAYER VI3 ;
  RECT 2618.820 6.340 2619.020 6.540 ;
  LAYER VI3 ;
  RECT 2618.820 5.940 2619.020 6.140 ;
  LAYER VI3 ;
  RECT 2618.420 6.340 2618.620 6.540 ;
  LAYER VI3 ;
  RECT 2618.420 5.940 2618.620 6.140 ;
  LAYER VI3 ;
  RECT 2618.020 6.340 2618.220 6.540 ;
  LAYER VI3 ;
  RECT 2618.020 5.940 2618.220 6.140 ;
  LAYER VI3 ;
  RECT 2617.620 6.340 2617.820 6.540 ;
  LAYER VI3 ;
  RECT 2617.620 5.940 2617.820 6.140 ;
  LAYER VI3 ;
  RECT 2638.700 5.880 2646.700 6.740 ;
  LAYER VI3 ;
  RECT 2646.300 6.340 2646.500 6.540 ;
  LAYER VI3 ;
  RECT 2646.300 5.940 2646.500 6.140 ;
  LAYER VI3 ;
  RECT 2645.900 6.340 2646.100 6.540 ;
  LAYER VI3 ;
  RECT 2645.900 5.940 2646.100 6.140 ;
  LAYER VI3 ;
  RECT 2645.500 6.340 2645.700 6.540 ;
  LAYER VI3 ;
  RECT 2645.500 5.940 2645.700 6.140 ;
  LAYER VI3 ;
  RECT 2645.100 6.340 2645.300 6.540 ;
  LAYER VI3 ;
  RECT 2645.100 5.940 2645.300 6.140 ;
  LAYER VI3 ;
  RECT 2644.700 6.340 2644.900 6.540 ;
  LAYER VI3 ;
  RECT 2644.700 5.940 2644.900 6.140 ;
  LAYER VI3 ;
  RECT 2644.300 6.340 2644.500 6.540 ;
  LAYER VI3 ;
  RECT 2644.300 5.940 2644.500 6.140 ;
  LAYER VI3 ;
  RECT 2643.900 6.340 2644.100 6.540 ;
  LAYER VI3 ;
  RECT 2643.900 5.940 2644.100 6.140 ;
  LAYER VI3 ;
  RECT 2643.500 6.340 2643.700 6.540 ;
  LAYER VI3 ;
  RECT 2643.500 5.940 2643.700 6.140 ;
  LAYER VI3 ;
  RECT 2643.100 6.340 2643.300 6.540 ;
  LAYER VI3 ;
  RECT 2643.100 5.940 2643.300 6.140 ;
  LAYER VI3 ;
  RECT 2642.700 6.340 2642.900 6.540 ;
  LAYER VI3 ;
  RECT 2642.700 5.940 2642.900 6.140 ;
  LAYER VI3 ;
  RECT 2642.300 6.340 2642.500 6.540 ;
  LAYER VI3 ;
  RECT 2642.300 5.940 2642.500 6.140 ;
  LAYER VI3 ;
  RECT 2641.900 6.340 2642.100 6.540 ;
  LAYER VI3 ;
  RECT 2641.900 5.940 2642.100 6.140 ;
  LAYER VI3 ;
  RECT 2641.500 6.340 2641.700 6.540 ;
  LAYER VI3 ;
  RECT 2641.500 5.940 2641.700 6.140 ;
  LAYER VI3 ;
  RECT 2641.100 6.340 2641.300 6.540 ;
  LAYER VI3 ;
  RECT 2641.100 5.940 2641.300 6.140 ;
  LAYER VI3 ;
  RECT 2640.700 6.340 2640.900 6.540 ;
  LAYER VI3 ;
  RECT 2640.700 5.940 2640.900 6.140 ;
  LAYER VI3 ;
  RECT 2640.300 6.340 2640.500 6.540 ;
  LAYER VI3 ;
  RECT 2640.300 5.940 2640.500 6.140 ;
  LAYER VI3 ;
  RECT 2639.900 6.340 2640.100 6.540 ;
  LAYER VI3 ;
  RECT 2639.900 5.940 2640.100 6.140 ;
  LAYER VI3 ;
  RECT 2639.500 6.340 2639.700 6.540 ;
  LAYER VI3 ;
  RECT 2639.500 5.940 2639.700 6.140 ;
  LAYER VI3 ;
  RECT 2639.100 6.340 2639.300 6.540 ;
  LAYER VI3 ;
  RECT 2639.100 5.940 2639.300 6.140 ;
  LAYER VI3 ;
  RECT 2638.700 6.340 2638.900 6.540 ;
  LAYER VI3 ;
  RECT 2638.700 5.940 2638.900 6.140 ;
  LAYER VI3 ;
  RECT 2658.540 5.880 2666.540 6.740 ;
  LAYER VI3 ;
  RECT 2666.140 6.340 2666.340 6.540 ;
  LAYER VI3 ;
  RECT 2666.140 5.940 2666.340 6.140 ;
  LAYER VI3 ;
  RECT 2665.740 6.340 2665.940 6.540 ;
  LAYER VI3 ;
  RECT 2665.740 5.940 2665.940 6.140 ;
  LAYER VI3 ;
  RECT 2665.340 6.340 2665.540 6.540 ;
  LAYER VI3 ;
  RECT 2665.340 5.940 2665.540 6.140 ;
  LAYER VI3 ;
  RECT 2664.940 6.340 2665.140 6.540 ;
  LAYER VI3 ;
  RECT 2664.940 5.940 2665.140 6.140 ;
  LAYER VI3 ;
  RECT 2664.540 6.340 2664.740 6.540 ;
  LAYER VI3 ;
  RECT 2664.540 5.940 2664.740 6.140 ;
  LAYER VI3 ;
  RECT 2664.140 6.340 2664.340 6.540 ;
  LAYER VI3 ;
  RECT 2664.140 5.940 2664.340 6.140 ;
  LAYER VI3 ;
  RECT 2663.740 6.340 2663.940 6.540 ;
  LAYER VI3 ;
  RECT 2663.740 5.940 2663.940 6.140 ;
  LAYER VI3 ;
  RECT 2663.340 6.340 2663.540 6.540 ;
  LAYER VI3 ;
  RECT 2663.340 5.940 2663.540 6.140 ;
  LAYER VI3 ;
  RECT 2662.940 6.340 2663.140 6.540 ;
  LAYER VI3 ;
  RECT 2662.940 5.940 2663.140 6.140 ;
  LAYER VI3 ;
  RECT 2662.540 6.340 2662.740 6.540 ;
  LAYER VI3 ;
  RECT 2662.540 5.940 2662.740 6.140 ;
  LAYER VI3 ;
  RECT 2662.140 6.340 2662.340 6.540 ;
  LAYER VI3 ;
  RECT 2662.140 5.940 2662.340 6.140 ;
  LAYER VI3 ;
  RECT 2661.740 6.340 2661.940 6.540 ;
  LAYER VI3 ;
  RECT 2661.740 5.940 2661.940 6.140 ;
  LAYER VI3 ;
  RECT 2661.340 6.340 2661.540 6.540 ;
  LAYER VI3 ;
  RECT 2661.340 5.940 2661.540 6.140 ;
  LAYER VI3 ;
  RECT 2660.940 6.340 2661.140 6.540 ;
  LAYER VI3 ;
  RECT 2660.940 5.940 2661.140 6.140 ;
  LAYER VI3 ;
  RECT 2660.540 6.340 2660.740 6.540 ;
  LAYER VI3 ;
  RECT 2660.540 5.940 2660.740 6.140 ;
  LAYER VI3 ;
  RECT 2660.140 6.340 2660.340 6.540 ;
  LAYER VI3 ;
  RECT 2660.140 5.940 2660.340 6.140 ;
  LAYER VI3 ;
  RECT 2659.740 6.340 2659.940 6.540 ;
  LAYER VI3 ;
  RECT 2659.740 5.940 2659.940 6.140 ;
  LAYER VI3 ;
  RECT 2659.340 6.340 2659.540 6.540 ;
  LAYER VI3 ;
  RECT 2659.340 5.940 2659.540 6.140 ;
  LAYER VI3 ;
  RECT 2658.940 6.340 2659.140 6.540 ;
  LAYER VI3 ;
  RECT 2658.940 5.940 2659.140 6.140 ;
  LAYER VI3 ;
  RECT 2658.540 6.340 2658.740 6.540 ;
  LAYER VI3 ;
  RECT 2658.540 5.940 2658.740 6.140 ;
  LAYER VI3 ;
  RECT 1335.440 5.880 1338.890 6.740 ;
  LAYER VI3 ;
  RECT 1338.640 6.340 1338.840 6.540 ;
  LAYER VI3 ;
  RECT 1338.640 5.940 1338.840 6.140 ;
  LAYER VI3 ;
  RECT 1338.240 6.340 1338.440 6.540 ;
  LAYER VI3 ;
  RECT 1338.240 5.940 1338.440 6.140 ;
  LAYER VI3 ;
  RECT 1337.840 6.340 1338.040 6.540 ;
  LAYER VI3 ;
  RECT 1337.840 5.940 1338.040 6.140 ;
  LAYER VI3 ;
  RECT 1337.440 6.340 1337.640 6.540 ;
  LAYER VI3 ;
  RECT 1337.440 5.940 1337.640 6.140 ;
  LAYER VI3 ;
  RECT 1337.040 6.340 1337.240 6.540 ;
  LAYER VI3 ;
  RECT 1337.040 5.940 1337.240 6.140 ;
  LAYER VI3 ;
  RECT 1336.640 6.340 1336.840 6.540 ;
  LAYER VI3 ;
  RECT 1336.640 5.940 1336.840 6.140 ;
  LAYER VI3 ;
  RECT 1336.240 6.340 1336.440 6.540 ;
  LAYER VI3 ;
  RECT 1336.240 5.940 1336.440 6.140 ;
  LAYER VI3 ;
  RECT 1335.840 6.340 1336.040 6.540 ;
  LAYER VI3 ;
  RECT 1335.840 5.940 1336.040 6.140 ;
  LAYER VI3 ;
  RECT 1335.440 6.340 1335.640 6.540 ;
  LAYER VI3 ;
  RECT 1335.440 5.940 1335.640 6.140 ;
  LAYER VI3 ;
  RECT 1344.290 5.880 1350.210 6.740 ;
  LAYER VI3 ;
  RECT 1349.890 6.340 1350.090 6.540 ;
  LAYER VI3 ;
  RECT 1349.890 5.940 1350.090 6.140 ;
  LAYER VI3 ;
  RECT 1349.490 6.340 1349.690 6.540 ;
  LAYER VI3 ;
  RECT 1349.490 5.940 1349.690 6.140 ;
  LAYER VI3 ;
  RECT 1349.090 6.340 1349.290 6.540 ;
  LAYER VI3 ;
  RECT 1349.090 5.940 1349.290 6.140 ;
  LAYER VI3 ;
  RECT 1348.690 6.340 1348.890 6.540 ;
  LAYER VI3 ;
  RECT 1348.690 5.940 1348.890 6.140 ;
  LAYER VI3 ;
  RECT 1348.290 6.340 1348.490 6.540 ;
  LAYER VI3 ;
  RECT 1348.290 5.940 1348.490 6.140 ;
  LAYER VI3 ;
  RECT 1347.890 6.340 1348.090 6.540 ;
  LAYER VI3 ;
  RECT 1347.890 5.940 1348.090 6.140 ;
  LAYER VI3 ;
  RECT 1347.490 6.340 1347.690 6.540 ;
  LAYER VI3 ;
  RECT 1347.490 5.940 1347.690 6.140 ;
  LAYER VI3 ;
  RECT 1347.090 6.340 1347.290 6.540 ;
  LAYER VI3 ;
  RECT 1347.090 5.940 1347.290 6.140 ;
  LAYER VI3 ;
  RECT 1346.690 6.340 1346.890 6.540 ;
  LAYER VI3 ;
  RECT 1346.690 5.940 1346.890 6.140 ;
  LAYER VI3 ;
  RECT 1346.290 6.340 1346.490 6.540 ;
  LAYER VI3 ;
  RECT 1346.290 5.940 1346.490 6.140 ;
  LAYER VI3 ;
  RECT 1345.890 6.340 1346.090 6.540 ;
  LAYER VI3 ;
  RECT 1345.890 5.940 1346.090 6.140 ;
  LAYER VI3 ;
  RECT 1345.490 6.340 1345.690 6.540 ;
  LAYER VI3 ;
  RECT 1345.490 5.940 1345.690 6.140 ;
  LAYER VI3 ;
  RECT 1345.090 6.340 1345.290 6.540 ;
  LAYER VI3 ;
  RECT 1345.090 5.940 1345.290 6.140 ;
  LAYER VI3 ;
  RECT 1344.690 6.340 1344.890 6.540 ;
  LAYER VI3 ;
  RECT 1344.690 5.940 1344.890 6.140 ;
  LAYER VI3 ;
  RECT 1344.290 6.340 1344.490 6.540 ;
  LAYER VI3 ;
  RECT 1344.290 5.940 1344.490 6.140 ;
  LAYER VI3 ;
  RECT 1327.160 5.880 1328.920 6.740 ;
  LAYER VI3 ;
  RECT 1328.360 6.340 1328.560 6.540 ;
  LAYER VI3 ;
  RECT 1328.360 5.940 1328.560 6.140 ;
  LAYER VI3 ;
  RECT 1327.960 6.340 1328.160 6.540 ;
  LAYER VI3 ;
  RECT 1327.960 5.940 1328.160 6.140 ;
  LAYER VI3 ;
  RECT 1327.560 6.340 1327.760 6.540 ;
  LAYER VI3 ;
  RECT 1327.560 5.940 1327.760 6.140 ;
  LAYER VI3 ;
  RECT 1327.160 6.340 1327.360 6.540 ;
  LAYER VI3 ;
  RECT 1327.160 5.940 1327.360 6.140 ;
  LAYER VI3 ;
  RECT 1321.820 5.880 1323.580 6.740 ;
  LAYER VI3 ;
  RECT 1323.020 6.340 1323.220 6.540 ;
  LAYER VI3 ;
  RECT 1323.020 5.940 1323.220 6.140 ;
  LAYER VI3 ;
  RECT 1322.620 6.340 1322.820 6.540 ;
  LAYER VI3 ;
  RECT 1322.620 5.940 1322.820 6.140 ;
  LAYER VI3 ;
  RECT 1322.220 6.340 1322.420 6.540 ;
  LAYER VI3 ;
  RECT 1322.220 5.940 1322.420 6.140 ;
  LAYER VI3 ;
  RECT 1321.820 6.340 1322.020 6.540 ;
  LAYER VI3 ;
  RECT 1321.820 5.940 1322.020 6.140 ;
  LAYER VI3 ;
  RECT 1317.820 5.880 1319.580 6.740 ;
  LAYER VI3 ;
  RECT 1319.020 6.340 1319.220 6.540 ;
  LAYER VI3 ;
  RECT 1319.020 5.940 1319.220 6.140 ;
  LAYER VI3 ;
  RECT 1318.620 6.340 1318.820 6.540 ;
  LAYER VI3 ;
  RECT 1318.620 5.940 1318.820 6.140 ;
  LAYER VI3 ;
  RECT 1318.220 6.340 1318.420 6.540 ;
  LAYER VI3 ;
  RECT 1318.220 5.940 1318.420 6.140 ;
  LAYER VI3 ;
  RECT 1317.820 6.340 1318.020 6.540 ;
  LAYER VI3 ;
  RECT 1317.820 5.940 1318.020 6.140 ;
  LAYER VI3 ;
  RECT 4.280 57.100 5.140 61.420 ;
  LAYER VI3 ;
  RECT 4.740 61.100 4.940 61.300 ;
  LAYER VI3 ;
  RECT 4.740 60.700 4.940 60.900 ;
  LAYER VI3 ;
  RECT 4.740 60.300 4.940 60.500 ;
  LAYER VI3 ;
  RECT 4.740 59.900 4.940 60.100 ;
  LAYER VI3 ;
  RECT 4.740 59.500 4.940 59.700 ;
  LAYER VI3 ;
  RECT 4.740 59.100 4.940 59.300 ;
  LAYER VI3 ;
  RECT 4.740 58.700 4.940 58.900 ;
  LAYER VI3 ;
  RECT 4.740 58.300 4.940 58.500 ;
  LAYER VI3 ;
  RECT 4.740 57.900 4.940 58.100 ;
  LAYER VI3 ;
  RECT 4.740 57.500 4.940 57.700 ;
  LAYER VI3 ;
  RECT 4.740 57.100 4.940 57.300 ;
  LAYER VI3 ;
  RECT 4.340 61.100 4.540 61.300 ;
  LAYER VI3 ;
  RECT 4.340 60.700 4.540 60.900 ;
  LAYER VI3 ;
  RECT 4.340 60.300 4.540 60.500 ;
  LAYER VI3 ;
  RECT 4.340 59.900 4.540 60.100 ;
  LAYER VI3 ;
  RECT 4.340 59.500 4.540 59.700 ;
  LAYER VI3 ;
  RECT 4.340 59.100 4.540 59.300 ;
  LAYER VI3 ;
  RECT 4.340 58.700 4.540 58.900 ;
  LAYER VI3 ;
  RECT 4.340 58.300 4.540 58.500 ;
  LAYER VI3 ;
  RECT 4.340 57.900 4.540 58.100 ;
  LAYER VI3 ;
  RECT 4.340 57.500 4.540 57.700 ;
  LAYER VI3 ;
  RECT 4.340 57.100 4.540 57.300 ;
  LAYER VI2 ;
  RECT 4.280 57.100 5.140 61.420 ;
  LAYER VI2 ;
  RECT 4.740 61.100 4.940 61.300 ;
  LAYER VI2 ;
  RECT 4.740 60.700 4.940 60.900 ;
  LAYER VI2 ;
  RECT 4.740 60.300 4.940 60.500 ;
  LAYER VI2 ;
  RECT 4.740 59.900 4.940 60.100 ;
  LAYER VI2 ;
  RECT 4.740 59.500 4.940 59.700 ;
  LAYER VI2 ;
  RECT 4.740 59.100 4.940 59.300 ;
  LAYER VI2 ;
  RECT 4.740 58.700 4.940 58.900 ;
  LAYER VI2 ;
  RECT 4.740 58.300 4.940 58.500 ;
  LAYER VI2 ;
  RECT 4.740 57.900 4.940 58.100 ;
  LAYER VI2 ;
  RECT 4.740 57.500 4.940 57.700 ;
  LAYER VI2 ;
  RECT 4.740 57.100 4.940 57.300 ;
  LAYER VI2 ;
  RECT 4.340 61.100 4.540 61.300 ;
  LAYER VI2 ;
  RECT 4.340 60.700 4.540 60.900 ;
  LAYER VI2 ;
  RECT 4.340 60.300 4.540 60.500 ;
  LAYER VI2 ;
  RECT 4.340 59.900 4.540 60.100 ;
  LAYER VI2 ;
  RECT 4.340 59.500 4.540 59.700 ;
  LAYER VI2 ;
  RECT 4.340 59.100 4.540 59.300 ;
  LAYER VI2 ;
  RECT 4.340 58.700 4.540 58.900 ;
  LAYER VI2 ;
  RECT 4.340 58.300 4.540 58.500 ;
  LAYER VI2 ;
  RECT 4.340 57.900 4.540 58.100 ;
  LAYER VI2 ;
  RECT 4.340 57.500 4.540 57.700 ;
  LAYER VI2 ;
  RECT 4.340 57.100 4.540 57.300 ;
  LAYER VI3 ;
  RECT 4.280 45.560 5.140 46.160 ;
  LAYER VI3 ;
  RECT 4.680 45.620 4.880 45.820 ;
  LAYER VI3 ;
  RECT 4.280 45.620 4.480 45.820 ;
  LAYER VI2 ;
  RECT 4.280 45.560 5.140 46.160 ;
  LAYER VI2 ;
  RECT 4.680 45.620 4.880 45.820 ;
  LAYER VI2 ;
  RECT 4.280 45.620 4.480 45.820 ;
  LAYER VI3 ;
  RECT 4.280 39.480 5.140 40.080 ;
  LAYER VI3 ;
  RECT 4.680 39.540 4.880 39.740 ;
  LAYER VI3 ;
  RECT 4.280 39.540 4.480 39.740 ;
  LAYER VI2 ;
  RECT 4.280 39.480 5.140 40.080 ;
  LAYER VI2 ;
  RECT 4.680 39.540 4.880 39.740 ;
  LAYER VI2 ;
  RECT 4.280 39.540 4.480 39.740 ;
  LAYER VI3 ;
  RECT 4.280 36.320 5.140 37.320 ;
  LAYER VI3 ;
  RECT 4.740 36.720 4.940 36.920 ;
  LAYER VI3 ;
  RECT 4.740 36.320 4.940 36.520 ;
  LAYER VI3 ;
  RECT 4.340 36.720 4.540 36.920 ;
  LAYER VI3 ;
  RECT 4.340 36.320 4.540 36.520 ;
  LAYER VI2 ;
  RECT 4.280 36.320 5.140 37.320 ;
  LAYER VI2 ;
  RECT 4.740 36.720 4.940 36.920 ;
  LAYER VI2 ;
  RECT 4.740 36.320 4.940 36.520 ;
  LAYER VI2 ;
  RECT 4.340 36.720 4.540 36.920 ;
  LAYER VI2 ;
  RECT 4.340 36.320 4.540 36.520 ;
  LAYER VI3 ;
  RECT 4.280 24.170 5.140 25.170 ;
  LAYER VI3 ;
  RECT 4.740 24.570 4.940 24.770 ;
  LAYER VI3 ;
  RECT 4.740 24.170 4.940 24.370 ;
  LAYER VI3 ;
  RECT 4.340 24.570 4.540 24.770 ;
  LAYER VI3 ;
  RECT 4.340 24.170 4.540 24.370 ;
  LAYER VI2 ;
  RECT 4.280 24.170 5.140 25.170 ;
  LAYER VI2 ;
  RECT 4.740 24.570 4.940 24.770 ;
  LAYER VI2 ;
  RECT 4.740 24.170 4.940 24.370 ;
  LAYER VI2 ;
  RECT 4.340 24.570 4.540 24.770 ;
  LAYER VI2 ;
  RECT 4.340 24.170 4.540 24.370 ;
  LAYER VI3 ;
  RECT 4.280 21.230 5.140 22.070 ;
  LAYER VI3 ;
  RECT 4.680 21.690 4.880 21.890 ;
  LAYER VI3 ;
  RECT 4.680 21.290 4.880 21.490 ;
  LAYER VI3 ;
  RECT 4.280 21.690 4.480 21.890 ;
  LAYER VI3 ;
  RECT 4.280 21.290 4.480 21.490 ;
  LAYER VI2 ;
  RECT 4.280 21.230 5.140 22.070 ;
  LAYER VI2 ;
  RECT 4.680 21.690 4.880 21.890 ;
  LAYER VI2 ;
  RECT 4.680 21.290 4.880 21.490 ;
  LAYER VI2 ;
  RECT 4.280 21.690 4.480 21.890 ;
  LAYER VI2 ;
  RECT 4.280 21.290 4.480 21.490 ;
  LAYER VI3 ;
  RECT 4.280 18.730 5.140 19.730 ;
  LAYER VI3 ;
  RECT 4.740 19.130 4.940 19.330 ;
  LAYER VI3 ;
  RECT 4.740 18.730 4.940 18.930 ;
  LAYER VI3 ;
  RECT 4.340 19.130 4.540 19.330 ;
  LAYER VI3 ;
  RECT 4.340 18.730 4.540 18.930 ;
  LAYER VI2 ;
  RECT 4.280 18.730 5.140 19.730 ;
  LAYER VI2 ;
  RECT 4.740 19.130 4.940 19.330 ;
  LAYER VI2 ;
  RECT 4.740 18.730 4.940 18.930 ;
  LAYER VI2 ;
  RECT 4.340 19.130 4.540 19.330 ;
  LAYER VI2 ;
  RECT 4.340 18.730 4.540 18.930 ;
  LAYER VI3 ;
  RECT 4.280 14.200 5.140 15.200 ;
  LAYER VI3 ;
  RECT 4.740 14.600 4.940 14.800 ;
  LAYER VI3 ;
  RECT 4.740 14.200 4.940 14.400 ;
  LAYER VI3 ;
  RECT 4.340 14.600 4.540 14.800 ;
  LAYER VI3 ;
  RECT 4.340 14.200 4.540 14.400 ;
  LAYER VI2 ;
  RECT 4.280 14.200 5.140 15.200 ;
  LAYER VI2 ;
  RECT 4.740 14.600 4.940 14.800 ;
  LAYER VI2 ;
  RECT 4.740 14.200 4.940 14.400 ;
  LAYER VI2 ;
  RECT 4.340 14.600 4.540 14.800 ;
  LAYER VI2 ;
  RECT 4.340 14.200 4.540 14.400 ;
  LAYER VI3 ;
  RECT 4.280 9.570 5.140 11.170 ;
  LAYER VI3 ;
  RECT 4.740 10.770 4.940 10.970 ;
  LAYER VI3 ;
  RECT 4.740 10.370 4.940 10.570 ;
  LAYER VI3 ;
  RECT 4.740 9.970 4.940 10.170 ;
  LAYER VI3 ;
  RECT 4.740 9.570 4.940 9.770 ;
  LAYER VI3 ;
  RECT 4.340 10.770 4.540 10.970 ;
  LAYER VI3 ;
  RECT 4.340 10.370 4.540 10.570 ;
  LAYER VI3 ;
  RECT 4.340 9.970 4.540 10.170 ;
  LAYER VI3 ;
  RECT 4.340 9.570 4.540 9.770 ;
  LAYER VI2 ;
  RECT 4.280 9.570 5.140 11.170 ;
  LAYER VI2 ;
  RECT 4.740 10.770 4.940 10.970 ;
  LAYER VI2 ;
  RECT 4.740 10.370 4.940 10.570 ;
  LAYER VI2 ;
  RECT 4.740 9.970 4.940 10.170 ;
  LAYER VI2 ;
  RECT 4.740 9.570 4.940 9.770 ;
  LAYER VI2 ;
  RECT 4.340 10.770 4.540 10.970 ;
  LAYER VI2 ;
  RECT 4.340 10.370 4.540 10.570 ;
  LAYER VI2 ;
  RECT 4.340 9.970 4.540 10.170 ;
  LAYER VI2 ;
  RECT 4.340 9.570 4.540 9.770 ;
  LAYER VI3 ;
  RECT 5.420 5.880 6.560 6.740 ;
  LAYER VI3 ;
  RECT 6.220 6.340 6.420 6.540 ;
  LAYER VI3 ;
  RECT 6.220 5.940 6.420 6.140 ;
  LAYER VI3 ;
  RECT 5.820 6.340 6.020 6.540 ;
  LAYER VI3 ;
  RECT 5.820 5.940 6.020 6.140 ;
  LAYER VI3 ;
  RECT 5.420 6.340 5.620 6.540 ;
  LAYER VI3 ;
  RECT 5.420 5.940 5.620 6.140 ;
  LAYER VI3 ;
  RECT 8.360 5.880 16.360 6.740 ;
  LAYER VI3 ;
  RECT 15.960 6.340 16.160 6.540 ;
  LAYER VI3 ;
  RECT 15.960 5.940 16.160 6.140 ;
  LAYER VI3 ;
  RECT 15.560 6.340 15.760 6.540 ;
  LAYER VI3 ;
  RECT 15.560 5.940 15.760 6.140 ;
  LAYER VI3 ;
  RECT 15.160 6.340 15.360 6.540 ;
  LAYER VI3 ;
  RECT 15.160 5.940 15.360 6.140 ;
  LAYER VI3 ;
  RECT 14.760 6.340 14.960 6.540 ;
  LAYER VI3 ;
  RECT 14.760 5.940 14.960 6.140 ;
  LAYER VI3 ;
  RECT 14.360 6.340 14.560 6.540 ;
  LAYER VI3 ;
  RECT 14.360 5.940 14.560 6.140 ;
  LAYER VI3 ;
  RECT 13.960 6.340 14.160 6.540 ;
  LAYER VI3 ;
  RECT 13.960 5.940 14.160 6.140 ;
  LAYER VI3 ;
  RECT 13.560 6.340 13.760 6.540 ;
  LAYER VI3 ;
  RECT 13.560 5.940 13.760 6.140 ;
  LAYER VI3 ;
  RECT 13.160 6.340 13.360 6.540 ;
  LAYER VI3 ;
  RECT 13.160 5.940 13.360 6.140 ;
  LAYER VI3 ;
  RECT 12.760 6.340 12.960 6.540 ;
  LAYER VI3 ;
  RECT 12.760 5.940 12.960 6.140 ;
  LAYER VI3 ;
  RECT 12.360 6.340 12.560 6.540 ;
  LAYER VI3 ;
  RECT 12.360 5.940 12.560 6.140 ;
  LAYER VI3 ;
  RECT 11.960 6.340 12.160 6.540 ;
  LAYER VI3 ;
  RECT 11.960 5.940 12.160 6.140 ;
  LAYER VI3 ;
  RECT 11.560 6.340 11.760 6.540 ;
  LAYER VI3 ;
  RECT 11.560 5.940 11.760 6.140 ;
  LAYER VI3 ;
  RECT 11.160 6.340 11.360 6.540 ;
  LAYER VI3 ;
  RECT 11.160 5.940 11.360 6.140 ;
  LAYER VI3 ;
  RECT 10.760 6.340 10.960 6.540 ;
  LAYER VI3 ;
  RECT 10.760 5.940 10.960 6.140 ;
  LAYER VI3 ;
  RECT 10.360 6.340 10.560 6.540 ;
  LAYER VI3 ;
  RECT 10.360 5.940 10.560 6.140 ;
  LAYER VI3 ;
  RECT 9.960 6.340 10.160 6.540 ;
  LAYER VI3 ;
  RECT 9.960 5.940 10.160 6.140 ;
  LAYER VI3 ;
  RECT 9.560 6.340 9.760 6.540 ;
  LAYER VI3 ;
  RECT 9.560 5.940 9.760 6.140 ;
  LAYER VI3 ;
  RECT 9.160 6.340 9.360 6.540 ;
  LAYER VI3 ;
  RECT 9.160 5.940 9.360 6.140 ;
  LAYER VI3 ;
  RECT 8.760 6.340 8.960 6.540 ;
  LAYER VI3 ;
  RECT 8.760 5.940 8.960 6.140 ;
  LAYER VI3 ;
  RECT 8.360 6.340 8.560 6.540 ;
  LAYER VI3 ;
  RECT 8.360 5.940 8.560 6.140 ;
  LAYER VI3 ;
  RECT 28.200 5.880 36.200 6.740 ;
  LAYER VI3 ;
  RECT 35.800 6.340 36.000 6.540 ;
  LAYER VI3 ;
  RECT 35.800 5.940 36.000 6.140 ;
  LAYER VI3 ;
  RECT 35.400 6.340 35.600 6.540 ;
  LAYER VI3 ;
  RECT 35.400 5.940 35.600 6.140 ;
  LAYER VI3 ;
  RECT 35.000 6.340 35.200 6.540 ;
  LAYER VI3 ;
  RECT 35.000 5.940 35.200 6.140 ;
  LAYER VI3 ;
  RECT 34.600 6.340 34.800 6.540 ;
  LAYER VI3 ;
  RECT 34.600 5.940 34.800 6.140 ;
  LAYER VI3 ;
  RECT 34.200 6.340 34.400 6.540 ;
  LAYER VI3 ;
  RECT 34.200 5.940 34.400 6.140 ;
  LAYER VI3 ;
  RECT 33.800 6.340 34.000 6.540 ;
  LAYER VI3 ;
  RECT 33.800 5.940 34.000 6.140 ;
  LAYER VI3 ;
  RECT 33.400 6.340 33.600 6.540 ;
  LAYER VI3 ;
  RECT 33.400 5.940 33.600 6.140 ;
  LAYER VI3 ;
  RECT 33.000 6.340 33.200 6.540 ;
  LAYER VI3 ;
  RECT 33.000 5.940 33.200 6.140 ;
  LAYER VI3 ;
  RECT 32.600 6.340 32.800 6.540 ;
  LAYER VI3 ;
  RECT 32.600 5.940 32.800 6.140 ;
  LAYER VI3 ;
  RECT 32.200 6.340 32.400 6.540 ;
  LAYER VI3 ;
  RECT 32.200 5.940 32.400 6.140 ;
  LAYER VI3 ;
  RECT 31.800 6.340 32.000 6.540 ;
  LAYER VI3 ;
  RECT 31.800 5.940 32.000 6.140 ;
  LAYER VI3 ;
  RECT 31.400 6.340 31.600 6.540 ;
  LAYER VI3 ;
  RECT 31.400 5.940 31.600 6.140 ;
  LAYER VI3 ;
  RECT 31.000 6.340 31.200 6.540 ;
  LAYER VI3 ;
  RECT 31.000 5.940 31.200 6.140 ;
  LAYER VI3 ;
  RECT 30.600 6.340 30.800 6.540 ;
  LAYER VI3 ;
  RECT 30.600 5.940 30.800 6.140 ;
  LAYER VI3 ;
  RECT 30.200 6.340 30.400 6.540 ;
  LAYER VI3 ;
  RECT 30.200 5.940 30.400 6.140 ;
  LAYER VI3 ;
  RECT 29.800 6.340 30.000 6.540 ;
  LAYER VI3 ;
  RECT 29.800 5.940 30.000 6.140 ;
  LAYER VI3 ;
  RECT 29.400 6.340 29.600 6.540 ;
  LAYER VI3 ;
  RECT 29.400 5.940 29.600 6.140 ;
  LAYER VI3 ;
  RECT 29.000 6.340 29.200 6.540 ;
  LAYER VI3 ;
  RECT 29.000 5.940 29.200 6.140 ;
  LAYER VI3 ;
  RECT 28.600 6.340 28.800 6.540 ;
  LAYER VI3 ;
  RECT 28.600 5.940 28.800 6.140 ;
  LAYER VI3 ;
  RECT 28.200 6.340 28.400 6.540 ;
  LAYER VI3 ;
  RECT 28.200 5.940 28.400 6.140 ;
  LAYER VI3 ;
  RECT 49.280 5.880 57.280 6.740 ;
  LAYER VI3 ;
  RECT 56.880 6.340 57.080 6.540 ;
  LAYER VI3 ;
  RECT 56.880 5.940 57.080 6.140 ;
  LAYER VI3 ;
  RECT 56.480 6.340 56.680 6.540 ;
  LAYER VI3 ;
  RECT 56.480 5.940 56.680 6.140 ;
  LAYER VI3 ;
  RECT 56.080 6.340 56.280 6.540 ;
  LAYER VI3 ;
  RECT 56.080 5.940 56.280 6.140 ;
  LAYER VI3 ;
  RECT 55.680 6.340 55.880 6.540 ;
  LAYER VI3 ;
  RECT 55.680 5.940 55.880 6.140 ;
  LAYER VI3 ;
  RECT 55.280 6.340 55.480 6.540 ;
  LAYER VI3 ;
  RECT 55.280 5.940 55.480 6.140 ;
  LAYER VI3 ;
  RECT 54.880 6.340 55.080 6.540 ;
  LAYER VI3 ;
  RECT 54.880 5.940 55.080 6.140 ;
  LAYER VI3 ;
  RECT 54.480 6.340 54.680 6.540 ;
  LAYER VI3 ;
  RECT 54.480 5.940 54.680 6.140 ;
  LAYER VI3 ;
  RECT 54.080 6.340 54.280 6.540 ;
  LAYER VI3 ;
  RECT 54.080 5.940 54.280 6.140 ;
  LAYER VI3 ;
  RECT 53.680 6.340 53.880 6.540 ;
  LAYER VI3 ;
  RECT 53.680 5.940 53.880 6.140 ;
  LAYER VI3 ;
  RECT 53.280 6.340 53.480 6.540 ;
  LAYER VI3 ;
  RECT 53.280 5.940 53.480 6.140 ;
  LAYER VI3 ;
  RECT 52.880 6.340 53.080 6.540 ;
  LAYER VI3 ;
  RECT 52.880 5.940 53.080 6.140 ;
  LAYER VI3 ;
  RECT 52.480 6.340 52.680 6.540 ;
  LAYER VI3 ;
  RECT 52.480 5.940 52.680 6.140 ;
  LAYER VI3 ;
  RECT 52.080 6.340 52.280 6.540 ;
  LAYER VI3 ;
  RECT 52.080 5.940 52.280 6.140 ;
  LAYER VI3 ;
  RECT 51.680 6.340 51.880 6.540 ;
  LAYER VI3 ;
  RECT 51.680 5.940 51.880 6.140 ;
  LAYER VI3 ;
  RECT 51.280 6.340 51.480 6.540 ;
  LAYER VI3 ;
  RECT 51.280 5.940 51.480 6.140 ;
  LAYER VI3 ;
  RECT 50.880 6.340 51.080 6.540 ;
  LAYER VI3 ;
  RECT 50.880 5.940 51.080 6.140 ;
  LAYER VI3 ;
  RECT 50.480 6.340 50.680 6.540 ;
  LAYER VI3 ;
  RECT 50.480 5.940 50.680 6.140 ;
  LAYER VI3 ;
  RECT 50.080 6.340 50.280 6.540 ;
  LAYER VI3 ;
  RECT 50.080 5.940 50.280 6.140 ;
  LAYER VI3 ;
  RECT 49.680 6.340 49.880 6.540 ;
  LAYER VI3 ;
  RECT 49.680 5.940 49.880 6.140 ;
  LAYER VI3 ;
  RECT 49.280 6.340 49.480 6.540 ;
  LAYER VI3 ;
  RECT 49.280 5.940 49.480 6.140 ;
  LAYER VI3 ;
  RECT 69.120 5.880 77.120 6.740 ;
  LAYER VI3 ;
  RECT 76.720 6.340 76.920 6.540 ;
  LAYER VI3 ;
  RECT 76.720 5.940 76.920 6.140 ;
  LAYER VI3 ;
  RECT 76.320 6.340 76.520 6.540 ;
  LAYER VI3 ;
  RECT 76.320 5.940 76.520 6.140 ;
  LAYER VI3 ;
  RECT 75.920 6.340 76.120 6.540 ;
  LAYER VI3 ;
  RECT 75.920 5.940 76.120 6.140 ;
  LAYER VI3 ;
  RECT 75.520 6.340 75.720 6.540 ;
  LAYER VI3 ;
  RECT 75.520 5.940 75.720 6.140 ;
  LAYER VI3 ;
  RECT 75.120 6.340 75.320 6.540 ;
  LAYER VI3 ;
  RECT 75.120 5.940 75.320 6.140 ;
  LAYER VI3 ;
  RECT 74.720 6.340 74.920 6.540 ;
  LAYER VI3 ;
  RECT 74.720 5.940 74.920 6.140 ;
  LAYER VI3 ;
  RECT 74.320 6.340 74.520 6.540 ;
  LAYER VI3 ;
  RECT 74.320 5.940 74.520 6.140 ;
  LAYER VI3 ;
  RECT 73.920 6.340 74.120 6.540 ;
  LAYER VI3 ;
  RECT 73.920 5.940 74.120 6.140 ;
  LAYER VI3 ;
  RECT 73.520 6.340 73.720 6.540 ;
  LAYER VI3 ;
  RECT 73.520 5.940 73.720 6.140 ;
  LAYER VI3 ;
  RECT 73.120 6.340 73.320 6.540 ;
  LAYER VI3 ;
  RECT 73.120 5.940 73.320 6.140 ;
  LAYER VI3 ;
  RECT 72.720 6.340 72.920 6.540 ;
  LAYER VI3 ;
  RECT 72.720 5.940 72.920 6.140 ;
  LAYER VI3 ;
  RECT 72.320 6.340 72.520 6.540 ;
  LAYER VI3 ;
  RECT 72.320 5.940 72.520 6.140 ;
  LAYER VI3 ;
  RECT 71.920 6.340 72.120 6.540 ;
  LAYER VI3 ;
  RECT 71.920 5.940 72.120 6.140 ;
  LAYER VI3 ;
  RECT 71.520 6.340 71.720 6.540 ;
  LAYER VI3 ;
  RECT 71.520 5.940 71.720 6.140 ;
  LAYER VI3 ;
  RECT 71.120 6.340 71.320 6.540 ;
  LAYER VI3 ;
  RECT 71.120 5.940 71.320 6.140 ;
  LAYER VI3 ;
  RECT 70.720 6.340 70.920 6.540 ;
  LAYER VI3 ;
  RECT 70.720 5.940 70.920 6.140 ;
  LAYER VI3 ;
  RECT 70.320 6.340 70.520 6.540 ;
  LAYER VI3 ;
  RECT 70.320 5.940 70.520 6.140 ;
  LAYER VI3 ;
  RECT 69.920 6.340 70.120 6.540 ;
  LAYER VI3 ;
  RECT 69.920 5.940 70.120 6.140 ;
  LAYER VI3 ;
  RECT 69.520 6.340 69.720 6.540 ;
  LAYER VI3 ;
  RECT 69.520 5.940 69.720 6.140 ;
  LAYER VI3 ;
  RECT 69.120 6.340 69.320 6.540 ;
  LAYER VI3 ;
  RECT 69.120 5.940 69.320 6.140 ;
  LAYER VI3 ;
  RECT 90.200 5.880 98.200 6.740 ;
  LAYER VI3 ;
  RECT 97.800 6.340 98.000 6.540 ;
  LAYER VI3 ;
  RECT 97.800 5.940 98.000 6.140 ;
  LAYER VI3 ;
  RECT 97.400 6.340 97.600 6.540 ;
  LAYER VI3 ;
  RECT 97.400 5.940 97.600 6.140 ;
  LAYER VI3 ;
  RECT 97.000 6.340 97.200 6.540 ;
  LAYER VI3 ;
  RECT 97.000 5.940 97.200 6.140 ;
  LAYER VI3 ;
  RECT 96.600 6.340 96.800 6.540 ;
  LAYER VI3 ;
  RECT 96.600 5.940 96.800 6.140 ;
  LAYER VI3 ;
  RECT 96.200 6.340 96.400 6.540 ;
  LAYER VI3 ;
  RECT 96.200 5.940 96.400 6.140 ;
  LAYER VI3 ;
  RECT 95.800 6.340 96.000 6.540 ;
  LAYER VI3 ;
  RECT 95.800 5.940 96.000 6.140 ;
  LAYER VI3 ;
  RECT 95.400 6.340 95.600 6.540 ;
  LAYER VI3 ;
  RECT 95.400 5.940 95.600 6.140 ;
  LAYER VI3 ;
  RECT 95.000 6.340 95.200 6.540 ;
  LAYER VI3 ;
  RECT 95.000 5.940 95.200 6.140 ;
  LAYER VI3 ;
  RECT 94.600 6.340 94.800 6.540 ;
  LAYER VI3 ;
  RECT 94.600 5.940 94.800 6.140 ;
  LAYER VI3 ;
  RECT 94.200 6.340 94.400 6.540 ;
  LAYER VI3 ;
  RECT 94.200 5.940 94.400 6.140 ;
  LAYER VI3 ;
  RECT 93.800 6.340 94.000 6.540 ;
  LAYER VI3 ;
  RECT 93.800 5.940 94.000 6.140 ;
  LAYER VI3 ;
  RECT 93.400 6.340 93.600 6.540 ;
  LAYER VI3 ;
  RECT 93.400 5.940 93.600 6.140 ;
  LAYER VI3 ;
  RECT 93.000 6.340 93.200 6.540 ;
  LAYER VI3 ;
  RECT 93.000 5.940 93.200 6.140 ;
  LAYER VI3 ;
  RECT 92.600 6.340 92.800 6.540 ;
  LAYER VI3 ;
  RECT 92.600 5.940 92.800 6.140 ;
  LAYER VI3 ;
  RECT 92.200 6.340 92.400 6.540 ;
  LAYER VI3 ;
  RECT 92.200 5.940 92.400 6.140 ;
  LAYER VI3 ;
  RECT 91.800 6.340 92.000 6.540 ;
  LAYER VI3 ;
  RECT 91.800 5.940 92.000 6.140 ;
  LAYER VI3 ;
  RECT 91.400 6.340 91.600 6.540 ;
  LAYER VI3 ;
  RECT 91.400 5.940 91.600 6.140 ;
  LAYER VI3 ;
  RECT 91.000 6.340 91.200 6.540 ;
  LAYER VI3 ;
  RECT 91.000 5.940 91.200 6.140 ;
  LAYER VI3 ;
  RECT 90.600 6.340 90.800 6.540 ;
  LAYER VI3 ;
  RECT 90.600 5.940 90.800 6.140 ;
  LAYER VI3 ;
  RECT 90.200 6.340 90.400 6.540 ;
  LAYER VI3 ;
  RECT 90.200 5.940 90.400 6.140 ;
  LAYER VI3 ;
  RECT 110.040 5.880 118.040 6.740 ;
  LAYER VI3 ;
  RECT 117.640 6.340 117.840 6.540 ;
  LAYER VI3 ;
  RECT 117.640 5.940 117.840 6.140 ;
  LAYER VI3 ;
  RECT 117.240 6.340 117.440 6.540 ;
  LAYER VI3 ;
  RECT 117.240 5.940 117.440 6.140 ;
  LAYER VI3 ;
  RECT 116.840 6.340 117.040 6.540 ;
  LAYER VI3 ;
  RECT 116.840 5.940 117.040 6.140 ;
  LAYER VI3 ;
  RECT 116.440 6.340 116.640 6.540 ;
  LAYER VI3 ;
  RECT 116.440 5.940 116.640 6.140 ;
  LAYER VI3 ;
  RECT 116.040 6.340 116.240 6.540 ;
  LAYER VI3 ;
  RECT 116.040 5.940 116.240 6.140 ;
  LAYER VI3 ;
  RECT 115.640 6.340 115.840 6.540 ;
  LAYER VI3 ;
  RECT 115.640 5.940 115.840 6.140 ;
  LAYER VI3 ;
  RECT 115.240 6.340 115.440 6.540 ;
  LAYER VI3 ;
  RECT 115.240 5.940 115.440 6.140 ;
  LAYER VI3 ;
  RECT 114.840 6.340 115.040 6.540 ;
  LAYER VI3 ;
  RECT 114.840 5.940 115.040 6.140 ;
  LAYER VI3 ;
  RECT 114.440 6.340 114.640 6.540 ;
  LAYER VI3 ;
  RECT 114.440 5.940 114.640 6.140 ;
  LAYER VI3 ;
  RECT 114.040 6.340 114.240 6.540 ;
  LAYER VI3 ;
  RECT 114.040 5.940 114.240 6.140 ;
  LAYER VI3 ;
  RECT 113.640 6.340 113.840 6.540 ;
  LAYER VI3 ;
  RECT 113.640 5.940 113.840 6.140 ;
  LAYER VI3 ;
  RECT 113.240 6.340 113.440 6.540 ;
  LAYER VI3 ;
  RECT 113.240 5.940 113.440 6.140 ;
  LAYER VI3 ;
  RECT 112.840 6.340 113.040 6.540 ;
  LAYER VI3 ;
  RECT 112.840 5.940 113.040 6.140 ;
  LAYER VI3 ;
  RECT 112.440 6.340 112.640 6.540 ;
  LAYER VI3 ;
  RECT 112.440 5.940 112.640 6.140 ;
  LAYER VI3 ;
  RECT 112.040 6.340 112.240 6.540 ;
  LAYER VI3 ;
  RECT 112.040 5.940 112.240 6.140 ;
  LAYER VI3 ;
  RECT 111.640 6.340 111.840 6.540 ;
  LAYER VI3 ;
  RECT 111.640 5.940 111.840 6.140 ;
  LAYER VI3 ;
  RECT 111.240 6.340 111.440 6.540 ;
  LAYER VI3 ;
  RECT 111.240 5.940 111.440 6.140 ;
  LAYER VI3 ;
  RECT 110.840 6.340 111.040 6.540 ;
  LAYER VI3 ;
  RECT 110.840 5.940 111.040 6.140 ;
  LAYER VI3 ;
  RECT 110.440 6.340 110.640 6.540 ;
  LAYER VI3 ;
  RECT 110.440 5.940 110.640 6.140 ;
  LAYER VI3 ;
  RECT 110.040 6.340 110.240 6.540 ;
  LAYER VI3 ;
  RECT 110.040 5.940 110.240 6.140 ;
  LAYER VI3 ;
  RECT 131.120 5.880 139.120 6.740 ;
  LAYER VI3 ;
  RECT 138.720 6.340 138.920 6.540 ;
  LAYER VI3 ;
  RECT 138.720 5.940 138.920 6.140 ;
  LAYER VI3 ;
  RECT 138.320 6.340 138.520 6.540 ;
  LAYER VI3 ;
  RECT 138.320 5.940 138.520 6.140 ;
  LAYER VI3 ;
  RECT 137.920 6.340 138.120 6.540 ;
  LAYER VI3 ;
  RECT 137.920 5.940 138.120 6.140 ;
  LAYER VI3 ;
  RECT 137.520 6.340 137.720 6.540 ;
  LAYER VI3 ;
  RECT 137.520 5.940 137.720 6.140 ;
  LAYER VI3 ;
  RECT 137.120 6.340 137.320 6.540 ;
  LAYER VI3 ;
  RECT 137.120 5.940 137.320 6.140 ;
  LAYER VI3 ;
  RECT 136.720 6.340 136.920 6.540 ;
  LAYER VI3 ;
  RECT 136.720 5.940 136.920 6.140 ;
  LAYER VI3 ;
  RECT 136.320 6.340 136.520 6.540 ;
  LAYER VI3 ;
  RECT 136.320 5.940 136.520 6.140 ;
  LAYER VI3 ;
  RECT 135.920 6.340 136.120 6.540 ;
  LAYER VI3 ;
  RECT 135.920 5.940 136.120 6.140 ;
  LAYER VI3 ;
  RECT 135.520 6.340 135.720 6.540 ;
  LAYER VI3 ;
  RECT 135.520 5.940 135.720 6.140 ;
  LAYER VI3 ;
  RECT 135.120 6.340 135.320 6.540 ;
  LAYER VI3 ;
  RECT 135.120 5.940 135.320 6.140 ;
  LAYER VI3 ;
  RECT 134.720 6.340 134.920 6.540 ;
  LAYER VI3 ;
  RECT 134.720 5.940 134.920 6.140 ;
  LAYER VI3 ;
  RECT 134.320 6.340 134.520 6.540 ;
  LAYER VI3 ;
  RECT 134.320 5.940 134.520 6.140 ;
  LAYER VI3 ;
  RECT 133.920 6.340 134.120 6.540 ;
  LAYER VI3 ;
  RECT 133.920 5.940 134.120 6.140 ;
  LAYER VI3 ;
  RECT 133.520 6.340 133.720 6.540 ;
  LAYER VI3 ;
  RECT 133.520 5.940 133.720 6.140 ;
  LAYER VI3 ;
  RECT 133.120 6.340 133.320 6.540 ;
  LAYER VI3 ;
  RECT 133.120 5.940 133.320 6.140 ;
  LAYER VI3 ;
  RECT 132.720 6.340 132.920 6.540 ;
  LAYER VI3 ;
  RECT 132.720 5.940 132.920 6.140 ;
  LAYER VI3 ;
  RECT 132.320 6.340 132.520 6.540 ;
  LAYER VI3 ;
  RECT 132.320 5.940 132.520 6.140 ;
  LAYER VI3 ;
  RECT 131.920 6.340 132.120 6.540 ;
  LAYER VI3 ;
  RECT 131.920 5.940 132.120 6.140 ;
  LAYER VI3 ;
  RECT 131.520 6.340 131.720 6.540 ;
  LAYER VI3 ;
  RECT 131.520 5.940 131.720 6.140 ;
  LAYER VI3 ;
  RECT 131.120 6.340 131.320 6.540 ;
  LAYER VI3 ;
  RECT 131.120 5.940 131.320 6.140 ;
  LAYER VI3 ;
  RECT 150.960 5.880 158.960 6.740 ;
  LAYER VI3 ;
  RECT 158.560 6.340 158.760 6.540 ;
  LAYER VI3 ;
  RECT 158.560 5.940 158.760 6.140 ;
  LAYER VI3 ;
  RECT 158.160 6.340 158.360 6.540 ;
  LAYER VI3 ;
  RECT 158.160 5.940 158.360 6.140 ;
  LAYER VI3 ;
  RECT 157.760 6.340 157.960 6.540 ;
  LAYER VI3 ;
  RECT 157.760 5.940 157.960 6.140 ;
  LAYER VI3 ;
  RECT 157.360 6.340 157.560 6.540 ;
  LAYER VI3 ;
  RECT 157.360 5.940 157.560 6.140 ;
  LAYER VI3 ;
  RECT 156.960 6.340 157.160 6.540 ;
  LAYER VI3 ;
  RECT 156.960 5.940 157.160 6.140 ;
  LAYER VI3 ;
  RECT 156.560 6.340 156.760 6.540 ;
  LAYER VI3 ;
  RECT 156.560 5.940 156.760 6.140 ;
  LAYER VI3 ;
  RECT 156.160 6.340 156.360 6.540 ;
  LAYER VI3 ;
  RECT 156.160 5.940 156.360 6.140 ;
  LAYER VI3 ;
  RECT 155.760 6.340 155.960 6.540 ;
  LAYER VI3 ;
  RECT 155.760 5.940 155.960 6.140 ;
  LAYER VI3 ;
  RECT 155.360 6.340 155.560 6.540 ;
  LAYER VI3 ;
  RECT 155.360 5.940 155.560 6.140 ;
  LAYER VI3 ;
  RECT 154.960 6.340 155.160 6.540 ;
  LAYER VI3 ;
  RECT 154.960 5.940 155.160 6.140 ;
  LAYER VI3 ;
  RECT 154.560 6.340 154.760 6.540 ;
  LAYER VI3 ;
  RECT 154.560 5.940 154.760 6.140 ;
  LAYER VI3 ;
  RECT 154.160 6.340 154.360 6.540 ;
  LAYER VI3 ;
  RECT 154.160 5.940 154.360 6.140 ;
  LAYER VI3 ;
  RECT 153.760 6.340 153.960 6.540 ;
  LAYER VI3 ;
  RECT 153.760 5.940 153.960 6.140 ;
  LAYER VI3 ;
  RECT 153.360 6.340 153.560 6.540 ;
  LAYER VI3 ;
  RECT 153.360 5.940 153.560 6.140 ;
  LAYER VI3 ;
  RECT 152.960 6.340 153.160 6.540 ;
  LAYER VI3 ;
  RECT 152.960 5.940 153.160 6.140 ;
  LAYER VI3 ;
  RECT 152.560 6.340 152.760 6.540 ;
  LAYER VI3 ;
  RECT 152.560 5.940 152.760 6.140 ;
  LAYER VI3 ;
  RECT 152.160 6.340 152.360 6.540 ;
  LAYER VI3 ;
  RECT 152.160 5.940 152.360 6.140 ;
  LAYER VI3 ;
  RECT 151.760 6.340 151.960 6.540 ;
  LAYER VI3 ;
  RECT 151.760 5.940 151.960 6.140 ;
  LAYER VI3 ;
  RECT 151.360 6.340 151.560 6.540 ;
  LAYER VI3 ;
  RECT 151.360 5.940 151.560 6.140 ;
  LAYER VI3 ;
  RECT 150.960 6.340 151.160 6.540 ;
  LAYER VI3 ;
  RECT 150.960 5.940 151.160 6.140 ;
  LAYER VI3 ;
  RECT 172.040 5.880 180.040 6.740 ;
  LAYER VI3 ;
  RECT 179.640 6.340 179.840 6.540 ;
  LAYER VI3 ;
  RECT 179.640 5.940 179.840 6.140 ;
  LAYER VI3 ;
  RECT 179.240 6.340 179.440 6.540 ;
  LAYER VI3 ;
  RECT 179.240 5.940 179.440 6.140 ;
  LAYER VI3 ;
  RECT 178.840 6.340 179.040 6.540 ;
  LAYER VI3 ;
  RECT 178.840 5.940 179.040 6.140 ;
  LAYER VI3 ;
  RECT 178.440 6.340 178.640 6.540 ;
  LAYER VI3 ;
  RECT 178.440 5.940 178.640 6.140 ;
  LAYER VI3 ;
  RECT 178.040 6.340 178.240 6.540 ;
  LAYER VI3 ;
  RECT 178.040 5.940 178.240 6.140 ;
  LAYER VI3 ;
  RECT 177.640 6.340 177.840 6.540 ;
  LAYER VI3 ;
  RECT 177.640 5.940 177.840 6.140 ;
  LAYER VI3 ;
  RECT 177.240 6.340 177.440 6.540 ;
  LAYER VI3 ;
  RECT 177.240 5.940 177.440 6.140 ;
  LAYER VI3 ;
  RECT 176.840 6.340 177.040 6.540 ;
  LAYER VI3 ;
  RECT 176.840 5.940 177.040 6.140 ;
  LAYER VI3 ;
  RECT 176.440 6.340 176.640 6.540 ;
  LAYER VI3 ;
  RECT 176.440 5.940 176.640 6.140 ;
  LAYER VI3 ;
  RECT 176.040 6.340 176.240 6.540 ;
  LAYER VI3 ;
  RECT 176.040 5.940 176.240 6.140 ;
  LAYER VI3 ;
  RECT 175.640 6.340 175.840 6.540 ;
  LAYER VI3 ;
  RECT 175.640 5.940 175.840 6.140 ;
  LAYER VI3 ;
  RECT 175.240 6.340 175.440 6.540 ;
  LAYER VI3 ;
  RECT 175.240 5.940 175.440 6.140 ;
  LAYER VI3 ;
  RECT 174.840 6.340 175.040 6.540 ;
  LAYER VI3 ;
  RECT 174.840 5.940 175.040 6.140 ;
  LAYER VI3 ;
  RECT 174.440 6.340 174.640 6.540 ;
  LAYER VI3 ;
  RECT 174.440 5.940 174.640 6.140 ;
  LAYER VI3 ;
  RECT 174.040 6.340 174.240 6.540 ;
  LAYER VI3 ;
  RECT 174.040 5.940 174.240 6.140 ;
  LAYER VI3 ;
  RECT 173.640 6.340 173.840 6.540 ;
  LAYER VI3 ;
  RECT 173.640 5.940 173.840 6.140 ;
  LAYER VI3 ;
  RECT 173.240 6.340 173.440 6.540 ;
  LAYER VI3 ;
  RECT 173.240 5.940 173.440 6.140 ;
  LAYER VI3 ;
  RECT 172.840 6.340 173.040 6.540 ;
  LAYER VI3 ;
  RECT 172.840 5.940 173.040 6.140 ;
  LAYER VI3 ;
  RECT 172.440 6.340 172.640 6.540 ;
  LAYER VI3 ;
  RECT 172.440 5.940 172.640 6.140 ;
  LAYER VI3 ;
  RECT 172.040 6.340 172.240 6.540 ;
  LAYER VI3 ;
  RECT 172.040 5.940 172.240 6.140 ;
  LAYER VI3 ;
  RECT 191.880 5.880 199.880 6.740 ;
  LAYER VI3 ;
  RECT 199.480 6.340 199.680 6.540 ;
  LAYER VI3 ;
  RECT 199.480 5.940 199.680 6.140 ;
  LAYER VI3 ;
  RECT 199.080 6.340 199.280 6.540 ;
  LAYER VI3 ;
  RECT 199.080 5.940 199.280 6.140 ;
  LAYER VI3 ;
  RECT 198.680 6.340 198.880 6.540 ;
  LAYER VI3 ;
  RECT 198.680 5.940 198.880 6.140 ;
  LAYER VI3 ;
  RECT 198.280 6.340 198.480 6.540 ;
  LAYER VI3 ;
  RECT 198.280 5.940 198.480 6.140 ;
  LAYER VI3 ;
  RECT 197.880 6.340 198.080 6.540 ;
  LAYER VI3 ;
  RECT 197.880 5.940 198.080 6.140 ;
  LAYER VI3 ;
  RECT 197.480 6.340 197.680 6.540 ;
  LAYER VI3 ;
  RECT 197.480 5.940 197.680 6.140 ;
  LAYER VI3 ;
  RECT 197.080 6.340 197.280 6.540 ;
  LAYER VI3 ;
  RECT 197.080 5.940 197.280 6.140 ;
  LAYER VI3 ;
  RECT 196.680 6.340 196.880 6.540 ;
  LAYER VI3 ;
  RECT 196.680 5.940 196.880 6.140 ;
  LAYER VI3 ;
  RECT 196.280 6.340 196.480 6.540 ;
  LAYER VI3 ;
  RECT 196.280 5.940 196.480 6.140 ;
  LAYER VI3 ;
  RECT 195.880 6.340 196.080 6.540 ;
  LAYER VI3 ;
  RECT 195.880 5.940 196.080 6.140 ;
  LAYER VI3 ;
  RECT 195.480 6.340 195.680 6.540 ;
  LAYER VI3 ;
  RECT 195.480 5.940 195.680 6.140 ;
  LAYER VI3 ;
  RECT 195.080 6.340 195.280 6.540 ;
  LAYER VI3 ;
  RECT 195.080 5.940 195.280 6.140 ;
  LAYER VI3 ;
  RECT 194.680 6.340 194.880 6.540 ;
  LAYER VI3 ;
  RECT 194.680 5.940 194.880 6.140 ;
  LAYER VI3 ;
  RECT 194.280 6.340 194.480 6.540 ;
  LAYER VI3 ;
  RECT 194.280 5.940 194.480 6.140 ;
  LAYER VI3 ;
  RECT 193.880 6.340 194.080 6.540 ;
  LAYER VI3 ;
  RECT 193.880 5.940 194.080 6.140 ;
  LAYER VI3 ;
  RECT 193.480 6.340 193.680 6.540 ;
  LAYER VI3 ;
  RECT 193.480 5.940 193.680 6.140 ;
  LAYER VI3 ;
  RECT 193.080 6.340 193.280 6.540 ;
  LAYER VI3 ;
  RECT 193.080 5.940 193.280 6.140 ;
  LAYER VI3 ;
  RECT 192.680 6.340 192.880 6.540 ;
  LAYER VI3 ;
  RECT 192.680 5.940 192.880 6.140 ;
  LAYER VI3 ;
  RECT 192.280 6.340 192.480 6.540 ;
  LAYER VI3 ;
  RECT 192.280 5.940 192.480 6.140 ;
  LAYER VI3 ;
  RECT 191.880 6.340 192.080 6.540 ;
  LAYER VI3 ;
  RECT 191.880 5.940 192.080 6.140 ;
  LAYER VI3 ;
  RECT 212.960 5.880 220.960 6.740 ;
  LAYER VI3 ;
  RECT 220.560 6.340 220.760 6.540 ;
  LAYER VI3 ;
  RECT 220.560 5.940 220.760 6.140 ;
  LAYER VI3 ;
  RECT 220.160 6.340 220.360 6.540 ;
  LAYER VI3 ;
  RECT 220.160 5.940 220.360 6.140 ;
  LAYER VI3 ;
  RECT 219.760 6.340 219.960 6.540 ;
  LAYER VI3 ;
  RECT 219.760 5.940 219.960 6.140 ;
  LAYER VI3 ;
  RECT 219.360 6.340 219.560 6.540 ;
  LAYER VI3 ;
  RECT 219.360 5.940 219.560 6.140 ;
  LAYER VI3 ;
  RECT 218.960 6.340 219.160 6.540 ;
  LAYER VI3 ;
  RECT 218.960 5.940 219.160 6.140 ;
  LAYER VI3 ;
  RECT 218.560 6.340 218.760 6.540 ;
  LAYER VI3 ;
  RECT 218.560 5.940 218.760 6.140 ;
  LAYER VI3 ;
  RECT 218.160 6.340 218.360 6.540 ;
  LAYER VI3 ;
  RECT 218.160 5.940 218.360 6.140 ;
  LAYER VI3 ;
  RECT 217.760 6.340 217.960 6.540 ;
  LAYER VI3 ;
  RECT 217.760 5.940 217.960 6.140 ;
  LAYER VI3 ;
  RECT 217.360 6.340 217.560 6.540 ;
  LAYER VI3 ;
  RECT 217.360 5.940 217.560 6.140 ;
  LAYER VI3 ;
  RECT 216.960 6.340 217.160 6.540 ;
  LAYER VI3 ;
  RECT 216.960 5.940 217.160 6.140 ;
  LAYER VI3 ;
  RECT 216.560 6.340 216.760 6.540 ;
  LAYER VI3 ;
  RECT 216.560 5.940 216.760 6.140 ;
  LAYER VI3 ;
  RECT 216.160 6.340 216.360 6.540 ;
  LAYER VI3 ;
  RECT 216.160 5.940 216.360 6.140 ;
  LAYER VI3 ;
  RECT 215.760 6.340 215.960 6.540 ;
  LAYER VI3 ;
  RECT 215.760 5.940 215.960 6.140 ;
  LAYER VI3 ;
  RECT 215.360 6.340 215.560 6.540 ;
  LAYER VI3 ;
  RECT 215.360 5.940 215.560 6.140 ;
  LAYER VI3 ;
  RECT 214.960 6.340 215.160 6.540 ;
  LAYER VI3 ;
  RECT 214.960 5.940 215.160 6.140 ;
  LAYER VI3 ;
  RECT 214.560 6.340 214.760 6.540 ;
  LAYER VI3 ;
  RECT 214.560 5.940 214.760 6.140 ;
  LAYER VI3 ;
  RECT 214.160 6.340 214.360 6.540 ;
  LAYER VI3 ;
  RECT 214.160 5.940 214.360 6.140 ;
  LAYER VI3 ;
  RECT 213.760 6.340 213.960 6.540 ;
  LAYER VI3 ;
  RECT 213.760 5.940 213.960 6.140 ;
  LAYER VI3 ;
  RECT 213.360 6.340 213.560 6.540 ;
  LAYER VI3 ;
  RECT 213.360 5.940 213.560 6.140 ;
  LAYER VI3 ;
  RECT 212.960 6.340 213.160 6.540 ;
  LAYER VI3 ;
  RECT 212.960 5.940 213.160 6.140 ;
  LAYER VI3 ;
  RECT 232.800 5.880 240.800 6.740 ;
  LAYER VI3 ;
  RECT 240.400 6.340 240.600 6.540 ;
  LAYER VI3 ;
  RECT 240.400 5.940 240.600 6.140 ;
  LAYER VI3 ;
  RECT 240.000 6.340 240.200 6.540 ;
  LAYER VI3 ;
  RECT 240.000 5.940 240.200 6.140 ;
  LAYER VI3 ;
  RECT 239.600 6.340 239.800 6.540 ;
  LAYER VI3 ;
  RECT 239.600 5.940 239.800 6.140 ;
  LAYER VI3 ;
  RECT 239.200 6.340 239.400 6.540 ;
  LAYER VI3 ;
  RECT 239.200 5.940 239.400 6.140 ;
  LAYER VI3 ;
  RECT 238.800 6.340 239.000 6.540 ;
  LAYER VI3 ;
  RECT 238.800 5.940 239.000 6.140 ;
  LAYER VI3 ;
  RECT 238.400 6.340 238.600 6.540 ;
  LAYER VI3 ;
  RECT 238.400 5.940 238.600 6.140 ;
  LAYER VI3 ;
  RECT 238.000 6.340 238.200 6.540 ;
  LAYER VI3 ;
  RECT 238.000 5.940 238.200 6.140 ;
  LAYER VI3 ;
  RECT 237.600 6.340 237.800 6.540 ;
  LAYER VI3 ;
  RECT 237.600 5.940 237.800 6.140 ;
  LAYER VI3 ;
  RECT 237.200 6.340 237.400 6.540 ;
  LAYER VI3 ;
  RECT 237.200 5.940 237.400 6.140 ;
  LAYER VI3 ;
  RECT 236.800 6.340 237.000 6.540 ;
  LAYER VI3 ;
  RECT 236.800 5.940 237.000 6.140 ;
  LAYER VI3 ;
  RECT 236.400 6.340 236.600 6.540 ;
  LAYER VI3 ;
  RECT 236.400 5.940 236.600 6.140 ;
  LAYER VI3 ;
  RECT 236.000 6.340 236.200 6.540 ;
  LAYER VI3 ;
  RECT 236.000 5.940 236.200 6.140 ;
  LAYER VI3 ;
  RECT 235.600 6.340 235.800 6.540 ;
  LAYER VI3 ;
  RECT 235.600 5.940 235.800 6.140 ;
  LAYER VI3 ;
  RECT 235.200 6.340 235.400 6.540 ;
  LAYER VI3 ;
  RECT 235.200 5.940 235.400 6.140 ;
  LAYER VI3 ;
  RECT 234.800 6.340 235.000 6.540 ;
  LAYER VI3 ;
  RECT 234.800 5.940 235.000 6.140 ;
  LAYER VI3 ;
  RECT 234.400 6.340 234.600 6.540 ;
  LAYER VI3 ;
  RECT 234.400 5.940 234.600 6.140 ;
  LAYER VI3 ;
  RECT 234.000 6.340 234.200 6.540 ;
  LAYER VI3 ;
  RECT 234.000 5.940 234.200 6.140 ;
  LAYER VI3 ;
  RECT 233.600 6.340 233.800 6.540 ;
  LAYER VI3 ;
  RECT 233.600 5.940 233.800 6.140 ;
  LAYER VI3 ;
  RECT 233.200 6.340 233.400 6.540 ;
  LAYER VI3 ;
  RECT 233.200 5.940 233.400 6.140 ;
  LAYER VI3 ;
  RECT 232.800 6.340 233.000 6.540 ;
  LAYER VI3 ;
  RECT 232.800 5.940 233.000 6.140 ;
  LAYER VI3 ;
  RECT 253.880 5.880 261.880 6.740 ;
  LAYER VI3 ;
  RECT 261.480 6.340 261.680 6.540 ;
  LAYER VI3 ;
  RECT 261.480 5.940 261.680 6.140 ;
  LAYER VI3 ;
  RECT 261.080 6.340 261.280 6.540 ;
  LAYER VI3 ;
  RECT 261.080 5.940 261.280 6.140 ;
  LAYER VI3 ;
  RECT 260.680 6.340 260.880 6.540 ;
  LAYER VI3 ;
  RECT 260.680 5.940 260.880 6.140 ;
  LAYER VI3 ;
  RECT 260.280 6.340 260.480 6.540 ;
  LAYER VI3 ;
  RECT 260.280 5.940 260.480 6.140 ;
  LAYER VI3 ;
  RECT 259.880 6.340 260.080 6.540 ;
  LAYER VI3 ;
  RECT 259.880 5.940 260.080 6.140 ;
  LAYER VI3 ;
  RECT 259.480 6.340 259.680 6.540 ;
  LAYER VI3 ;
  RECT 259.480 5.940 259.680 6.140 ;
  LAYER VI3 ;
  RECT 259.080 6.340 259.280 6.540 ;
  LAYER VI3 ;
  RECT 259.080 5.940 259.280 6.140 ;
  LAYER VI3 ;
  RECT 258.680 6.340 258.880 6.540 ;
  LAYER VI3 ;
  RECT 258.680 5.940 258.880 6.140 ;
  LAYER VI3 ;
  RECT 258.280 6.340 258.480 6.540 ;
  LAYER VI3 ;
  RECT 258.280 5.940 258.480 6.140 ;
  LAYER VI3 ;
  RECT 257.880 6.340 258.080 6.540 ;
  LAYER VI3 ;
  RECT 257.880 5.940 258.080 6.140 ;
  LAYER VI3 ;
  RECT 257.480 6.340 257.680 6.540 ;
  LAYER VI3 ;
  RECT 257.480 5.940 257.680 6.140 ;
  LAYER VI3 ;
  RECT 257.080 6.340 257.280 6.540 ;
  LAYER VI3 ;
  RECT 257.080 5.940 257.280 6.140 ;
  LAYER VI3 ;
  RECT 256.680 6.340 256.880 6.540 ;
  LAYER VI3 ;
  RECT 256.680 5.940 256.880 6.140 ;
  LAYER VI3 ;
  RECT 256.280 6.340 256.480 6.540 ;
  LAYER VI3 ;
  RECT 256.280 5.940 256.480 6.140 ;
  LAYER VI3 ;
  RECT 255.880 6.340 256.080 6.540 ;
  LAYER VI3 ;
  RECT 255.880 5.940 256.080 6.140 ;
  LAYER VI3 ;
  RECT 255.480 6.340 255.680 6.540 ;
  LAYER VI3 ;
  RECT 255.480 5.940 255.680 6.140 ;
  LAYER VI3 ;
  RECT 255.080 6.340 255.280 6.540 ;
  LAYER VI3 ;
  RECT 255.080 5.940 255.280 6.140 ;
  LAYER VI3 ;
  RECT 254.680 6.340 254.880 6.540 ;
  LAYER VI3 ;
  RECT 254.680 5.940 254.880 6.140 ;
  LAYER VI3 ;
  RECT 254.280 6.340 254.480 6.540 ;
  LAYER VI3 ;
  RECT 254.280 5.940 254.480 6.140 ;
  LAYER VI3 ;
  RECT 253.880 6.340 254.080 6.540 ;
  LAYER VI3 ;
  RECT 253.880 5.940 254.080 6.140 ;
  LAYER VI3 ;
  RECT 273.720 5.880 281.720 6.740 ;
  LAYER VI3 ;
  RECT 281.320 6.340 281.520 6.540 ;
  LAYER VI3 ;
  RECT 281.320 5.940 281.520 6.140 ;
  LAYER VI3 ;
  RECT 280.920 6.340 281.120 6.540 ;
  LAYER VI3 ;
  RECT 280.920 5.940 281.120 6.140 ;
  LAYER VI3 ;
  RECT 280.520 6.340 280.720 6.540 ;
  LAYER VI3 ;
  RECT 280.520 5.940 280.720 6.140 ;
  LAYER VI3 ;
  RECT 280.120 6.340 280.320 6.540 ;
  LAYER VI3 ;
  RECT 280.120 5.940 280.320 6.140 ;
  LAYER VI3 ;
  RECT 279.720 6.340 279.920 6.540 ;
  LAYER VI3 ;
  RECT 279.720 5.940 279.920 6.140 ;
  LAYER VI3 ;
  RECT 279.320 6.340 279.520 6.540 ;
  LAYER VI3 ;
  RECT 279.320 5.940 279.520 6.140 ;
  LAYER VI3 ;
  RECT 278.920 6.340 279.120 6.540 ;
  LAYER VI3 ;
  RECT 278.920 5.940 279.120 6.140 ;
  LAYER VI3 ;
  RECT 278.520 6.340 278.720 6.540 ;
  LAYER VI3 ;
  RECT 278.520 5.940 278.720 6.140 ;
  LAYER VI3 ;
  RECT 278.120 6.340 278.320 6.540 ;
  LAYER VI3 ;
  RECT 278.120 5.940 278.320 6.140 ;
  LAYER VI3 ;
  RECT 277.720 6.340 277.920 6.540 ;
  LAYER VI3 ;
  RECT 277.720 5.940 277.920 6.140 ;
  LAYER VI3 ;
  RECT 277.320 6.340 277.520 6.540 ;
  LAYER VI3 ;
  RECT 277.320 5.940 277.520 6.140 ;
  LAYER VI3 ;
  RECT 276.920 6.340 277.120 6.540 ;
  LAYER VI3 ;
  RECT 276.920 5.940 277.120 6.140 ;
  LAYER VI3 ;
  RECT 276.520 6.340 276.720 6.540 ;
  LAYER VI3 ;
  RECT 276.520 5.940 276.720 6.140 ;
  LAYER VI3 ;
  RECT 276.120 6.340 276.320 6.540 ;
  LAYER VI3 ;
  RECT 276.120 5.940 276.320 6.140 ;
  LAYER VI3 ;
  RECT 275.720 6.340 275.920 6.540 ;
  LAYER VI3 ;
  RECT 275.720 5.940 275.920 6.140 ;
  LAYER VI3 ;
  RECT 275.320 6.340 275.520 6.540 ;
  LAYER VI3 ;
  RECT 275.320 5.940 275.520 6.140 ;
  LAYER VI3 ;
  RECT 274.920 6.340 275.120 6.540 ;
  LAYER VI3 ;
  RECT 274.920 5.940 275.120 6.140 ;
  LAYER VI3 ;
  RECT 274.520 6.340 274.720 6.540 ;
  LAYER VI3 ;
  RECT 274.520 5.940 274.720 6.140 ;
  LAYER VI3 ;
  RECT 274.120 6.340 274.320 6.540 ;
  LAYER VI3 ;
  RECT 274.120 5.940 274.320 6.140 ;
  LAYER VI3 ;
  RECT 273.720 6.340 273.920 6.540 ;
  LAYER VI3 ;
  RECT 273.720 5.940 273.920 6.140 ;
  LAYER VI3 ;
  RECT 294.800 5.880 302.800 6.740 ;
  LAYER VI3 ;
  RECT 302.400 6.340 302.600 6.540 ;
  LAYER VI3 ;
  RECT 302.400 5.940 302.600 6.140 ;
  LAYER VI3 ;
  RECT 302.000 6.340 302.200 6.540 ;
  LAYER VI3 ;
  RECT 302.000 5.940 302.200 6.140 ;
  LAYER VI3 ;
  RECT 301.600 6.340 301.800 6.540 ;
  LAYER VI3 ;
  RECT 301.600 5.940 301.800 6.140 ;
  LAYER VI3 ;
  RECT 301.200 6.340 301.400 6.540 ;
  LAYER VI3 ;
  RECT 301.200 5.940 301.400 6.140 ;
  LAYER VI3 ;
  RECT 300.800 6.340 301.000 6.540 ;
  LAYER VI3 ;
  RECT 300.800 5.940 301.000 6.140 ;
  LAYER VI3 ;
  RECT 300.400 6.340 300.600 6.540 ;
  LAYER VI3 ;
  RECT 300.400 5.940 300.600 6.140 ;
  LAYER VI3 ;
  RECT 300.000 6.340 300.200 6.540 ;
  LAYER VI3 ;
  RECT 300.000 5.940 300.200 6.140 ;
  LAYER VI3 ;
  RECT 299.600 6.340 299.800 6.540 ;
  LAYER VI3 ;
  RECT 299.600 5.940 299.800 6.140 ;
  LAYER VI3 ;
  RECT 299.200 6.340 299.400 6.540 ;
  LAYER VI3 ;
  RECT 299.200 5.940 299.400 6.140 ;
  LAYER VI3 ;
  RECT 298.800 6.340 299.000 6.540 ;
  LAYER VI3 ;
  RECT 298.800 5.940 299.000 6.140 ;
  LAYER VI3 ;
  RECT 298.400 6.340 298.600 6.540 ;
  LAYER VI3 ;
  RECT 298.400 5.940 298.600 6.140 ;
  LAYER VI3 ;
  RECT 298.000 6.340 298.200 6.540 ;
  LAYER VI3 ;
  RECT 298.000 5.940 298.200 6.140 ;
  LAYER VI3 ;
  RECT 297.600 6.340 297.800 6.540 ;
  LAYER VI3 ;
  RECT 297.600 5.940 297.800 6.140 ;
  LAYER VI3 ;
  RECT 297.200 6.340 297.400 6.540 ;
  LAYER VI3 ;
  RECT 297.200 5.940 297.400 6.140 ;
  LAYER VI3 ;
  RECT 296.800 6.340 297.000 6.540 ;
  LAYER VI3 ;
  RECT 296.800 5.940 297.000 6.140 ;
  LAYER VI3 ;
  RECT 296.400 6.340 296.600 6.540 ;
  LAYER VI3 ;
  RECT 296.400 5.940 296.600 6.140 ;
  LAYER VI3 ;
  RECT 296.000 6.340 296.200 6.540 ;
  LAYER VI3 ;
  RECT 296.000 5.940 296.200 6.140 ;
  LAYER VI3 ;
  RECT 295.600 6.340 295.800 6.540 ;
  LAYER VI3 ;
  RECT 295.600 5.940 295.800 6.140 ;
  LAYER VI3 ;
  RECT 295.200 6.340 295.400 6.540 ;
  LAYER VI3 ;
  RECT 295.200 5.940 295.400 6.140 ;
  LAYER VI3 ;
  RECT 294.800 6.340 295.000 6.540 ;
  LAYER VI3 ;
  RECT 294.800 5.940 295.000 6.140 ;
  LAYER VI3 ;
  RECT 314.640 5.880 322.640 6.740 ;
  LAYER VI3 ;
  RECT 322.240 6.340 322.440 6.540 ;
  LAYER VI3 ;
  RECT 322.240 5.940 322.440 6.140 ;
  LAYER VI3 ;
  RECT 321.840 6.340 322.040 6.540 ;
  LAYER VI3 ;
  RECT 321.840 5.940 322.040 6.140 ;
  LAYER VI3 ;
  RECT 321.440 6.340 321.640 6.540 ;
  LAYER VI3 ;
  RECT 321.440 5.940 321.640 6.140 ;
  LAYER VI3 ;
  RECT 321.040 6.340 321.240 6.540 ;
  LAYER VI3 ;
  RECT 321.040 5.940 321.240 6.140 ;
  LAYER VI3 ;
  RECT 320.640 6.340 320.840 6.540 ;
  LAYER VI3 ;
  RECT 320.640 5.940 320.840 6.140 ;
  LAYER VI3 ;
  RECT 320.240 6.340 320.440 6.540 ;
  LAYER VI3 ;
  RECT 320.240 5.940 320.440 6.140 ;
  LAYER VI3 ;
  RECT 319.840 6.340 320.040 6.540 ;
  LAYER VI3 ;
  RECT 319.840 5.940 320.040 6.140 ;
  LAYER VI3 ;
  RECT 319.440 6.340 319.640 6.540 ;
  LAYER VI3 ;
  RECT 319.440 5.940 319.640 6.140 ;
  LAYER VI3 ;
  RECT 319.040 6.340 319.240 6.540 ;
  LAYER VI3 ;
  RECT 319.040 5.940 319.240 6.140 ;
  LAYER VI3 ;
  RECT 318.640 6.340 318.840 6.540 ;
  LAYER VI3 ;
  RECT 318.640 5.940 318.840 6.140 ;
  LAYER VI3 ;
  RECT 318.240 6.340 318.440 6.540 ;
  LAYER VI3 ;
  RECT 318.240 5.940 318.440 6.140 ;
  LAYER VI3 ;
  RECT 317.840 6.340 318.040 6.540 ;
  LAYER VI3 ;
  RECT 317.840 5.940 318.040 6.140 ;
  LAYER VI3 ;
  RECT 317.440 6.340 317.640 6.540 ;
  LAYER VI3 ;
  RECT 317.440 5.940 317.640 6.140 ;
  LAYER VI3 ;
  RECT 317.040 6.340 317.240 6.540 ;
  LAYER VI3 ;
  RECT 317.040 5.940 317.240 6.140 ;
  LAYER VI3 ;
  RECT 316.640 6.340 316.840 6.540 ;
  LAYER VI3 ;
  RECT 316.640 5.940 316.840 6.140 ;
  LAYER VI3 ;
  RECT 316.240 6.340 316.440 6.540 ;
  LAYER VI3 ;
  RECT 316.240 5.940 316.440 6.140 ;
  LAYER VI3 ;
  RECT 315.840 6.340 316.040 6.540 ;
  LAYER VI3 ;
  RECT 315.840 5.940 316.040 6.140 ;
  LAYER VI3 ;
  RECT 315.440 6.340 315.640 6.540 ;
  LAYER VI3 ;
  RECT 315.440 5.940 315.640 6.140 ;
  LAYER VI3 ;
  RECT 315.040 6.340 315.240 6.540 ;
  LAYER VI3 ;
  RECT 315.040 5.940 315.240 6.140 ;
  LAYER VI3 ;
  RECT 314.640 6.340 314.840 6.540 ;
  LAYER VI3 ;
  RECT 314.640 5.940 314.840 6.140 ;
  LAYER VI3 ;
  RECT 335.720 5.880 343.720 6.740 ;
  LAYER VI3 ;
  RECT 343.320 6.340 343.520 6.540 ;
  LAYER VI3 ;
  RECT 343.320 5.940 343.520 6.140 ;
  LAYER VI3 ;
  RECT 342.920 6.340 343.120 6.540 ;
  LAYER VI3 ;
  RECT 342.920 5.940 343.120 6.140 ;
  LAYER VI3 ;
  RECT 342.520 6.340 342.720 6.540 ;
  LAYER VI3 ;
  RECT 342.520 5.940 342.720 6.140 ;
  LAYER VI3 ;
  RECT 342.120 6.340 342.320 6.540 ;
  LAYER VI3 ;
  RECT 342.120 5.940 342.320 6.140 ;
  LAYER VI3 ;
  RECT 341.720 6.340 341.920 6.540 ;
  LAYER VI3 ;
  RECT 341.720 5.940 341.920 6.140 ;
  LAYER VI3 ;
  RECT 341.320 6.340 341.520 6.540 ;
  LAYER VI3 ;
  RECT 341.320 5.940 341.520 6.140 ;
  LAYER VI3 ;
  RECT 340.920 6.340 341.120 6.540 ;
  LAYER VI3 ;
  RECT 340.920 5.940 341.120 6.140 ;
  LAYER VI3 ;
  RECT 340.520 6.340 340.720 6.540 ;
  LAYER VI3 ;
  RECT 340.520 5.940 340.720 6.140 ;
  LAYER VI3 ;
  RECT 340.120 6.340 340.320 6.540 ;
  LAYER VI3 ;
  RECT 340.120 5.940 340.320 6.140 ;
  LAYER VI3 ;
  RECT 339.720 6.340 339.920 6.540 ;
  LAYER VI3 ;
  RECT 339.720 5.940 339.920 6.140 ;
  LAYER VI3 ;
  RECT 339.320 6.340 339.520 6.540 ;
  LAYER VI3 ;
  RECT 339.320 5.940 339.520 6.140 ;
  LAYER VI3 ;
  RECT 338.920 6.340 339.120 6.540 ;
  LAYER VI3 ;
  RECT 338.920 5.940 339.120 6.140 ;
  LAYER VI3 ;
  RECT 338.520 6.340 338.720 6.540 ;
  LAYER VI3 ;
  RECT 338.520 5.940 338.720 6.140 ;
  LAYER VI3 ;
  RECT 338.120 6.340 338.320 6.540 ;
  LAYER VI3 ;
  RECT 338.120 5.940 338.320 6.140 ;
  LAYER VI3 ;
  RECT 337.720 6.340 337.920 6.540 ;
  LAYER VI3 ;
  RECT 337.720 5.940 337.920 6.140 ;
  LAYER VI3 ;
  RECT 337.320 6.340 337.520 6.540 ;
  LAYER VI3 ;
  RECT 337.320 5.940 337.520 6.140 ;
  LAYER VI3 ;
  RECT 336.920 6.340 337.120 6.540 ;
  LAYER VI3 ;
  RECT 336.920 5.940 337.120 6.140 ;
  LAYER VI3 ;
  RECT 336.520 6.340 336.720 6.540 ;
  LAYER VI3 ;
  RECT 336.520 5.940 336.720 6.140 ;
  LAYER VI3 ;
  RECT 336.120 6.340 336.320 6.540 ;
  LAYER VI3 ;
  RECT 336.120 5.940 336.320 6.140 ;
  LAYER VI3 ;
  RECT 335.720 6.340 335.920 6.540 ;
  LAYER VI3 ;
  RECT 335.720 5.940 335.920 6.140 ;
  LAYER VI3 ;
  RECT 355.560 5.880 363.560 6.740 ;
  LAYER VI3 ;
  RECT 363.160 6.340 363.360 6.540 ;
  LAYER VI3 ;
  RECT 363.160 5.940 363.360 6.140 ;
  LAYER VI3 ;
  RECT 362.760 6.340 362.960 6.540 ;
  LAYER VI3 ;
  RECT 362.760 5.940 362.960 6.140 ;
  LAYER VI3 ;
  RECT 362.360 6.340 362.560 6.540 ;
  LAYER VI3 ;
  RECT 362.360 5.940 362.560 6.140 ;
  LAYER VI3 ;
  RECT 361.960 6.340 362.160 6.540 ;
  LAYER VI3 ;
  RECT 361.960 5.940 362.160 6.140 ;
  LAYER VI3 ;
  RECT 361.560 6.340 361.760 6.540 ;
  LAYER VI3 ;
  RECT 361.560 5.940 361.760 6.140 ;
  LAYER VI3 ;
  RECT 361.160 6.340 361.360 6.540 ;
  LAYER VI3 ;
  RECT 361.160 5.940 361.360 6.140 ;
  LAYER VI3 ;
  RECT 360.760 6.340 360.960 6.540 ;
  LAYER VI3 ;
  RECT 360.760 5.940 360.960 6.140 ;
  LAYER VI3 ;
  RECT 360.360 6.340 360.560 6.540 ;
  LAYER VI3 ;
  RECT 360.360 5.940 360.560 6.140 ;
  LAYER VI3 ;
  RECT 359.960 6.340 360.160 6.540 ;
  LAYER VI3 ;
  RECT 359.960 5.940 360.160 6.140 ;
  LAYER VI3 ;
  RECT 359.560 6.340 359.760 6.540 ;
  LAYER VI3 ;
  RECT 359.560 5.940 359.760 6.140 ;
  LAYER VI3 ;
  RECT 359.160 6.340 359.360 6.540 ;
  LAYER VI3 ;
  RECT 359.160 5.940 359.360 6.140 ;
  LAYER VI3 ;
  RECT 358.760 6.340 358.960 6.540 ;
  LAYER VI3 ;
  RECT 358.760 5.940 358.960 6.140 ;
  LAYER VI3 ;
  RECT 358.360 6.340 358.560 6.540 ;
  LAYER VI3 ;
  RECT 358.360 5.940 358.560 6.140 ;
  LAYER VI3 ;
  RECT 357.960 6.340 358.160 6.540 ;
  LAYER VI3 ;
  RECT 357.960 5.940 358.160 6.140 ;
  LAYER VI3 ;
  RECT 357.560 6.340 357.760 6.540 ;
  LAYER VI3 ;
  RECT 357.560 5.940 357.760 6.140 ;
  LAYER VI3 ;
  RECT 357.160 6.340 357.360 6.540 ;
  LAYER VI3 ;
  RECT 357.160 5.940 357.360 6.140 ;
  LAYER VI3 ;
  RECT 356.760 6.340 356.960 6.540 ;
  LAYER VI3 ;
  RECT 356.760 5.940 356.960 6.140 ;
  LAYER VI3 ;
  RECT 356.360 6.340 356.560 6.540 ;
  LAYER VI3 ;
  RECT 356.360 5.940 356.560 6.140 ;
  LAYER VI3 ;
  RECT 355.960 6.340 356.160 6.540 ;
  LAYER VI3 ;
  RECT 355.960 5.940 356.160 6.140 ;
  LAYER VI3 ;
  RECT 355.560 6.340 355.760 6.540 ;
  LAYER VI3 ;
  RECT 355.560 5.940 355.760 6.140 ;
  LAYER VI3 ;
  RECT 376.640 5.880 384.640 6.740 ;
  LAYER VI3 ;
  RECT 384.240 6.340 384.440 6.540 ;
  LAYER VI3 ;
  RECT 384.240 5.940 384.440 6.140 ;
  LAYER VI3 ;
  RECT 383.840 6.340 384.040 6.540 ;
  LAYER VI3 ;
  RECT 383.840 5.940 384.040 6.140 ;
  LAYER VI3 ;
  RECT 383.440 6.340 383.640 6.540 ;
  LAYER VI3 ;
  RECT 383.440 5.940 383.640 6.140 ;
  LAYER VI3 ;
  RECT 383.040 6.340 383.240 6.540 ;
  LAYER VI3 ;
  RECT 383.040 5.940 383.240 6.140 ;
  LAYER VI3 ;
  RECT 382.640 6.340 382.840 6.540 ;
  LAYER VI3 ;
  RECT 382.640 5.940 382.840 6.140 ;
  LAYER VI3 ;
  RECT 382.240 6.340 382.440 6.540 ;
  LAYER VI3 ;
  RECT 382.240 5.940 382.440 6.140 ;
  LAYER VI3 ;
  RECT 381.840 6.340 382.040 6.540 ;
  LAYER VI3 ;
  RECT 381.840 5.940 382.040 6.140 ;
  LAYER VI3 ;
  RECT 381.440 6.340 381.640 6.540 ;
  LAYER VI3 ;
  RECT 381.440 5.940 381.640 6.140 ;
  LAYER VI3 ;
  RECT 381.040 6.340 381.240 6.540 ;
  LAYER VI3 ;
  RECT 381.040 5.940 381.240 6.140 ;
  LAYER VI3 ;
  RECT 380.640 6.340 380.840 6.540 ;
  LAYER VI3 ;
  RECT 380.640 5.940 380.840 6.140 ;
  LAYER VI3 ;
  RECT 380.240 6.340 380.440 6.540 ;
  LAYER VI3 ;
  RECT 380.240 5.940 380.440 6.140 ;
  LAYER VI3 ;
  RECT 379.840 6.340 380.040 6.540 ;
  LAYER VI3 ;
  RECT 379.840 5.940 380.040 6.140 ;
  LAYER VI3 ;
  RECT 379.440 6.340 379.640 6.540 ;
  LAYER VI3 ;
  RECT 379.440 5.940 379.640 6.140 ;
  LAYER VI3 ;
  RECT 379.040 6.340 379.240 6.540 ;
  LAYER VI3 ;
  RECT 379.040 5.940 379.240 6.140 ;
  LAYER VI3 ;
  RECT 378.640 6.340 378.840 6.540 ;
  LAYER VI3 ;
  RECT 378.640 5.940 378.840 6.140 ;
  LAYER VI3 ;
  RECT 378.240 6.340 378.440 6.540 ;
  LAYER VI3 ;
  RECT 378.240 5.940 378.440 6.140 ;
  LAYER VI3 ;
  RECT 377.840 6.340 378.040 6.540 ;
  LAYER VI3 ;
  RECT 377.840 5.940 378.040 6.140 ;
  LAYER VI3 ;
  RECT 377.440 6.340 377.640 6.540 ;
  LAYER VI3 ;
  RECT 377.440 5.940 377.640 6.140 ;
  LAYER VI3 ;
  RECT 377.040 6.340 377.240 6.540 ;
  LAYER VI3 ;
  RECT 377.040 5.940 377.240 6.140 ;
  LAYER VI3 ;
  RECT 376.640 6.340 376.840 6.540 ;
  LAYER VI3 ;
  RECT 376.640 5.940 376.840 6.140 ;
  LAYER VI3 ;
  RECT 396.480 5.880 404.480 6.740 ;
  LAYER VI3 ;
  RECT 404.080 6.340 404.280 6.540 ;
  LAYER VI3 ;
  RECT 404.080 5.940 404.280 6.140 ;
  LAYER VI3 ;
  RECT 403.680 6.340 403.880 6.540 ;
  LAYER VI3 ;
  RECT 403.680 5.940 403.880 6.140 ;
  LAYER VI3 ;
  RECT 403.280 6.340 403.480 6.540 ;
  LAYER VI3 ;
  RECT 403.280 5.940 403.480 6.140 ;
  LAYER VI3 ;
  RECT 402.880 6.340 403.080 6.540 ;
  LAYER VI3 ;
  RECT 402.880 5.940 403.080 6.140 ;
  LAYER VI3 ;
  RECT 402.480 6.340 402.680 6.540 ;
  LAYER VI3 ;
  RECT 402.480 5.940 402.680 6.140 ;
  LAYER VI3 ;
  RECT 402.080 6.340 402.280 6.540 ;
  LAYER VI3 ;
  RECT 402.080 5.940 402.280 6.140 ;
  LAYER VI3 ;
  RECT 401.680 6.340 401.880 6.540 ;
  LAYER VI3 ;
  RECT 401.680 5.940 401.880 6.140 ;
  LAYER VI3 ;
  RECT 401.280 6.340 401.480 6.540 ;
  LAYER VI3 ;
  RECT 401.280 5.940 401.480 6.140 ;
  LAYER VI3 ;
  RECT 400.880 6.340 401.080 6.540 ;
  LAYER VI3 ;
  RECT 400.880 5.940 401.080 6.140 ;
  LAYER VI3 ;
  RECT 400.480 6.340 400.680 6.540 ;
  LAYER VI3 ;
  RECT 400.480 5.940 400.680 6.140 ;
  LAYER VI3 ;
  RECT 400.080 6.340 400.280 6.540 ;
  LAYER VI3 ;
  RECT 400.080 5.940 400.280 6.140 ;
  LAYER VI3 ;
  RECT 399.680 6.340 399.880 6.540 ;
  LAYER VI3 ;
  RECT 399.680 5.940 399.880 6.140 ;
  LAYER VI3 ;
  RECT 399.280 6.340 399.480 6.540 ;
  LAYER VI3 ;
  RECT 399.280 5.940 399.480 6.140 ;
  LAYER VI3 ;
  RECT 398.880 6.340 399.080 6.540 ;
  LAYER VI3 ;
  RECT 398.880 5.940 399.080 6.140 ;
  LAYER VI3 ;
  RECT 398.480 6.340 398.680 6.540 ;
  LAYER VI3 ;
  RECT 398.480 5.940 398.680 6.140 ;
  LAYER VI3 ;
  RECT 398.080 6.340 398.280 6.540 ;
  LAYER VI3 ;
  RECT 398.080 5.940 398.280 6.140 ;
  LAYER VI3 ;
  RECT 397.680 6.340 397.880 6.540 ;
  LAYER VI3 ;
  RECT 397.680 5.940 397.880 6.140 ;
  LAYER VI3 ;
  RECT 397.280 6.340 397.480 6.540 ;
  LAYER VI3 ;
  RECT 397.280 5.940 397.480 6.140 ;
  LAYER VI3 ;
  RECT 396.880 6.340 397.080 6.540 ;
  LAYER VI3 ;
  RECT 396.880 5.940 397.080 6.140 ;
  LAYER VI3 ;
  RECT 396.480 6.340 396.680 6.540 ;
  LAYER VI3 ;
  RECT 396.480 5.940 396.680 6.140 ;
  LAYER VI3 ;
  RECT 417.560 5.880 425.560 6.740 ;
  LAYER VI3 ;
  RECT 425.160 6.340 425.360 6.540 ;
  LAYER VI3 ;
  RECT 425.160 5.940 425.360 6.140 ;
  LAYER VI3 ;
  RECT 424.760 6.340 424.960 6.540 ;
  LAYER VI3 ;
  RECT 424.760 5.940 424.960 6.140 ;
  LAYER VI3 ;
  RECT 424.360 6.340 424.560 6.540 ;
  LAYER VI3 ;
  RECT 424.360 5.940 424.560 6.140 ;
  LAYER VI3 ;
  RECT 423.960 6.340 424.160 6.540 ;
  LAYER VI3 ;
  RECT 423.960 5.940 424.160 6.140 ;
  LAYER VI3 ;
  RECT 423.560 6.340 423.760 6.540 ;
  LAYER VI3 ;
  RECT 423.560 5.940 423.760 6.140 ;
  LAYER VI3 ;
  RECT 423.160 6.340 423.360 6.540 ;
  LAYER VI3 ;
  RECT 423.160 5.940 423.360 6.140 ;
  LAYER VI3 ;
  RECT 422.760 6.340 422.960 6.540 ;
  LAYER VI3 ;
  RECT 422.760 5.940 422.960 6.140 ;
  LAYER VI3 ;
  RECT 422.360 6.340 422.560 6.540 ;
  LAYER VI3 ;
  RECT 422.360 5.940 422.560 6.140 ;
  LAYER VI3 ;
  RECT 421.960 6.340 422.160 6.540 ;
  LAYER VI3 ;
  RECT 421.960 5.940 422.160 6.140 ;
  LAYER VI3 ;
  RECT 421.560 6.340 421.760 6.540 ;
  LAYER VI3 ;
  RECT 421.560 5.940 421.760 6.140 ;
  LAYER VI3 ;
  RECT 421.160 6.340 421.360 6.540 ;
  LAYER VI3 ;
  RECT 421.160 5.940 421.360 6.140 ;
  LAYER VI3 ;
  RECT 420.760 6.340 420.960 6.540 ;
  LAYER VI3 ;
  RECT 420.760 5.940 420.960 6.140 ;
  LAYER VI3 ;
  RECT 420.360 6.340 420.560 6.540 ;
  LAYER VI3 ;
  RECT 420.360 5.940 420.560 6.140 ;
  LAYER VI3 ;
  RECT 419.960 6.340 420.160 6.540 ;
  LAYER VI3 ;
  RECT 419.960 5.940 420.160 6.140 ;
  LAYER VI3 ;
  RECT 419.560 6.340 419.760 6.540 ;
  LAYER VI3 ;
  RECT 419.560 5.940 419.760 6.140 ;
  LAYER VI3 ;
  RECT 419.160 6.340 419.360 6.540 ;
  LAYER VI3 ;
  RECT 419.160 5.940 419.360 6.140 ;
  LAYER VI3 ;
  RECT 418.760 6.340 418.960 6.540 ;
  LAYER VI3 ;
  RECT 418.760 5.940 418.960 6.140 ;
  LAYER VI3 ;
  RECT 418.360 6.340 418.560 6.540 ;
  LAYER VI3 ;
  RECT 418.360 5.940 418.560 6.140 ;
  LAYER VI3 ;
  RECT 417.960 6.340 418.160 6.540 ;
  LAYER VI3 ;
  RECT 417.960 5.940 418.160 6.140 ;
  LAYER VI3 ;
  RECT 417.560 6.340 417.760 6.540 ;
  LAYER VI3 ;
  RECT 417.560 5.940 417.760 6.140 ;
  LAYER VI3 ;
  RECT 437.400 5.880 445.400 6.740 ;
  LAYER VI3 ;
  RECT 445.000 6.340 445.200 6.540 ;
  LAYER VI3 ;
  RECT 445.000 5.940 445.200 6.140 ;
  LAYER VI3 ;
  RECT 444.600 6.340 444.800 6.540 ;
  LAYER VI3 ;
  RECT 444.600 5.940 444.800 6.140 ;
  LAYER VI3 ;
  RECT 444.200 6.340 444.400 6.540 ;
  LAYER VI3 ;
  RECT 444.200 5.940 444.400 6.140 ;
  LAYER VI3 ;
  RECT 443.800 6.340 444.000 6.540 ;
  LAYER VI3 ;
  RECT 443.800 5.940 444.000 6.140 ;
  LAYER VI3 ;
  RECT 443.400 6.340 443.600 6.540 ;
  LAYER VI3 ;
  RECT 443.400 5.940 443.600 6.140 ;
  LAYER VI3 ;
  RECT 443.000 6.340 443.200 6.540 ;
  LAYER VI3 ;
  RECT 443.000 5.940 443.200 6.140 ;
  LAYER VI3 ;
  RECT 442.600 6.340 442.800 6.540 ;
  LAYER VI3 ;
  RECT 442.600 5.940 442.800 6.140 ;
  LAYER VI3 ;
  RECT 442.200 6.340 442.400 6.540 ;
  LAYER VI3 ;
  RECT 442.200 5.940 442.400 6.140 ;
  LAYER VI3 ;
  RECT 441.800 6.340 442.000 6.540 ;
  LAYER VI3 ;
  RECT 441.800 5.940 442.000 6.140 ;
  LAYER VI3 ;
  RECT 441.400 6.340 441.600 6.540 ;
  LAYER VI3 ;
  RECT 441.400 5.940 441.600 6.140 ;
  LAYER VI3 ;
  RECT 441.000 6.340 441.200 6.540 ;
  LAYER VI3 ;
  RECT 441.000 5.940 441.200 6.140 ;
  LAYER VI3 ;
  RECT 440.600 6.340 440.800 6.540 ;
  LAYER VI3 ;
  RECT 440.600 5.940 440.800 6.140 ;
  LAYER VI3 ;
  RECT 440.200 6.340 440.400 6.540 ;
  LAYER VI3 ;
  RECT 440.200 5.940 440.400 6.140 ;
  LAYER VI3 ;
  RECT 439.800 6.340 440.000 6.540 ;
  LAYER VI3 ;
  RECT 439.800 5.940 440.000 6.140 ;
  LAYER VI3 ;
  RECT 439.400 6.340 439.600 6.540 ;
  LAYER VI3 ;
  RECT 439.400 5.940 439.600 6.140 ;
  LAYER VI3 ;
  RECT 439.000 6.340 439.200 6.540 ;
  LAYER VI3 ;
  RECT 439.000 5.940 439.200 6.140 ;
  LAYER VI3 ;
  RECT 438.600 6.340 438.800 6.540 ;
  LAYER VI3 ;
  RECT 438.600 5.940 438.800 6.140 ;
  LAYER VI3 ;
  RECT 438.200 6.340 438.400 6.540 ;
  LAYER VI3 ;
  RECT 438.200 5.940 438.400 6.140 ;
  LAYER VI3 ;
  RECT 437.800 6.340 438.000 6.540 ;
  LAYER VI3 ;
  RECT 437.800 5.940 438.000 6.140 ;
  LAYER VI3 ;
  RECT 437.400 6.340 437.600 6.540 ;
  LAYER VI3 ;
  RECT 437.400 5.940 437.600 6.140 ;
  LAYER VI3 ;
  RECT 458.480 5.880 466.480 6.740 ;
  LAYER VI3 ;
  RECT 466.080 6.340 466.280 6.540 ;
  LAYER VI3 ;
  RECT 466.080 5.940 466.280 6.140 ;
  LAYER VI3 ;
  RECT 465.680 6.340 465.880 6.540 ;
  LAYER VI3 ;
  RECT 465.680 5.940 465.880 6.140 ;
  LAYER VI3 ;
  RECT 465.280 6.340 465.480 6.540 ;
  LAYER VI3 ;
  RECT 465.280 5.940 465.480 6.140 ;
  LAYER VI3 ;
  RECT 464.880 6.340 465.080 6.540 ;
  LAYER VI3 ;
  RECT 464.880 5.940 465.080 6.140 ;
  LAYER VI3 ;
  RECT 464.480 6.340 464.680 6.540 ;
  LAYER VI3 ;
  RECT 464.480 5.940 464.680 6.140 ;
  LAYER VI3 ;
  RECT 464.080 6.340 464.280 6.540 ;
  LAYER VI3 ;
  RECT 464.080 5.940 464.280 6.140 ;
  LAYER VI3 ;
  RECT 463.680 6.340 463.880 6.540 ;
  LAYER VI3 ;
  RECT 463.680 5.940 463.880 6.140 ;
  LAYER VI3 ;
  RECT 463.280 6.340 463.480 6.540 ;
  LAYER VI3 ;
  RECT 463.280 5.940 463.480 6.140 ;
  LAYER VI3 ;
  RECT 462.880 6.340 463.080 6.540 ;
  LAYER VI3 ;
  RECT 462.880 5.940 463.080 6.140 ;
  LAYER VI3 ;
  RECT 462.480 6.340 462.680 6.540 ;
  LAYER VI3 ;
  RECT 462.480 5.940 462.680 6.140 ;
  LAYER VI3 ;
  RECT 462.080 6.340 462.280 6.540 ;
  LAYER VI3 ;
  RECT 462.080 5.940 462.280 6.140 ;
  LAYER VI3 ;
  RECT 461.680 6.340 461.880 6.540 ;
  LAYER VI3 ;
  RECT 461.680 5.940 461.880 6.140 ;
  LAYER VI3 ;
  RECT 461.280 6.340 461.480 6.540 ;
  LAYER VI3 ;
  RECT 461.280 5.940 461.480 6.140 ;
  LAYER VI3 ;
  RECT 460.880 6.340 461.080 6.540 ;
  LAYER VI3 ;
  RECT 460.880 5.940 461.080 6.140 ;
  LAYER VI3 ;
  RECT 460.480 6.340 460.680 6.540 ;
  LAYER VI3 ;
  RECT 460.480 5.940 460.680 6.140 ;
  LAYER VI3 ;
  RECT 460.080 6.340 460.280 6.540 ;
  LAYER VI3 ;
  RECT 460.080 5.940 460.280 6.140 ;
  LAYER VI3 ;
  RECT 459.680 6.340 459.880 6.540 ;
  LAYER VI3 ;
  RECT 459.680 5.940 459.880 6.140 ;
  LAYER VI3 ;
  RECT 459.280 6.340 459.480 6.540 ;
  LAYER VI3 ;
  RECT 459.280 5.940 459.480 6.140 ;
  LAYER VI3 ;
  RECT 458.880 6.340 459.080 6.540 ;
  LAYER VI3 ;
  RECT 458.880 5.940 459.080 6.140 ;
  LAYER VI3 ;
  RECT 458.480 6.340 458.680 6.540 ;
  LAYER VI3 ;
  RECT 458.480 5.940 458.680 6.140 ;
  LAYER VI3 ;
  RECT 478.320 5.880 486.320 6.740 ;
  LAYER VI3 ;
  RECT 485.920 6.340 486.120 6.540 ;
  LAYER VI3 ;
  RECT 485.920 5.940 486.120 6.140 ;
  LAYER VI3 ;
  RECT 485.520 6.340 485.720 6.540 ;
  LAYER VI3 ;
  RECT 485.520 5.940 485.720 6.140 ;
  LAYER VI3 ;
  RECT 485.120 6.340 485.320 6.540 ;
  LAYER VI3 ;
  RECT 485.120 5.940 485.320 6.140 ;
  LAYER VI3 ;
  RECT 484.720 6.340 484.920 6.540 ;
  LAYER VI3 ;
  RECT 484.720 5.940 484.920 6.140 ;
  LAYER VI3 ;
  RECT 484.320 6.340 484.520 6.540 ;
  LAYER VI3 ;
  RECT 484.320 5.940 484.520 6.140 ;
  LAYER VI3 ;
  RECT 483.920 6.340 484.120 6.540 ;
  LAYER VI3 ;
  RECT 483.920 5.940 484.120 6.140 ;
  LAYER VI3 ;
  RECT 483.520 6.340 483.720 6.540 ;
  LAYER VI3 ;
  RECT 483.520 5.940 483.720 6.140 ;
  LAYER VI3 ;
  RECT 483.120 6.340 483.320 6.540 ;
  LAYER VI3 ;
  RECT 483.120 5.940 483.320 6.140 ;
  LAYER VI3 ;
  RECT 482.720 6.340 482.920 6.540 ;
  LAYER VI3 ;
  RECT 482.720 5.940 482.920 6.140 ;
  LAYER VI3 ;
  RECT 482.320 6.340 482.520 6.540 ;
  LAYER VI3 ;
  RECT 482.320 5.940 482.520 6.140 ;
  LAYER VI3 ;
  RECT 481.920 6.340 482.120 6.540 ;
  LAYER VI3 ;
  RECT 481.920 5.940 482.120 6.140 ;
  LAYER VI3 ;
  RECT 481.520 6.340 481.720 6.540 ;
  LAYER VI3 ;
  RECT 481.520 5.940 481.720 6.140 ;
  LAYER VI3 ;
  RECT 481.120 6.340 481.320 6.540 ;
  LAYER VI3 ;
  RECT 481.120 5.940 481.320 6.140 ;
  LAYER VI3 ;
  RECT 480.720 6.340 480.920 6.540 ;
  LAYER VI3 ;
  RECT 480.720 5.940 480.920 6.140 ;
  LAYER VI3 ;
  RECT 480.320 6.340 480.520 6.540 ;
  LAYER VI3 ;
  RECT 480.320 5.940 480.520 6.140 ;
  LAYER VI3 ;
  RECT 479.920 6.340 480.120 6.540 ;
  LAYER VI3 ;
  RECT 479.920 5.940 480.120 6.140 ;
  LAYER VI3 ;
  RECT 479.520 6.340 479.720 6.540 ;
  LAYER VI3 ;
  RECT 479.520 5.940 479.720 6.140 ;
  LAYER VI3 ;
  RECT 479.120 6.340 479.320 6.540 ;
  LAYER VI3 ;
  RECT 479.120 5.940 479.320 6.140 ;
  LAYER VI3 ;
  RECT 478.720 6.340 478.920 6.540 ;
  LAYER VI3 ;
  RECT 478.720 5.940 478.920 6.140 ;
  LAYER VI3 ;
  RECT 478.320 6.340 478.520 6.540 ;
  LAYER VI3 ;
  RECT 478.320 5.940 478.520 6.140 ;
  LAYER VI3 ;
  RECT 499.400 5.880 507.400 6.740 ;
  LAYER VI3 ;
  RECT 507.000 6.340 507.200 6.540 ;
  LAYER VI3 ;
  RECT 507.000 5.940 507.200 6.140 ;
  LAYER VI3 ;
  RECT 506.600 6.340 506.800 6.540 ;
  LAYER VI3 ;
  RECT 506.600 5.940 506.800 6.140 ;
  LAYER VI3 ;
  RECT 506.200 6.340 506.400 6.540 ;
  LAYER VI3 ;
  RECT 506.200 5.940 506.400 6.140 ;
  LAYER VI3 ;
  RECT 505.800 6.340 506.000 6.540 ;
  LAYER VI3 ;
  RECT 505.800 5.940 506.000 6.140 ;
  LAYER VI3 ;
  RECT 505.400 6.340 505.600 6.540 ;
  LAYER VI3 ;
  RECT 505.400 5.940 505.600 6.140 ;
  LAYER VI3 ;
  RECT 505.000 6.340 505.200 6.540 ;
  LAYER VI3 ;
  RECT 505.000 5.940 505.200 6.140 ;
  LAYER VI3 ;
  RECT 504.600 6.340 504.800 6.540 ;
  LAYER VI3 ;
  RECT 504.600 5.940 504.800 6.140 ;
  LAYER VI3 ;
  RECT 504.200 6.340 504.400 6.540 ;
  LAYER VI3 ;
  RECT 504.200 5.940 504.400 6.140 ;
  LAYER VI3 ;
  RECT 503.800 6.340 504.000 6.540 ;
  LAYER VI3 ;
  RECT 503.800 5.940 504.000 6.140 ;
  LAYER VI3 ;
  RECT 503.400 6.340 503.600 6.540 ;
  LAYER VI3 ;
  RECT 503.400 5.940 503.600 6.140 ;
  LAYER VI3 ;
  RECT 503.000 6.340 503.200 6.540 ;
  LAYER VI3 ;
  RECT 503.000 5.940 503.200 6.140 ;
  LAYER VI3 ;
  RECT 502.600 6.340 502.800 6.540 ;
  LAYER VI3 ;
  RECT 502.600 5.940 502.800 6.140 ;
  LAYER VI3 ;
  RECT 502.200 6.340 502.400 6.540 ;
  LAYER VI3 ;
  RECT 502.200 5.940 502.400 6.140 ;
  LAYER VI3 ;
  RECT 501.800 6.340 502.000 6.540 ;
  LAYER VI3 ;
  RECT 501.800 5.940 502.000 6.140 ;
  LAYER VI3 ;
  RECT 501.400 6.340 501.600 6.540 ;
  LAYER VI3 ;
  RECT 501.400 5.940 501.600 6.140 ;
  LAYER VI3 ;
  RECT 501.000 6.340 501.200 6.540 ;
  LAYER VI3 ;
  RECT 501.000 5.940 501.200 6.140 ;
  LAYER VI3 ;
  RECT 500.600 6.340 500.800 6.540 ;
  LAYER VI3 ;
  RECT 500.600 5.940 500.800 6.140 ;
  LAYER VI3 ;
  RECT 500.200 6.340 500.400 6.540 ;
  LAYER VI3 ;
  RECT 500.200 5.940 500.400 6.140 ;
  LAYER VI3 ;
  RECT 499.800 6.340 500.000 6.540 ;
  LAYER VI3 ;
  RECT 499.800 5.940 500.000 6.140 ;
  LAYER VI3 ;
  RECT 499.400 6.340 499.600 6.540 ;
  LAYER VI3 ;
  RECT 499.400 5.940 499.600 6.140 ;
  LAYER VI3 ;
  RECT 519.240 5.880 527.240 6.740 ;
  LAYER VI3 ;
  RECT 526.840 6.340 527.040 6.540 ;
  LAYER VI3 ;
  RECT 526.840 5.940 527.040 6.140 ;
  LAYER VI3 ;
  RECT 526.440 6.340 526.640 6.540 ;
  LAYER VI3 ;
  RECT 526.440 5.940 526.640 6.140 ;
  LAYER VI3 ;
  RECT 526.040 6.340 526.240 6.540 ;
  LAYER VI3 ;
  RECT 526.040 5.940 526.240 6.140 ;
  LAYER VI3 ;
  RECT 525.640 6.340 525.840 6.540 ;
  LAYER VI3 ;
  RECT 525.640 5.940 525.840 6.140 ;
  LAYER VI3 ;
  RECT 525.240 6.340 525.440 6.540 ;
  LAYER VI3 ;
  RECT 525.240 5.940 525.440 6.140 ;
  LAYER VI3 ;
  RECT 524.840 6.340 525.040 6.540 ;
  LAYER VI3 ;
  RECT 524.840 5.940 525.040 6.140 ;
  LAYER VI3 ;
  RECT 524.440 6.340 524.640 6.540 ;
  LAYER VI3 ;
  RECT 524.440 5.940 524.640 6.140 ;
  LAYER VI3 ;
  RECT 524.040 6.340 524.240 6.540 ;
  LAYER VI3 ;
  RECT 524.040 5.940 524.240 6.140 ;
  LAYER VI3 ;
  RECT 523.640 6.340 523.840 6.540 ;
  LAYER VI3 ;
  RECT 523.640 5.940 523.840 6.140 ;
  LAYER VI3 ;
  RECT 523.240 6.340 523.440 6.540 ;
  LAYER VI3 ;
  RECT 523.240 5.940 523.440 6.140 ;
  LAYER VI3 ;
  RECT 522.840 6.340 523.040 6.540 ;
  LAYER VI3 ;
  RECT 522.840 5.940 523.040 6.140 ;
  LAYER VI3 ;
  RECT 522.440 6.340 522.640 6.540 ;
  LAYER VI3 ;
  RECT 522.440 5.940 522.640 6.140 ;
  LAYER VI3 ;
  RECT 522.040 6.340 522.240 6.540 ;
  LAYER VI3 ;
  RECT 522.040 5.940 522.240 6.140 ;
  LAYER VI3 ;
  RECT 521.640 6.340 521.840 6.540 ;
  LAYER VI3 ;
  RECT 521.640 5.940 521.840 6.140 ;
  LAYER VI3 ;
  RECT 521.240 6.340 521.440 6.540 ;
  LAYER VI3 ;
  RECT 521.240 5.940 521.440 6.140 ;
  LAYER VI3 ;
  RECT 520.840 6.340 521.040 6.540 ;
  LAYER VI3 ;
  RECT 520.840 5.940 521.040 6.140 ;
  LAYER VI3 ;
  RECT 520.440 6.340 520.640 6.540 ;
  LAYER VI3 ;
  RECT 520.440 5.940 520.640 6.140 ;
  LAYER VI3 ;
  RECT 520.040 6.340 520.240 6.540 ;
  LAYER VI3 ;
  RECT 520.040 5.940 520.240 6.140 ;
  LAYER VI3 ;
  RECT 519.640 6.340 519.840 6.540 ;
  LAYER VI3 ;
  RECT 519.640 5.940 519.840 6.140 ;
  LAYER VI3 ;
  RECT 519.240 6.340 519.440 6.540 ;
  LAYER VI3 ;
  RECT 519.240 5.940 519.440 6.140 ;
  LAYER VI3 ;
  RECT 540.320 5.880 548.320 6.740 ;
  LAYER VI3 ;
  RECT 547.920 6.340 548.120 6.540 ;
  LAYER VI3 ;
  RECT 547.920 5.940 548.120 6.140 ;
  LAYER VI3 ;
  RECT 547.520 6.340 547.720 6.540 ;
  LAYER VI3 ;
  RECT 547.520 5.940 547.720 6.140 ;
  LAYER VI3 ;
  RECT 547.120 6.340 547.320 6.540 ;
  LAYER VI3 ;
  RECT 547.120 5.940 547.320 6.140 ;
  LAYER VI3 ;
  RECT 546.720 6.340 546.920 6.540 ;
  LAYER VI3 ;
  RECT 546.720 5.940 546.920 6.140 ;
  LAYER VI3 ;
  RECT 546.320 6.340 546.520 6.540 ;
  LAYER VI3 ;
  RECT 546.320 5.940 546.520 6.140 ;
  LAYER VI3 ;
  RECT 545.920 6.340 546.120 6.540 ;
  LAYER VI3 ;
  RECT 545.920 5.940 546.120 6.140 ;
  LAYER VI3 ;
  RECT 545.520 6.340 545.720 6.540 ;
  LAYER VI3 ;
  RECT 545.520 5.940 545.720 6.140 ;
  LAYER VI3 ;
  RECT 545.120 6.340 545.320 6.540 ;
  LAYER VI3 ;
  RECT 545.120 5.940 545.320 6.140 ;
  LAYER VI3 ;
  RECT 544.720 6.340 544.920 6.540 ;
  LAYER VI3 ;
  RECT 544.720 5.940 544.920 6.140 ;
  LAYER VI3 ;
  RECT 544.320 6.340 544.520 6.540 ;
  LAYER VI3 ;
  RECT 544.320 5.940 544.520 6.140 ;
  LAYER VI3 ;
  RECT 543.920 6.340 544.120 6.540 ;
  LAYER VI3 ;
  RECT 543.920 5.940 544.120 6.140 ;
  LAYER VI3 ;
  RECT 543.520 6.340 543.720 6.540 ;
  LAYER VI3 ;
  RECT 543.520 5.940 543.720 6.140 ;
  LAYER VI3 ;
  RECT 543.120 6.340 543.320 6.540 ;
  LAYER VI3 ;
  RECT 543.120 5.940 543.320 6.140 ;
  LAYER VI3 ;
  RECT 542.720 6.340 542.920 6.540 ;
  LAYER VI3 ;
  RECT 542.720 5.940 542.920 6.140 ;
  LAYER VI3 ;
  RECT 542.320 6.340 542.520 6.540 ;
  LAYER VI3 ;
  RECT 542.320 5.940 542.520 6.140 ;
  LAYER VI3 ;
  RECT 541.920 6.340 542.120 6.540 ;
  LAYER VI3 ;
  RECT 541.920 5.940 542.120 6.140 ;
  LAYER VI3 ;
  RECT 541.520 6.340 541.720 6.540 ;
  LAYER VI3 ;
  RECT 541.520 5.940 541.720 6.140 ;
  LAYER VI3 ;
  RECT 541.120 6.340 541.320 6.540 ;
  LAYER VI3 ;
  RECT 541.120 5.940 541.320 6.140 ;
  LAYER VI3 ;
  RECT 540.720 6.340 540.920 6.540 ;
  LAYER VI3 ;
  RECT 540.720 5.940 540.920 6.140 ;
  LAYER VI3 ;
  RECT 540.320 6.340 540.520 6.540 ;
  LAYER VI3 ;
  RECT 540.320 5.940 540.520 6.140 ;
  LAYER VI3 ;
  RECT 560.160 5.880 568.160 6.740 ;
  LAYER VI3 ;
  RECT 567.760 6.340 567.960 6.540 ;
  LAYER VI3 ;
  RECT 567.760 5.940 567.960 6.140 ;
  LAYER VI3 ;
  RECT 567.360 6.340 567.560 6.540 ;
  LAYER VI3 ;
  RECT 567.360 5.940 567.560 6.140 ;
  LAYER VI3 ;
  RECT 566.960 6.340 567.160 6.540 ;
  LAYER VI3 ;
  RECT 566.960 5.940 567.160 6.140 ;
  LAYER VI3 ;
  RECT 566.560 6.340 566.760 6.540 ;
  LAYER VI3 ;
  RECT 566.560 5.940 566.760 6.140 ;
  LAYER VI3 ;
  RECT 566.160 6.340 566.360 6.540 ;
  LAYER VI3 ;
  RECT 566.160 5.940 566.360 6.140 ;
  LAYER VI3 ;
  RECT 565.760 6.340 565.960 6.540 ;
  LAYER VI3 ;
  RECT 565.760 5.940 565.960 6.140 ;
  LAYER VI3 ;
  RECT 565.360 6.340 565.560 6.540 ;
  LAYER VI3 ;
  RECT 565.360 5.940 565.560 6.140 ;
  LAYER VI3 ;
  RECT 564.960 6.340 565.160 6.540 ;
  LAYER VI3 ;
  RECT 564.960 5.940 565.160 6.140 ;
  LAYER VI3 ;
  RECT 564.560 6.340 564.760 6.540 ;
  LAYER VI3 ;
  RECT 564.560 5.940 564.760 6.140 ;
  LAYER VI3 ;
  RECT 564.160 6.340 564.360 6.540 ;
  LAYER VI3 ;
  RECT 564.160 5.940 564.360 6.140 ;
  LAYER VI3 ;
  RECT 563.760 6.340 563.960 6.540 ;
  LAYER VI3 ;
  RECT 563.760 5.940 563.960 6.140 ;
  LAYER VI3 ;
  RECT 563.360 6.340 563.560 6.540 ;
  LAYER VI3 ;
  RECT 563.360 5.940 563.560 6.140 ;
  LAYER VI3 ;
  RECT 562.960 6.340 563.160 6.540 ;
  LAYER VI3 ;
  RECT 562.960 5.940 563.160 6.140 ;
  LAYER VI3 ;
  RECT 562.560 6.340 562.760 6.540 ;
  LAYER VI3 ;
  RECT 562.560 5.940 562.760 6.140 ;
  LAYER VI3 ;
  RECT 562.160 6.340 562.360 6.540 ;
  LAYER VI3 ;
  RECT 562.160 5.940 562.360 6.140 ;
  LAYER VI3 ;
  RECT 561.760 6.340 561.960 6.540 ;
  LAYER VI3 ;
  RECT 561.760 5.940 561.960 6.140 ;
  LAYER VI3 ;
  RECT 561.360 6.340 561.560 6.540 ;
  LAYER VI3 ;
  RECT 561.360 5.940 561.560 6.140 ;
  LAYER VI3 ;
  RECT 560.960 6.340 561.160 6.540 ;
  LAYER VI3 ;
  RECT 560.960 5.940 561.160 6.140 ;
  LAYER VI3 ;
  RECT 560.560 6.340 560.760 6.540 ;
  LAYER VI3 ;
  RECT 560.560 5.940 560.760 6.140 ;
  LAYER VI3 ;
  RECT 560.160 6.340 560.360 6.540 ;
  LAYER VI3 ;
  RECT 560.160 5.940 560.360 6.140 ;
  LAYER VI3 ;
  RECT 581.240 5.880 589.240 6.740 ;
  LAYER VI3 ;
  RECT 588.840 6.340 589.040 6.540 ;
  LAYER VI3 ;
  RECT 588.840 5.940 589.040 6.140 ;
  LAYER VI3 ;
  RECT 588.440 6.340 588.640 6.540 ;
  LAYER VI3 ;
  RECT 588.440 5.940 588.640 6.140 ;
  LAYER VI3 ;
  RECT 588.040 6.340 588.240 6.540 ;
  LAYER VI3 ;
  RECT 588.040 5.940 588.240 6.140 ;
  LAYER VI3 ;
  RECT 587.640 6.340 587.840 6.540 ;
  LAYER VI3 ;
  RECT 587.640 5.940 587.840 6.140 ;
  LAYER VI3 ;
  RECT 587.240 6.340 587.440 6.540 ;
  LAYER VI3 ;
  RECT 587.240 5.940 587.440 6.140 ;
  LAYER VI3 ;
  RECT 586.840 6.340 587.040 6.540 ;
  LAYER VI3 ;
  RECT 586.840 5.940 587.040 6.140 ;
  LAYER VI3 ;
  RECT 586.440 6.340 586.640 6.540 ;
  LAYER VI3 ;
  RECT 586.440 5.940 586.640 6.140 ;
  LAYER VI3 ;
  RECT 586.040 6.340 586.240 6.540 ;
  LAYER VI3 ;
  RECT 586.040 5.940 586.240 6.140 ;
  LAYER VI3 ;
  RECT 585.640 6.340 585.840 6.540 ;
  LAYER VI3 ;
  RECT 585.640 5.940 585.840 6.140 ;
  LAYER VI3 ;
  RECT 585.240 6.340 585.440 6.540 ;
  LAYER VI3 ;
  RECT 585.240 5.940 585.440 6.140 ;
  LAYER VI3 ;
  RECT 584.840 6.340 585.040 6.540 ;
  LAYER VI3 ;
  RECT 584.840 5.940 585.040 6.140 ;
  LAYER VI3 ;
  RECT 584.440 6.340 584.640 6.540 ;
  LAYER VI3 ;
  RECT 584.440 5.940 584.640 6.140 ;
  LAYER VI3 ;
  RECT 584.040 6.340 584.240 6.540 ;
  LAYER VI3 ;
  RECT 584.040 5.940 584.240 6.140 ;
  LAYER VI3 ;
  RECT 583.640 6.340 583.840 6.540 ;
  LAYER VI3 ;
  RECT 583.640 5.940 583.840 6.140 ;
  LAYER VI3 ;
  RECT 583.240 6.340 583.440 6.540 ;
  LAYER VI3 ;
  RECT 583.240 5.940 583.440 6.140 ;
  LAYER VI3 ;
  RECT 582.840 6.340 583.040 6.540 ;
  LAYER VI3 ;
  RECT 582.840 5.940 583.040 6.140 ;
  LAYER VI3 ;
  RECT 582.440 6.340 582.640 6.540 ;
  LAYER VI3 ;
  RECT 582.440 5.940 582.640 6.140 ;
  LAYER VI3 ;
  RECT 582.040 6.340 582.240 6.540 ;
  LAYER VI3 ;
  RECT 582.040 5.940 582.240 6.140 ;
  LAYER VI3 ;
  RECT 581.640 6.340 581.840 6.540 ;
  LAYER VI3 ;
  RECT 581.640 5.940 581.840 6.140 ;
  LAYER VI3 ;
  RECT 581.240 6.340 581.440 6.540 ;
  LAYER VI3 ;
  RECT 581.240 5.940 581.440 6.140 ;
  LAYER VI3 ;
  RECT 601.080 5.880 609.080 6.740 ;
  LAYER VI3 ;
  RECT 608.680 6.340 608.880 6.540 ;
  LAYER VI3 ;
  RECT 608.680 5.940 608.880 6.140 ;
  LAYER VI3 ;
  RECT 608.280 6.340 608.480 6.540 ;
  LAYER VI3 ;
  RECT 608.280 5.940 608.480 6.140 ;
  LAYER VI3 ;
  RECT 607.880 6.340 608.080 6.540 ;
  LAYER VI3 ;
  RECT 607.880 5.940 608.080 6.140 ;
  LAYER VI3 ;
  RECT 607.480 6.340 607.680 6.540 ;
  LAYER VI3 ;
  RECT 607.480 5.940 607.680 6.140 ;
  LAYER VI3 ;
  RECT 607.080 6.340 607.280 6.540 ;
  LAYER VI3 ;
  RECT 607.080 5.940 607.280 6.140 ;
  LAYER VI3 ;
  RECT 606.680 6.340 606.880 6.540 ;
  LAYER VI3 ;
  RECT 606.680 5.940 606.880 6.140 ;
  LAYER VI3 ;
  RECT 606.280 6.340 606.480 6.540 ;
  LAYER VI3 ;
  RECT 606.280 5.940 606.480 6.140 ;
  LAYER VI3 ;
  RECT 605.880 6.340 606.080 6.540 ;
  LAYER VI3 ;
  RECT 605.880 5.940 606.080 6.140 ;
  LAYER VI3 ;
  RECT 605.480 6.340 605.680 6.540 ;
  LAYER VI3 ;
  RECT 605.480 5.940 605.680 6.140 ;
  LAYER VI3 ;
  RECT 605.080 6.340 605.280 6.540 ;
  LAYER VI3 ;
  RECT 605.080 5.940 605.280 6.140 ;
  LAYER VI3 ;
  RECT 604.680 6.340 604.880 6.540 ;
  LAYER VI3 ;
  RECT 604.680 5.940 604.880 6.140 ;
  LAYER VI3 ;
  RECT 604.280 6.340 604.480 6.540 ;
  LAYER VI3 ;
  RECT 604.280 5.940 604.480 6.140 ;
  LAYER VI3 ;
  RECT 603.880 6.340 604.080 6.540 ;
  LAYER VI3 ;
  RECT 603.880 5.940 604.080 6.140 ;
  LAYER VI3 ;
  RECT 603.480 6.340 603.680 6.540 ;
  LAYER VI3 ;
  RECT 603.480 5.940 603.680 6.140 ;
  LAYER VI3 ;
  RECT 603.080 6.340 603.280 6.540 ;
  LAYER VI3 ;
  RECT 603.080 5.940 603.280 6.140 ;
  LAYER VI3 ;
  RECT 602.680 6.340 602.880 6.540 ;
  LAYER VI3 ;
  RECT 602.680 5.940 602.880 6.140 ;
  LAYER VI3 ;
  RECT 602.280 6.340 602.480 6.540 ;
  LAYER VI3 ;
  RECT 602.280 5.940 602.480 6.140 ;
  LAYER VI3 ;
  RECT 601.880 6.340 602.080 6.540 ;
  LAYER VI3 ;
  RECT 601.880 5.940 602.080 6.140 ;
  LAYER VI3 ;
  RECT 601.480 6.340 601.680 6.540 ;
  LAYER VI3 ;
  RECT 601.480 5.940 601.680 6.140 ;
  LAYER VI3 ;
  RECT 601.080 6.340 601.280 6.540 ;
  LAYER VI3 ;
  RECT 601.080 5.940 601.280 6.140 ;
  LAYER VI3 ;
  RECT 622.160 5.880 630.160 6.740 ;
  LAYER VI3 ;
  RECT 629.760 6.340 629.960 6.540 ;
  LAYER VI3 ;
  RECT 629.760 5.940 629.960 6.140 ;
  LAYER VI3 ;
  RECT 629.360 6.340 629.560 6.540 ;
  LAYER VI3 ;
  RECT 629.360 5.940 629.560 6.140 ;
  LAYER VI3 ;
  RECT 628.960 6.340 629.160 6.540 ;
  LAYER VI3 ;
  RECT 628.960 5.940 629.160 6.140 ;
  LAYER VI3 ;
  RECT 628.560 6.340 628.760 6.540 ;
  LAYER VI3 ;
  RECT 628.560 5.940 628.760 6.140 ;
  LAYER VI3 ;
  RECT 628.160 6.340 628.360 6.540 ;
  LAYER VI3 ;
  RECT 628.160 5.940 628.360 6.140 ;
  LAYER VI3 ;
  RECT 627.760 6.340 627.960 6.540 ;
  LAYER VI3 ;
  RECT 627.760 5.940 627.960 6.140 ;
  LAYER VI3 ;
  RECT 627.360 6.340 627.560 6.540 ;
  LAYER VI3 ;
  RECT 627.360 5.940 627.560 6.140 ;
  LAYER VI3 ;
  RECT 626.960 6.340 627.160 6.540 ;
  LAYER VI3 ;
  RECT 626.960 5.940 627.160 6.140 ;
  LAYER VI3 ;
  RECT 626.560 6.340 626.760 6.540 ;
  LAYER VI3 ;
  RECT 626.560 5.940 626.760 6.140 ;
  LAYER VI3 ;
  RECT 626.160 6.340 626.360 6.540 ;
  LAYER VI3 ;
  RECT 626.160 5.940 626.360 6.140 ;
  LAYER VI3 ;
  RECT 625.760 6.340 625.960 6.540 ;
  LAYER VI3 ;
  RECT 625.760 5.940 625.960 6.140 ;
  LAYER VI3 ;
  RECT 625.360 6.340 625.560 6.540 ;
  LAYER VI3 ;
  RECT 625.360 5.940 625.560 6.140 ;
  LAYER VI3 ;
  RECT 624.960 6.340 625.160 6.540 ;
  LAYER VI3 ;
  RECT 624.960 5.940 625.160 6.140 ;
  LAYER VI3 ;
  RECT 624.560 6.340 624.760 6.540 ;
  LAYER VI3 ;
  RECT 624.560 5.940 624.760 6.140 ;
  LAYER VI3 ;
  RECT 624.160 6.340 624.360 6.540 ;
  LAYER VI3 ;
  RECT 624.160 5.940 624.360 6.140 ;
  LAYER VI3 ;
  RECT 623.760 6.340 623.960 6.540 ;
  LAYER VI3 ;
  RECT 623.760 5.940 623.960 6.140 ;
  LAYER VI3 ;
  RECT 623.360 6.340 623.560 6.540 ;
  LAYER VI3 ;
  RECT 623.360 5.940 623.560 6.140 ;
  LAYER VI3 ;
  RECT 622.960 6.340 623.160 6.540 ;
  LAYER VI3 ;
  RECT 622.960 5.940 623.160 6.140 ;
  LAYER VI3 ;
  RECT 622.560 6.340 622.760 6.540 ;
  LAYER VI3 ;
  RECT 622.560 5.940 622.760 6.140 ;
  LAYER VI3 ;
  RECT 622.160 6.340 622.360 6.540 ;
  LAYER VI3 ;
  RECT 622.160 5.940 622.360 6.140 ;
  LAYER VI3 ;
  RECT 642.000 5.880 650.000 6.740 ;
  LAYER VI3 ;
  RECT 649.600 6.340 649.800 6.540 ;
  LAYER VI3 ;
  RECT 649.600 5.940 649.800 6.140 ;
  LAYER VI3 ;
  RECT 649.200 6.340 649.400 6.540 ;
  LAYER VI3 ;
  RECT 649.200 5.940 649.400 6.140 ;
  LAYER VI3 ;
  RECT 648.800 6.340 649.000 6.540 ;
  LAYER VI3 ;
  RECT 648.800 5.940 649.000 6.140 ;
  LAYER VI3 ;
  RECT 648.400 6.340 648.600 6.540 ;
  LAYER VI3 ;
  RECT 648.400 5.940 648.600 6.140 ;
  LAYER VI3 ;
  RECT 648.000 6.340 648.200 6.540 ;
  LAYER VI3 ;
  RECT 648.000 5.940 648.200 6.140 ;
  LAYER VI3 ;
  RECT 647.600 6.340 647.800 6.540 ;
  LAYER VI3 ;
  RECT 647.600 5.940 647.800 6.140 ;
  LAYER VI3 ;
  RECT 647.200 6.340 647.400 6.540 ;
  LAYER VI3 ;
  RECT 647.200 5.940 647.400 6.140 ;
  LAYER VI3 ;
  RECT 646.800 6.340 647.000 6.540 ;
  LAYER VI3 ;
  RECT 646.800 5.940 647.000 6.140 ;
  LAYER VI3 ;
  RECT 646.400 6.340 646.600 6.540 ;
  LAYER VI3 ;
  RECT 646.400 5.940 646.600 6.140 ;
  LAYER VI3 ;
  RECT 646.000 6.340 646.200 6.540 ;
  LAYER VI3 ;
  RECT 646.000 5.940 646.200 6.140 ;
  LAYER VI3 ;
  RECT 645.600 6.340 645.800 6.540 ;
  LAYER VI3 ;
  RECT 645.600 5.940 645.800 6.140 ;
  LAYER VI3 ;
  RECT 645.200 6.340 645.400 6.540 ;
  LAYER VI3 ;
  RECT 645.200 5.940 645.400 6.140 ;
  LAYER VI3 ;
  RECT 644.800 6.340 645.000 6.540 ;
  LAYER VI3 ;
  RECT 644.800 5.940 645.000 6.140 ;
  LAYER VI3 ;
  RECT 644.400 6.340 644.600 6.540 ;
  LAYER VI3 ;
  RECT 644.400 5.940 644.600 6.140 ;
  LAYER VI3 ;
  RECT 644.000 6.340 644.200 6.540 ;
  LAYER VI3 ;
  RECT 644.000 5.940 644.200 6.140 ;
  LAYER VI3 ;
  RECT 643.600 6.340 643.800 6.540 ;
  LAYER VI3 ;
  RECT 643.600 5.940 643.800 6.140 ;
  LAYER VI3 ;
  RECT 643.200 6.340 643.400 6.540 ;
  LAYER VI3 ;
  RECT 643.200 5.940 643.400 6.140 ;
  LAYER VI3 ;
  RECT 642.800 6.340 643.000 6.540 ;
  LAYER VI3 ;
  RECT 642.800 5.940 643.000 6.140 ;
  LAYER VI3 ;
  RECT 642.400 6.340 642.600 6.540 ;
  LAYER VI3 ;
  RECT 642.400 5.940 642.600 6.140 ;
  LAYER VI3 ;
  RECT 642.000 6.340 642.200 6.540 ;
  LAYER VI3 ;
  RECT 642.000 5.940 642.200 6.140 ;
  LAYER VI3 ;
  RECT 663.080 5.880 671.080 6.740 ;
  LAYER VI3 ;
  RECT 670.680 6.340 670.880 6.540 ;
  LAYER VI3 ;
  RECT 670.680 5.940 670.880 6.140 ;
  LAYER VI3 ;
  RECT 670.280 6.340 670.480 6.540 ;
  LAYER VI3 ;
  RECT 670.280 5.940 670.480 6.140 ;
  LAYER VI3 ;
  RECT 669.880 6.340 670.080 6.540 ;
  LAYER VI3 ;
  RECT 669.880 5.940 670.080 6.140 ;
  LAYER VI3 ;
  RECT 669.480 6.340 669.680 6.540 ;
  LAYER VI3 ;
  RECT 669.480 5.940 669.680 6.140 ;
  LAYER VI3 ;
  RECT 669.080 6.340 669.280 6.540 ;
  LAYER VI3 ;
  RECT 669.080 5.940 669.280 6.140 ;
  LAYER VI3 ;
  RECT 668.680 6.340 668.880 6.540 ;
  LAYER VI3 ;
  RECT 668.680 5.940 668.880 6.140 ;
  LAYER VI3 ;
  RECT 668.280 6.340 668.480 6.540 ;
  LAYER VI3 ;
  RECT 668.280 5.940 668.480 6.140 ;
  LAYER VI3 ;
  RECT 667.880 6.340 668.080 6.540 ;
  LAYER VI3 ;
  RECT 667.880 5.940 668.080 6.140 ;
  LAYER VI3 ;
  RECT 667.480 6.340 667.680 6.540 ;
  LAYER VI3 ;
  RECT 667.480 5.940 667.680 6.140 ;
  LAYER VI3 ;
  RECT 667.080 6.340 667.280 6.540 ;
  LAYER VI3 ;
  RECT 667.080 5.940 667.280 6.140 ;
  LAYER VI3 ;
  RECT 666.680 6.340 666.880 6.540 ;
  LAYER VI3 ;
  RECT 666.680 5.940 666.880 6.140 ;
  LAYER VI3 ;
  RECT 666.280 6.340 666.480 6.540 ;
  LAYER VI3 ;
  RECT 666.280 5.940 666.480 6.140 ;
  LAYER VI3 ;
  RECT 665.880 6.340 666.080 6.540 ;
  LAYER VI3 ;
  RECT 665.880 5.940 666.080 6.140 ;
  LAYER VI3 ;
  RECT 665.480 6.340 665.680 6.540 ;
  LAYER VI3 ;
  RECT 665.480 5.940 665.680 6.140 ;
  LAYER VI3 ;
  RECT 665.080 6.340 665.280 6.540 ;
  LAYER VI3 ;
  RECT 665.080 5.940 665.280 6.140 ;
  LAYER VI3 ;
  RECT 664.680 6.340 664.880 6.540 ;
  LAYER VI3 ;
  RECT 664.680 5.940 664.880 6.140 ;
  LAYER VI3 ;
  RECT 664.280 6.340 664.480 6.540 ;
  LAYER VI3 ;
  RECT 664.280 5.940 664.480 6.140 ;
  LAYER VI3 ;
  RECT 663.880 6.340 664.080 6.540 ;
  LAYER VI3 ;
  RECT 663.880 5.940 664.080 6.140 ;
  LAYER VI3 ;
  RECT 663.480 6.340 663.680 6.540 ;
  LAYER VI3 ;
  RECT 663.480 5.940 663.680 6.140 ;
  LAYER VI3 ;
  RECT 663.080 6.340 663.280 6.540 ;
  LAYER VI3 ;
  RECT 663.080 5.940 663.280 6.140 ;
  LAYER VI3 ;
  RECT 682.920 5.880 690.920 6.740 ;
  LAYER VI3 ;
  RECT 690.520 6.340 690.720 6.540 ;
  LAYER VI3 ;
  RECT 690.520 5.940 690.720 6.140 ;
  LAYER VI3 ;
  RECT 690.120 6.340 690.320 6.540 ;
  LAYER VI3 ;
  RECT 690.120 5.940 690.320 6.140 ;
  LAYER VI3 ;
  RECT 689.720 6.340 689.920 6.540 ;
  LAYER VI3 ;
  RECT 689.720 5.940 689.920 6.140 ;
  LAYER VI3 ;
  RECT 689.320 6.340 689.520 6.540 ;
  LAYER VI3 ;
  RECT 689.320 5.940 689.520 6.140 ;
  LAYER VI3 ;
  RECT 688.920 6.340 689.120 6.540 ;
  LAYER VI3 ;
  RECT 688.920 5.940 689.120 6.140 ;
  LAYER VI3 ;
  RECT 688.520 6.340 688.720 6.540 ;
  LAYER VI3 ;
  RECT 688.520 5.940 688.720 6.140 ;
  LAYER VI3 ;
  RECT 688.120 6.340 688.320 6.540 ;
  LAYER VI3 ;
  RECT 688.120 5.940 688.320 6.140 ;
  LAYER VI3 ;
  RECT 687.720 6.340 687.920 6.540 ;
  LAYER VI3 ;
  RECT 687.720 5.940 687.920 6.140 ;
  LAYER VI3 ;
  RECT 687.320 6.340 687.520 6.540 ;
  LAYER VI3 ;
  RECT 687.320 5.940 687.520 6.140 ;
  LAYER VI3 ;
  RECT 686.920 6.340 687.120 6.540 ;
  LAYER VI3 ;
  RECT 686.920 5.940 687.120 6.140 ;
  LAYER VI3 ;
  RECT 686.520 6.340 686.720 6.540 ;
  LAYER VI3 ;
  RECT 686.520 5.940 686.720 6.140 ;
  LAYER VI3 ;
  RECT 686.120 6.340 686.320 6.540 ;
  LAYER VI3 ;
  RECT 686.120 5.940 686.320 6.140 ;
  LAYER VI3 ;
  RECT 685.720 6.340 685.920 6.540 ;
  LAYER VI3 ;
  RECT 685.720 5.940 685.920 6.140 ;
  LAYER VI3 ;
  RECT 685.320 6.340 685.520 6.540 ;
  LAYER VI3 ;
  RECT 685.320 5.940 685.520 6.140 ;
  LAYER VI3 ;
  RECT 684.920 6.340 685.120 6.540 ;
  LAYER VI3 ;
  RECT 684.920 5.940 685.120 6.140 ;
  LAYER VI3 ;
  RECT 684.520 6.340 684.720 6.540 ;
  LAYER VI3 ;
  RECT 684.520 5.940 684.720 6.140 ;
  LAYER VI3 ;
  RECT 684.120 6.340 684.320 6.540 ;
  LAYER VI3 ;
  RECT 684.120 5.940 684.320 6.140 ;
  LAYER VI3 ;
  RECT 683.720 6.340 683.920 6.540 ;
  LAYER VI3 ;
  RECT 683.720 5.940 683.920 6.140 ;
  LAYER VI3 ;
  RECT 683.320 6.340 683.520 6.540 ;
  LAYER VI3 ;
  RECT 683.320 5.940 683.520 6.140 ;
  LAYER VI3 ;
  RECT 682.920 6.340 683.120 6.540 ;
  LAYER VI3 ;
  RECT 682.920 5.940 683.120 6.140 ;
  LAYER VI3 ;
  RECT 704.000 5.880 712.000 6.740 ;
  LAYER VI3 ;
  RECT 711.600 6.340 711.800 6.540 ;
  LAYER VI3 ;
  RECT 711.600 5.940 711.800 6.140 ;
  LAYER VI3 ;
  RECT 711.200 6.340 711.400 6.540 ;
  LAYER VI3 ;
  RECT 711.200 5.940 711.400 6.140 ;
  LAYER VI3 ;
  RECT 710.800 6.340 711.000 6.540 ;
  LAYER VI3 ;
  RECT 710.800 5.940 711.000 6.140 ;
  LAYER VI3 ;
  RECT 710.400 6.340 710.600 6.540 ;
  LAYER VI3 ;
  RECT 710.400 5.940 710.600 6.140 ;
  LAYER VI3 ;
  RECT 710.000 6.340 710.200 6.540 ;
  LAYER VI3 ;
  RECT 710.000 5.940 710.200 6.140 ;
  LAYER VI3 ;
  RECT 709.600 6.340 709.800 6.540 ;
  LAYER VI3 ;
  RECT 709.600 5.940 709.800 6.140 ;
  LAYER VI3 ;
  RECT 709.200 6.340 709.400 6.540 ;
  LAYER VI3 ;
  RECT 709.200 5.940 709.400 6.140 ;
  LAYER VI3 ;
  RECT 708.800 6.340 709.000 6.540 ;
  LAYER VI3 ;
  RECT 708.800 5.940 709.000 6.140 ;
  LAYER VI3 ;
  RECT 708.400 6.340 708.600 6.540 ;
  LAYER VI3 ;
  RECT 708.400 5.940 708.600 6.140 ;
  LAYER VI3 ;
  RECT 708.000 6.340 708.200 6.540 ;
  LAYER VI3 ;
  RECT 708.000 5.940 708.200 6.140 ;
  LAYER VI3 ;
  RECT 707.600 6.340 707.800 6.540 ;
  LAYER VI3 ;
  RECT 707.600 5.940 707.800 6.140 ;
  LAYER VI3 ;
  RECT 707.200 6.340 707.400 6.540 ;
  LAYER VI3 ;
  RECT 707.200 5.940 707.400 6.140 ;
  LAYER VI3 ;
  RECT 706.800 6.340 707.000 6.540 ;
  LAYER VI3 ;
  RECT 706.800 5.940 707.000 6.140 ;
  LAYER VI3 ;
  RECT 706.400 6.340 706.600 6.540 ;
  LAYER VI3 ;
  RECT 706.400 5.940 706.600 6.140 ;
  LAYER VI3 ;
  RECT 706.000 6.340 706.200 6.540 ;
  LAYER VI3 ;
  RECT 706.000 5.940 706.200 6.140 ;
  LAYER VI3 ;
  RECT 705.600 6.340 705.800 6.540 ;
  LAYER VI3 ;
  RECT 705.600 5.940 705.800 6.140 ;
  LAYER VI3 ;
  RECT 705.200 6.340 705.400 6.540 ;
  LAYER VI3 ;
  RECT 705.200 5.940 705.400 6.140 ;
  LAYER VI3 ;
  RECT 704.800 6.340 705.000 6.540 ;
  LAYER VI3 ;
  RECT 704.800 5.940 705.000 6.140 ;
  LAYER VI3 ;
  RECT 704.400 6.340 704.600 6.540 ;
  LAYER VI3 ;
  RECT 704.400 5.940 704.600 6.140 ;
  LAYER VI3 ;
  RECT 704.000 6.340 704.200 6.540 ;
  LAYER VI3 ;
  RECT 704.000 5.940 704.200 6.140 ;
  LAYER VI3 ;
  RECT 723.840 5.880 731.840 6.740 ;
  LAYER VI3 ;
  RECT 731.440 6.340 731.640 6.540 ;
  LAYER VI3 ;
  RECT 731.440 5.940 731.640 6.140 ;
  LAYER VI3 ;
  RECT 731.040 6.340 731.240 6.540 ;
  LAYER VI3 ;
  RECT 731.040 5.940 731.240 6.140 ;
  LAYER VI3 ;
  RECT 730.640 6.340 730.840 6.540 ;
  LAYER VI3 ;
  RECT 730.640 5.940 730.840 6.140 ;
  LAYER VI3 ;
  RECT 730.240 6.340 730.440 6.540 ;
  LAYER VI3 ;
  RECT 730.240 5.940 730.440 6.140 ;
  LAYER VI3 ;
  RECT 729.840 6.340 730.040 6.540 ;
  LAYER VI3 ;
  RECT 729.840 5.940 730.040 6.140 ;
  LAYER VI3 ;
  RECT 729.440 6.340 729.640 6.540 ;
  LAYER VI3 ;
  RECT 729.440 5.940 729.640 6.140 ;
  LAYER VI3 ;
  RECT 729.040 6.340 729.240 6.540 ;
  LAYER VI3 ;
  RECT 729.040 5.940 729.240 6.140 ;
  LAYER VI3 ;
  RECT 728.640 6.340 728.840 6.540 ;
  LAYER VI3 ;
  RECT 728.640 5.940 728.840 6.140 ;
  LAYER VI3 ;
  RECT 728.240 6.340 728.440 6.540 ;
  LAYER VI3 ;
  RECT 728.240 5.940 728.440 6.140 ;
  LAYER VI3 ;
  RECT 727.840 6.340 728.040 6.540 ;
  LAYER VI3 ;
  RECT 727.840 5.940 728.040 6.140 ;
  LAYER VI3 ;
  RECT 727.440 6.340 727.640 6.540 ;
  LAYER VI3 ;
  RECT 727.440 5.940 727.640 6.140 ;
  LAYER VI3 ;
  RECT 727.040 6.340 727.240 6.540 ;
  LAYER VI3 ;
  RECT 727.040 5.940 727.240 6.140 ;
  LAYER VI3 ;
  RECT 726.640 6.340 726.840 6.540 ;
  LAYER VI3 ;
  RECT 726.640 5.940 726.840 6.140 ;
  LAYER VI3 ;
  RECT 726.240 6.340 726.440 6.540 ;
  LAYER VI3 ;
  RECT 726.240 5.940 726.440 6.140 ;
  LAYER VI3 ;
  RECT 725.840 6.340 726.040 6.540 ;
  LAYER VI3 ;
  RECT 725.840 5.940 726.040 6.140 ;
  LAYER VI3 ;
  RECT 725.440 6.340 725.640 6.540 ;
  LAYER VI3 ;
  RECT 725.440 5.940 725.640 6.140 ;
  LAYER VI3 ;
  RECT 725.040 6.340 725.240 6.540 ;
  LAYER VI3 ;
  RECT 725.040 5.940 725.240 6.140 ;
  LAYER VI3 ;
  RECT 724.640 6.340 724.840 6.540 ;
  LAYER VI3 ;
  RECT 724.640 5.940 724.840 6.140 ;
  LAYER VI3 ;
  RECT 724.240 6.340 724.440 6.540 ;
  LAYER VI3 ;
  RECT 724.240 5.940 724.440 6.140 ;
  LAYER VI3 ;
  RECT 723.840 6.340 724.040 6.540 ;
  LAYER VI3 ;
  RECT 723.840 5.940 724.040 6.140 ;
  LAYER VI3 ;
  RECT 744.920 5.880 752.920 6.740 ;
  LAYER VI3 ;
  RECT 752.520 6.340 752.720 6.540 ;
  LAYER VI3 ;
  RECT 752.520 5.940 752.720 6.140 ;
  LAYER VI3 ;
  RECT 752.120 6.340 752.320 6.540 ;
  LAYER VI3 ;
  RECT 752.120 5.940 752.320 6.140 ;
  LAYER VI3 ;
  RECT 751.720 6.340 751.920 6.540 ;
  LAYER VI3 ;
  RECT 751.720 5.940 751.920 6.140 ;
  LAYER VI3 ;
  RECT 751.320 6.340 751.520 6.540 ;
  LAYER VI3 ;
  RECT 751.320 5.940 751.520 6.140 ;
  LAYER VI3 ;
  RECT 750.920 6.340 751.120 6.540 ;
  LAYER VI3 ;
  RECT 750.920 5.940 751.120 6.140 ;
  LAYER VI3 ;
  RECT 750.520 6.340 750.720 6.540 ;
  LAYER VI3 ;
  RECT 750.520 5.940 750.720 6.140 ;
  LAYER VI3 ;
  RECT 750.120 6.340 750.320 6.540 ;
  LAYER VI3 ;
  RECT 750.120 5.940 750.320 6.140 ;
  LAYER VI3 ;
  RECT 749.720 6.340 749.920 6.540 ;
  LAYER VI3 ;
  RECT 749.720 5.940 749.920 6.140 ;
  LAYER VI3 ;
  RECT 749.320 6.340 749.520 6.540 ;
  LAYER VI3 ;
  RECT 749.320 5.940 749.520 6.140 ;
  LAYER VI3 ;
  RECT 748.920 6.340 749.120 6.540 ;
  LAYER VI3 ;
  RECT 748.920 5.940 749.120 6.140 ;
  LAYER VI3 ;
  RECT 748.520 6.340 748.720 6.540 ;
  LAYER VI3 ;
  RECT 748.520 5.940 748.720 6.140 ;
  LAYER VI3 ;
  RECT 748.120 6.340 748.320 6.540 ;
  LAYER VI3 ;
  RECT 748.120 5.940 748.320 6.140 ;
  LAYER VI3 ;
  RECT 747.720 6.340 747.920 6.540 ;
  LAYER VI3 ;
  RECT 747.720 5.940 747.920 6.140 ;
  LAYER VI3 ;
  RECT 747.320 6.340 747.520 6.540 ;
  LAYER VI3 ;
  RECT 747.320 5.940 747.520 6.140 ;
  LAYER VI3 ;
  RECT 746.920 6.340 747.120 6.540 ;
  LAYER VI3 ;
  RECT 746.920 5.940 747.120 6.140 ;
  LAYER VI3 ;
  RECT 746.520 6.340 746.720 6.540 ;
  LAYER VI3 ;
  RECT 746.520 5.940 746.720 6.140 ;
  LAYER VI3 ;
  RECT 746.120 6.340 746.320 6.540 ;
  LAYER VI3 ;
  RECT 746.120 5.940 746.320 6.140 ;
  LAYER VI3 ;
  RECT 745.720 6.340 745.920 6.540 ;
  LAYER VI3 ;
  RECT 745.720 5.940 745.920 6.140 ;
  LAYER VI3 ;
  RECT 745.320 6.340 745.520 6.540 ;
  LAYER VI3 ;
  RECT 745.320 5.940 745.520 6.140 ;
  LAYER VI3 ;
  RECT 744.920 6.340 745.120 6.540 ;
  LAYER VI3 ;
  RECT 744.920 5.940 745.120 6.140 ;
  LAYER VI3 ;
  RECT 764.760 5.880 772.760 6.740 ;
  LAYER VI3 ;
  RECT 772.360 6.340 772.560 6.540 ;
  LAYER VI3 ;
  RECT 772.360 5.940 772.560 6.140 ;
  LAYER VI3 ;
  RECT 771.960 6.340 772.160 6.540 ;
  LAYER VI3 ;
  RECT 771.960 5.940 772.160 6.140 ;
  LAYER VI3 ;
  RECT 771.560 6.340 771.760 6.540 ;
  LAYER VI3 ;
  RECT 771.560 5.940 771.760 6.140 ;
  LAYER VI3 ;
  RECT 771.160 6.340 771.360 6.540 ;
  LAYER VI3 ;
  RECT 771.160 5.940 771.360 6.140 ;
  LAYER VI3 ;
  RECT 770.760 6.340 770.960 6.540 ;
  LAYER VI3 ;
  RECT 770.760 5.940 770.960 6.140 ;
  LAYER VI3 ;
  RECT 770.360 6.340 770.560 6.540 ;
  LAYER VI3 ;
  RECT 770.360 5.940 770.560 6.140 ;
  LAYER VI3 ;
  RECT 769.960 6.340 770.160 6.540 ;
  LAYER VI3 ;
  RECT 769.960 5.940 770.160 6.140 ;
  LAYER VI3 ;
  RECT 769.560 6.340 769.760 6.540 ;
  LAYER VI3 ;
  RECT 769.560 5.940 769.760 6.140 ;
  LAYER VI3 ;
  RECT 769.160 6.340 769.360 6.540 ;
  LAYER VI3 ;
  RECT 769.160 5.940 769.360 6.140 ;
  LAYER VI3 ;
  RECT 768.760 6.340 768.960 6.540 ;
  LAYER VI3 ;
  RECT 768.760 5.940 768.960 6.140 ;
  LAYER VI3 ;
  RECT 768.360 6.340 768.560 6.540 ;
  LAYER VI3 ;
  RECT 768.360 5.940 768.560 6.140 ;
  LAYER VI3 ;
  RECT 767.960 6.340 768.160 6.540 ;
  LAYER VI3 ;
  RECT 767.960 5.940 768.160 6.140 ;
  LAYER VI3 ;
  RECT 767.560 6.340 767.760 6.540 ;
  LAYER VI3 ;
  RECT 767.560 5.940 767.760 6.140 ;
  LAYER VI3 ;
  RECT 767.160 6.340 767.360 6.540 ;
  LAYER VI3 ;
  RECT 767.160 5.940 767.360 6.140 ;
  LAYER VI3 ;
  RECT 766.760 6.340 766.960 6.540 ;
  LAYER VI3 ;
  RECT 766.760 5.940 766.960 6.140 ;
  LAYER VI3 ;
  RECT 766.360 6.340 766.560 6.540 ;
  LAYER VI3 ;
  RECT 766.360 5.940 766.560 6.140 ;
  LAYER VI3 ;
  RECT 765.960 6.340 766.160 6.540 ;
  LAYER VI3 ;
  RECT 765.960 5.940 766.160 6.140 ;
  LAYER VI3 ;
  RECT 765.560 6.340 765.760 6.540 ;
  LAYER VI3 ;
  RECT 765.560 5.940 765.760 6.140 ;
  LAYER VI3 ;
  RECT 765.160 6.340 765.360 6.540 ;
  LAYER VI3 ;
  RECT 765.160 5.940 765.360 6.140 ;
  LAYER VI3 ;
  RECT 764.760 6.340 764.960 6.540 ;
  LAYER VI3 ;
  RECT 764.760 5.940 764.960 6.140 ;
  LAYER VI3 ;
  RECT 785.840 5.880 793.840 6.740 ;
  LAYER VI3 ;
  RECT 793.440 6.340 793.640 6.540 ;
  LAYER VI3 ;
  RECT 793.440 5.940 793.640 6.140 ;
  LAYER VI3 ;
  RECT 793.040 6.340 793.240 6.540 ;
  LAYER VI3 ;
  RECT 793.040 5.940 793.240 6.140 ;
  LAYER VI3 ;
  RECT 792.640 6.340 792.840 6.540 ;
  LAYER VI3 ;
  RECT 792.640 5.940 792.840 6.140 ;
  LAYER VI3 ;
  RECT 792.240 6.340 792.440 6.540 ;
  LAYER VI3 ;
  RECT 792.240 5.940 792.440 6.140 ;
  LAYER VI3 ;
  RECT 791.840 6.340 792.040 6.540 ;
  LAYER VI3 ;
  RECT 791.840 5.940 792.040 6.140 ;
  LAYER VI3 ;
  RECT 791.440 6.340 791.640 6.540 ;
  LAYER VI3 ;
  RECT 791.440 5.940 791.640 6.140 ;
  LAYER VI3 ;
  RECT 791.040 6.340 791.240 6.540 ;
  LAYER VI3 ;
  RECT 791.040 5.940 791.240 6.140 ;
  LAYER VI3 ;
  RECT 790.640 6.340 790.840 6.540 ;
  LAYER VI3 ;
  RECT 790.640 5.940 790.840 6.140 ;
  LAYER VI3 ;
  RECT 790.240 6.340 790.440 6.540 ;
  LAYER VI3 ;
  RECT 790.240 5.940 790.440 6.140 ;
  LAYER VI3 ;
  RECT 789.840 6.340 790.040 6.540 ;
  LAYER VI3 ;
  RECT 789.840 5.940 790.040 6.140 ;
  LAYER VI3 ;
  RECT 789.440 6.340 789.640 6.540 ;
  LAYER VI3 ;
  RECT 789.440 5.940 789.640 6.140 ;
  LAYER VI3 ;
  RECT 789.040 6.340 789.240 6.540 ;
  LAYER VI3 ;
  RECT 789.040 5.940 789.240 6.140 ;
  LAYER VI3 ;
  RECT 788.640 6.340 788.840 6.540 ;
  LAYER VI3 ;
  RECT 788.640 5.940 788.840 6.140 ;
  LAYER VI3 ;
  RECT 788.240 6.340 788.440 6.540 ;
  LAYER VI3 ;
  RECT 788.240 5.940 788.440 6.140 ;
  LAYER VI3 ;
  RECT 787.840 6.340 788.040 6.540 ;
  LAYER VI3 ;
  RECT 787.840 5.940 788.040 6.140 ;
  LAYER VI3 ;
  RECT 787.440 6.340 787.640 6.540 ;
  LAYER VI3 ;
  RECT 787.440 5.940 787.640 6.140 ;
  LAYER VI3 ;
  RECT 787.040 6.340 787.240 6.540 ;
  LAYER VI3 ;
  RECT 787.040 5.940 787.240 6.140 ;
  LAYER VI3 ;
  RECT 786.640 6.340 786.840 6.540 ;
  LAYER VI3 ;
  RECT 786.640 5.940 786.840 6.140 ;
  LAYER VI3 ;
  RECT 786.240 6.340 786.440 6.540 ;
  LAYER VI3 ;
  RECT 786.240 5.940 786.440 6.140 ;
  LAYER VI3 ;
  RECT 785.840 6.340 786.040 6.540 ;
  LAYER VI3 ;
  RECT 785.840 5.940 786.040 6.140 ;
  LAYER VI3 ;
  RECT 805.680 5.880 813.680 6.740 ;
  LAYER VI3 ;
  RECT 813.280 6.340 813.480 6.540 ;
  LAYER VI3 ;
  RECT 813.280 5.940 813.480 6.140 ;
  LAYER VI3 ;
  RECT 812.880 6.340 813.080 6.540 ;
  LAYER VI3 ;
  RECT 812.880 5.940 813.080 6.140 ;
  LAYER VI3 ;
  RECT 812.480 6.340 812.680 6.540 ;
  LAYER VI3 ;
  RECT 812.480 5.940 812.680 6.140 ;
  LAYER VI3 ;
  RECT 812.080 6.340 812.280 6.540 ;
  LAYER VI3 ;
  RECT 812.080 5.940 812.280 6.140 ;
  LAYER VI3 ;
  RECT 811.680 6.340 811.880 6.540 ;
  LAYER VI3 ;
  RECT 811.680 5.940 811.880 6.140 ;
  LAYER VI3 ;
  RECT 811.280 6.340 811.480 6.540 ;
  LAYER VI3 ;
  RECT 811.280 5.940 811.480 6.140 ;
  LAYER VI3 ;
  RECT 810.880 6.340 811.080 6.540 ;
  LAYER VI3 ;
  RECT 810.880 5.940 811.080 6.140 ;
  LAYER VI3 ;
  RECT 810.480 6.340 810.680 6.540 ;
  LAYER VI3 ;
  RECT 810.480 5.940 810.680 6.140 ;
  LAYER VI3 ;
  RECT 810.080 6.340 810.280 6.540 ;
  LAYER VI3 ;
  RECT 810.080 5.940 810.280 6.140 ;
  LAYER VI3 ;
  RECT 809.680 6.340 809.880 6.540 ;
  LAYER VI3 ;
  RECT 809.680 5.940 809.880 6.140 ;
  LAYER VI3 ;
  RECT 809.280 6.340 809.480 6.540 ;
  LAYER VI3 ;
  RECT 809.280 5.940 809.480 6.140 ;
  LAYER VI3 ;
  RECT 808.880 6.340 809.080 6.540 ;
  LAYER VI3 ;
  RECT 808.880 5.940 809.080 6.140 ;
  LAYER VI3 ;
  RECT 808.480 6.340 808.680 6.540 ;
  LAYER VI3 ;
  RECT 808.480 5.940 808.680 6.140 ;
  LAYER VI3 ;
  RECT 808.080 6.340 808.280 6.540 ;
  LAYER VI3 ;
  RECT 808.080 5.940 808.280 6.140 ;
  LAYER VI3 ;
  RECT 807.680 6.340 807.880 6.540 ;
  LAYER VI3 ;
  RECT 807.680 5.940 807.880 6.140 ;
  LAYER VI3 ;
  RECT 807.280 6.340 807.480 6.540 ;
  LAYER VI3 ;
  RECT 807.280 5.940 807.480 6.140 ;
  LAYER VI3 ;
  RECT 806.880 6.340 807.080 6.540 ;
  LAYER VI3 ;
  RECT 806.880 5.940 807.080 6.140 ;
  LAYER VI3 ;
  RECT 806.480 6.340 806.680 6.540 ;
  LAYER VI3 ;
  RECT 806.480 5.940 806.680 6.140 ;
  LAYER VI3 ;
  RECT 806.080 6.340 806.280 6.540 ;
  LAYER VI3 ;
  RECT 806.080 5.940 806.280 6.140 ;
  LAYER VI3 ;
  RECT 805.680 6.340 805.880 6.540 ;
  LAYER VI3 ;
  RECT 805.680 5.940 805.880 6.140 ;
  LAYER VI3 ;
  RECT 826.760 5.880 834.760 6.740 ;
  LAYER VI3 ;
  RECT 834.360 6.340 834.560 6.540 ;
  LAYER VI3 ;
  RECT 834.360 5.940 834.560 6.140 ;
  LAYER VI3 ;
  RECT 833.960 6.340 834.160 6.540 ;
  LAYER VI3 ;
  RECT 833.960 5.940 834.160 6.140 ;
  LAYER VI3 ;
  RECT 833.560 6.340 833.760 6.540 ;
  LAYER VI3 ;
  RECT 833.560 5.940 833.760 6.140 ;
  LAYER VI3 ;
  RECT 833.160 6.340 833.360 6.540 ;
  LAYER VI3 ;
  RECT 833.160 5.940 833.360 6.140 ;
  LAYER VI3 ;
  RECT 832.760 6.340 832.960 6.540 ;
  LAYER VI3 ;
  RECT 832.760 5.940 832.960 6.140 ;
  LAYER VI3 ;
  RECT 832.360 6.340 832.560 6.540 ;
  LAYER VI3 ;
  RECT 832.360 5.940 832.560 6.140 ;
  LAYER VI3 ;
  RECT 831.960 6.340 832.160 6.540 ;
  LAYER VI3 ;
  RECT 831.960 5.940 832.160 6.140 ;
  LAYER VI3 ;
  RECT 831.560 6.340 831.760 6.540 ;
  LAYER VI3 ;
  RECT 831.560 5.940 831.760 6.140 ;
  LAYER VI3 ;
  RECT 831.160 6.340 831.360 6.540 ;
  LAYER VI3 ;
  RECT 831.160 5.940 831.360 6.140 ;
  LAYER VI3 ;
  RECT 830.760 6.340 830.960 6.540 ;
  LAYER VI3 ;
  RECT 830.760 5.940 830.960 6.140 ;
  LAYER VI3 ;
  RECT 830.360 6.340 830.560 6.540 ;
  LAYER VI3 ;
  RECT 830.360 5.940 830.560 6.140 ;
  LAYER VI3 ;
  RECT 829.960 6.340 830.160 6.540 ;
  LAYER VI3 ;
  RECT 829.960 5.940 830.160 6.140 ;
  LAYER VI3 ;
  RECT 829.560 6.340 829.760 6.540 ;
  LAYER VI3 ;
  RECT 829.560 5.940 829.760 6.140 ;
  LAYER VI3 ;
  RECT 829.160 6.340 829.360 6.540 ;
  LAYER VI3 ;
  RECT 829.160 5.940 829.360 6.140 ;
  LAYER VI3 ;
  RECT 828.760 6.340 828.960 6.540 ;
  LAYER VI3 ;
  RECT 828.760 5.940 828.960 6.140 ;
  LAYER VI3 ;
  RECT 828.360 6.340 828.560 6.540 ;
  LAYER VI3 ;
  RECT 828.360 5.940 828.560 6.140 ;
  LAYER VI3 ;
  RECT 827.960 6.340 828.160 6.540 ;
  LAYER VI3 ;
  RECT 827.960 5.940 828.160 6.140 ;
  LAYER VI3 ;
  RECT 827.560 6.340 827.760 6.540 ;
  LAYER VI3 ;
  RECT 827.560 5.940 827.760 6.140 ;
  LAYER VI3 ;
  RECT 827.160 6.340 827.360 6.540 ;
  LAYER VI3 ;
  RECT 827.160 5.940 827.360 6.140 ;
  LAYER VI3 ;
  RECT 826.760 6.340 826.960 6.540 ;
  LAYER VI3 ;
  RECT 826.760 5.940 826.960 6.140 ;
  LAYER VI3 ;
  RECT 846.600 5.880 854.600 6.740 ;
  LAYER VI3 ;
  RECT 854.200 6.340 854.400 6.540 ;
  LAYER VI3 ;
  RECT 854.200 5.940 854.400 6.140 ;
  LAYER VI3 ;
  RECT 853.800 6.340 854.000 6.540 ;
  LAYER VI3 ;
  RECT 853.800 5.940 854.000 6.140 ;
  LAYER VI3 ;
  RECT 853.400 6.340 853.600 6.540 ;
  LAYER VI3 ;
  RECT 853.400 5.940 853.600 6.140 ;
  LAYER VI3 ;
  RECT 853.000 6.340 853.200 6.540 ;
  LAYER VI3 ;
  RECT 853.000 5.940 853.200 6.140 ;
  LAYER VI3 ;
  RECT 852.600 6.340 852.800 6.540 ;
  LAYER VI3 ;
  RECT 852.600 5.940 852.800 6.140 ;
  LAYER VI3 ;
  RECT 852.200 6.340 852.400 6.540 ;
  LAYER VI3 ;
  RECT 852.200 5.940 852.400 6.140 ;
  LAYER VI3 ;
  RECT 851.800 6.340 852.000 6.540 ;
  LAYER VI3 ;
  RECT 851.800 5.940 852.000 6.140 ;
  LAYER VI3 ;
  RECT 851.400 6.340 851.600 6.540 ;
  LAYER VI3 ;
  RECT 851.400 5.940 851.600 6.140 ;
  LAYER VI3 ;
  RECT 851.000 6.340 851.200 6.540 ;
  LAYER VI3 ;
  RECT 851.000 5.940 851.200 6.140 ;
  LAYER VI3 ;
  RECT 850.600 6.340 850.800 6.540 ;
  LAYER VI3 ;
  RECT 850.600 5.940 850.800 6.140 ;
  LAYER VI3 ;
  RECT 850.200 6.340 850.400 6.540 ;
  LAYER VI3 ;
  RECT 850.200 5.940 850.400 6.140 ;
  LAYER VI3 ;
  RECT 849.800 6.340 850.000 6.540 ;
  LAYER VI3 ;
  RECT 849.800 5.940 850.000 6.140 ;
  LAYER VI3 ;
  RECT 849.400 6.340 849.600 6.540 ;
  LAYER VI3 ;
  RECT 849.400 5.940 849.600 6.140 ;
  LAYER VI3 ;
  RECT 849.000 6.340 849.200 6.540 ;
  LAYER VI3 ;
  RECT 849.000 5.940 849.200 6.140 ;
  LAYER VI3 ;
  RECT 848.600 6.340 848.800 6.540 ;
  LAYER VI3 ;
  RECT 848.600 5.940 848.800 6.140 ;
  LAYER VI3 ;
  RECT 848.200 6.340 848.400 6.540 ;
  LAYER VI3 ;
  RECT 848.200 5.940 848.400 6.140 ;
  LAYER VI3 ;
  RECT 847.800 6.340 848.000 6.540 ;
  LAYER VI3 ;
  RECT 847.800 5.940 848.000 6.140 ;
  LAYER VI3 ;
  RECT 847.400 6.340 847.600 6.540 ;
  LAYER VI3 ;
  RECT 847.400 5.940 847.600 6.140 ;
  LAYER VI3 ;
  RECT 847.000 6.340 847.200 6.540 ;
  LAYER VI3 ;
  RECT 847.000 5.940 847.200 6.140 ;
  LAYER VI3 ;
  RECT 846.600 6.340 846.800 6.540 ;
  LAYER VI3 ;
  RECT 846.600 5.940 846.800 6.140 ;
  LAYER VI3 ;
  RECT 867.680 5.880 875.680 6.740 ;
  LAYER VI3 ;
  RECT 875.280 6.340 875.480 6.540 ;
  LAYER VI3 ;
  RECT 875.280 5.940 875.480 6.140 ;
  LAYER VI3 ;
  RECT 874.880 6.340 875.080 6.540 ;
  LAYER VI3 ;
  RECT 874.880 5.940 875.080 6.140 ;
  LAYER VI3 ;
  RECT 874.480 6.340 874.680 6.540 ;
  LAYER VI3 ;
  RECT 874.480 5.940 874.680 6.140 ;
  LAYER VI3 ;
  RECT 874.080 6.340 874.280 6.540 ;
  LAYER VI3 ;
  RECT 874.080 5.940 874.280 6.140 ;
  LAYER VI3 ;
  RECT 873.680 6.340 873.880 6.540 ;
  LAYER VI3 ;
  RECT 873.680 5.940 873.880 6.140 ;
  LAYER VI3 ;
  RECT 873.280 6.340 873.480 6.540 ;
  LAYER VI3 ;
  RECT 873.280 5.940 873.480 6.140 ;
  LAYER VI3 ;
  RECT 872.880 6.340 873.080 6.540 ;
  LAYER VI3 ;
  RECT 872.880 5.940 873.080 6.140 ;
  LAYER VI3 ;
  RECT 872.480 6.340 872.680 6.540 ;
  LAYER VI3 ;
  RECT 872.480 5.940 872.680 6.140 ;
  LAYER VI3 ;
  RECT 872.080 6.340 872.280 6.540 ;
  LAYER VI3 ;
  RECT 872.080 5.940 872.280 6.140 ;
  LAYER VI3 ;
  RECT 871.680 6.340 871.880 6.540 ;
  LAYER VI3 ;
  RECT 871.680 5.940 871.880 6.140 ;
  LAYER VI3 ;
  RECT 871.280 6.340 871.480 6.540 ;
  LAYER VI3 ;
  RECT 871.280 5.940 871.480 6.140 ;
  LAYER VI3 ;
  RECT 870.880 6.340 871.080 6.540 ;
  LAYER VI3 ;
  RECT 870.880 5.940 871.080 6.140 ;
  LAYER VI3 ;
  RECT 870.480 6.340 870.680 6.540 ;
  LAYER VI3 ;
  RECT 870.480 5.940 870.680 6.140 ;
  LAYER VI3 ;
  RECT 870.080 6.340 870.280 6.540 ;
  LAYER VI3 ;
  RECT 870.080 5.940 870.280 6.140 ;
  LAYER VI3 ;
  RECT 869.680 6.340 869.880 6.540 ;
  LAYER VI3 ;
  RECT 869.680 5.940 869.880 6.140 ;
  LAYER VI3 ;
  RECT 869.280 6.340 869.480 6.540 ;
  LAYER VI3 ;
  RECT 869.280 5.940 869.480 6.140 ;
  LAYER VI3 ;
  RECT 868.880 6.340 869.080 6.540 ;
  LAYER VI3 ;
  RECT 868.880 5.940 869.080 6.140 ;
  LAYER VI3 ;
  RECT 868.480 6.340 868.680 6.540 ;
  LAYER VI3 ;
  RECT 868.480 5.940 868.680 6.140 ;
  LAYER VI3 ;
  RECT 868.080 6.340 868.280 6.540 ;
  LAYER VI3 ;
  RECT 868.080 5.940 868.280 6.140 ;
  LAYER VI3 ;
  RECT 867.680 6.340 867.880 6.540 ;
  LAYER VI3 ;
  RECT 867.680 5.940 867.880 6.140 ;
  LAYER VI3 ;
  RECT 887.520 5.880 895.520 6.740 ;
  LAYER VI3 ;
  RECT 895.120 6.340 895.320 6.540 ;
  LAYER VI3 ;
  RECT 895.120 5.940 895.320 6.140 ;
  LAYER VI3 ;
  RECT 894.720 6.340 894.920 6.540 ;
  LAYER VI3 ;
  RECT 894.720 5.940 894.920 6.140 ;
  LAYER VI3 ;
  RECT 894.320 6.340 894.520 6.540 ;
  LAYER VI3 ;
  RECT 894.320 5.940 894.520 6.140 ;
  LAYER VI3 ;
  RECT 893.920 6.340 894.120 6.540 ;
  LAYER VI3 ;
  RECT 893.920 5.940 894.120 6.140 ;
  LAYER VI3 ;
  RECT 893.520 6.340 893.720 6.540 ;
  LAYER VI3 ;
  RECT 893.520 5.940 893.720 6.140 ;
  LAYER VI3 ;
  RECT 893.120 6.340 893.320 6.540 ;
  LAYER VI3 ;
  RECT 893.120 5.940 893.320 6.140 ;
  LAYER VI3 ;
  RECT 892.720 6.340 892.920 6.540 ;
  LAYER VI3 ;
  RECT 892.720 5.940 892.920 6.140 ;
  LAYER VI3 ;
  RECT 892.320 6.340 892.520 6.540 ;
  LAYER VI3 ;
  RECT 892.320 5.940 892.520 6.140 ;
  LAYER VI3 ;
  RECT 891.920 6.340 892.120 6.540 ;
  LAYER VI3 ;
  RECT 891.920 5.940 892.120 6.140 ;
  LAYER VI3 ;
  RECT 891.520 6.340 891.720 6.540 ;
  LAYER VI3 ;
  RECT 891.520 5.940 891.720 6.140 ;
  LAYER VI3 ;
  RECT 891.120 6.340 891.320 6.540 ;
  LAYER VI3 ;
  RECT 891.120 5.940 891.320 6.140 ;
  LAYER VI3 ;
  RECT 890.720 6.340 890.920 6.540 ;
  LAYER VI3 ;
  RECT 890.720 5.940 890.920 6.140 ;
  LAYER VI3 ;
  RECT 890.320 6.340 890.520 6.540 ;
  LAYER VI3 ;
  RECT 890.320 5.940 890.520 6.140 ;
  LAYER VI3 ;
  RECT 889.920 6.340 890.120 6.540 ;
  LAYER VI3 ;
  RECT 889.920 5.940 890.120 6.140 ;
  LAYER VI3 ;
  RECT 889.520 6.340 889.720 6.540 ;
  LAYER VI3 ;
  RECT 889.520 5.940 889.720 6.140 ;
  LAYER VI3 ;
  RECT 889.120 6.340 889.320 6.540 ;
  LAYER VI3 ;
  RECT 889.120 5.940 889.320 6.140 ;
  LAYER VI3 ;
  RECT 888.720 6.340 888.920 6.540 ;
  LAYER VI3 ;
  RECT 888.720 5.940 888.920 6.140 ;
  LAYER VI3 ;
  RECT 888.320 6.340 888.520 6.540 ;
  LAYER VI3 ;
  RECT 888.320 5.940 888.520 6.140 ;
  LAYER VI3 ;
  RECT 887.920 6.340 888.120 6.540 ;
  LAYER VI3 ;
  RECT 887.920 5.940 888.120 6.140 ;
  LAYER VI3 ;
  RECT 887.520 6.340 887.720 6.540 ;
  LAYER VI3 ;
  RECT 887.520 5.940 887.720 6.140 ;
  LAYER VI3 ;
  RECT 908.600 5.880 916.600 6.740 ;
  LAYER VI3 ;
  RECT 916.200 6.340 916.400 6.540 ;
  LAYER VI3 ;
  RECT 916.200 5.940 916.400 6.140 ;
  LAYER VI3 ;
  RECT 915.800 6.340 916.000 6.540 ;
  LAYER VI3 ;
  RECT 915.800 5.940 916.000 6.140 ;
  LAYER VI3 ;
  RECT 915.400 6.340 915.600 6.540 ;
  LAYER VI3 ;
  RECT 915.400 5.940 915.600 6.140 ;
  LAYER VI3 ;
  RECT 915.000 6.340 915.200 6.540 ;
  LAYER VI3 ;
  RECT 915.000 5.940 915.200 6.140 ;
  LAYER VI3 ;
  RECT 914.600 6.340 914.800 6.540 ;
  LAYER VI3 ;
  RECT 914.600 5.940 914.800 6.140 ;
  LAYER VI3 ;
  RECT 914.200 6.340 914.400 6.540 ;
  LAYER VI3 ;
  RECT 914.200 5.940 914.400 6.140 ;
  LAYER VI3 ;
  RECT 913.800 6.340 914.000 6.540 ;
  LAYER VI3 ;
  RECT 913.800 5.940 914.000 6.140 ;
  LAYER VI3 ;
  RECT 913.400 6.340 913.600 6.540 ;
  LAYER VI3 ;
  RECT 913.400 5.940 913.600 6.140 ;
  LAYER VI3 ;
  RECT 913.000 6.340 913.200 6.540 ;
  LAYER VI3 ;
  RECT 913.000 5.940 913.200 6.140 ;
  LAYER VI3 ;
  RECT 912.600 6.340 912.800 6.540 ;
  LAYER VI3 ;
  RECT 912.600 5.940 912.800 6.140 ;
  LAYER VI3 ;
  RECT 912.200 6.340 912.400 6.540 ;
  LAYER VI3 ;
  RECT 912.200 5.940 912.400 6.140 ;
  LAYER VI3 ;
  RECT 911.800 6.340 912.000 6.540 ;
  LAYER VI3 ;
  RECT 911.800 5.940 912.000 6.140 ;
  LAYER VI3 ;
  RECT 911.400 6.340 911.600 6.540 ;
  LAYER VI3 ;
  RECT 911.400 5.940 911.600 6.140 ;
  LAYER VI3 ;
  RECT 911.000 6.340 911.200 6.540 ;
  LAYER VI3 ;
  RECT 911.000 5.940 911.200 6.140 ;
  LAYER VI3 ;
  RECT 910.600 6.340 910.800 6.540 ;
  LAYER VI3 ;
  RECT 910.600 5.940 910.800 6.140 ;
  LAYER VI3 ;
  RECT 910.200 6.340 910.400 6.540 ;
  LAYER VI3 ;
  RECT 910.200 5.940 910.400 6.140 ;
  LAYER VI3 ;
  RECT 909.800 6.340 910.000 6.540 ;
  LAYER VI3 ;
  RECT 909.800 5.940 910.000 6.140 ;
  LAYER VI3 ;
  RECT 909.400 6.340 909.600 6.540 ;
  LAYER VI3 ;
  RECT 909.400 5.940 909.600 6.140 ;
  LAYER VI3 ;
  RECT 909.000 6.340 909.200 6.540 ;
  LAYER VI3 ;
  RECT 909.000 5.940 909.200 6.140 ;
  LAYER VI3 ;
  RECT 908.600 6.340 908.800 6.540 ;
  LAYER VI3 ;
  RECT 908.600 5.940 908.800 6.140 ;
  LAYER VI3 ;
  RECT 928.440 5.880 936.440 6.740 ;
  LAYER VI3 ;
  RECT 936.040 6.340 936.240 6.540 ;
  LAYER VI3 ;
  RECT 936.040 5.940 936.240 6.140 ;
  LAYER VI3 ;
  RECT 935.640 6.340 935.840 6.540 ;
  LAYER VI3 ;
  RECT 935.640 5.940 935.840 6.140 ;
  LAYER VI3 ;
  RECT 935.240 6.340 935.440 6.540 ;
  LAYER VI3 ;
  RECT 935.240 5.940 935.440 6.140 ;
  LAYER VI3 ;
  RECT 934.840 6.340 935.040 6.540 ;
  LAYER VI3 ;
  RECT 934.840 5.940 935.040 6.140 ;
  LAYER VI3 ;
  RECT 934.440 6.340 934.640 6.540 ;
  LAYER VI3 ;
  RECT 934.440 5.940 934.640 6.140 ;
  LAYER VI3 ;
  RECT 934.040 6.340 934.240 6.540 ;
  LAYER VI3 ;
  RECT 934.040 5.940 934.240 6.140 ;
  LAYER VI3 ;
  RECT 933.640 6.340 933.840 6.540 ;
  LAYER VI3 ;
  RECT 933.640 5.940 933.840 6.140 ;
  LAYER VI3 ;
  RECT 933.240 6.340 933.440 6.540 ;
  LAYER VI3 ;
  RECT 933.240 5.940 933.440 6.140 ;
  LAYER VI3 ;
  RECT 932.840 6.340 933.040 6.540 ;
  LAYER VI3 ;
  RECT 932.840 5.940 933.040 6.140 ;
  LAYER VI3 ;
  RECT 932.440 6.340 932.640 6.540 ;
  LAYER VI3 ;
  RECT 932.440 5.940 932.640 6.140 ;
  LAYER VI3 ;
  RECT 932.040 6.340 932.240 6.540 ;
  LAYER VI3 ;
  RECT 932.040 5.940 932.240 6.140 ;
  LAYER VI3 ;
  RECT 931.640 6.340 931.840 6.540 ;
  LAYER VI3 ;
  RECT 931.640 5.940 931.840 6.140 ;
  LAYER VI3 ;
  RECT 931.240 6.340 931.440 6.540 ;
  LAYER VI3 ;
  RECT 931.240 5.940 931.440 6.140 ;
  LAYER VI3 ;
  RECT 930.840 6.340 931.040 6.540 ;
  LAYER VI3 ;
  RECT 930.840 5.940 931.040 6.140 ;
  LAYER VI3 ;
  RECT 930.440 6.340 930.640 6.540 ;
  LAYER VI3 ;
  RECT 930.440 5.940 930.640 6.140 ;
  LAYER VI3 ;
  RECT 930.040 6.340 930.240 6.540 ;
  LAYER VI3 ;
  RECT 930.040 5.940 930.240 6.140 ;
  LAYER VI3 ;
  RECT 929.640 6.340 929.840 6.540 ;
  LAYER VI3 ;
  RECT 929.640 5.940 929.840 6.140 ;
  LAYER VI3 ;
  RECT 929.240 6.340 929.440 6.540 ;
  LAYER VI3 ;
  RECT 929.240 5.940 929.440 6.140 ;
  LAYER VI3 ;
  RECT 928.840 6.340 929.040 6.540 ;
  LAYER VI3 ;
  RECT 928.840 5.940 929.040 6.140 ;
  LAYER VI3 ;
  RECT 928.440 6.340 928.640 6.540 ;
  LAYER VI3 ;
  RECT 928.440 5.940 928.640 6.140 ;
  LAYER VI3 ;
  RECT 949.520 5.880 957.520 6.740 ;
  LAYER VI3 ;
  RECT 957.120 6.340 957.320 6.540 ;
  LAYER VI3 ;
  RECT 957.120 5.940 957.320 6.140 ;
  LAYER VI3 ;
  RECT 956.720 6.340 956.920 6.540 ;
  LAYER VI3 ;
  RECT 956.720 5.940 956.920 6.140 ;
  LAYER VI3 ;
  RECT 956.320 6.340 956.520 6.540 ;
  LAYER VI3 ;
  RECT 956.320 5.940 956.520 6.140 ;
  LAYER VI3 ;
  RECT 955.920 6.340 956.120 6.540 ;
  LAYER VI3 ;
  RECT 955.920 5.940 956.120 6.140 ;
  LAYER VI3 ;
  RECT 955.520 6.340 955.720 6.540 ;
  LAYER VI3 ;
  RECT 955.520 5.940 955.720 6.140 ;
  LAYER VI3 ;
  RECT 955.120 6.340 955.320 6.540 ;
  LAYER VI3 ;
  RECT 955.120 5.940 955.320 6.140 ;
  LAYER VI3 ;
  RECT 954.720 6.340 954.920 6.540 ;
  LAYER VI3 ;
  RECT 954.720 5.940 954.920 6.140 ;
  LAYER VI3 ;
  RECT 954.320 6.340 954.520 6.540 ;
  LAYER VI3 ;
  RECT 954.320 5.940 954.520 6.140 ;
  LAYER VI3 ;
  RECT 953.920 6.340 954.120 6.540 ;
  LAYER VI3 ;
  RECT 953.920 5.940 954.120 6.140 ;
  LAYER VI3 ;
  RECT 953.520 6.340 953.720 6.540 ;
  LAYER VI3 ;
  RECT 953.520 5.940 953.720 6.140 ;
  LAYER VI3 ;
  RECT 953.120 6.340 953.320 6.540 ;
  LAYER VI3 ;
  RECT 953.120 5.940 953.320 6.140 ;
  LAYER VI3 ;
  RECT 952.720 6.340 952.920 6.540 ;
  LAYER VI3 ;
  RECT 952.720 5.940 952.920 6.140 ;
  LAYER VI3 ;
  RECT 952.320 6.340 952.520 6.540 ;
  LAYER VI3 ;
  RECT 952.320 5.940 952.520 6.140 ;
  LAYER VI3 ;
  RECT 951.920 6.340 952.120 6.540 ;
  LAYER VI3 ;
  RECT 951.920 5.940 952.120 6.140 ;
  LAYER VI3 ;
  RECT 951.520 6.340 951.720 6.540 ;
  LAYER VI3 ;
  RECT 951.520 5.940 951.720 6.140 ;
  LAYER VI3 ;
  RECT 951.120 6.340 951.320 6.540 ;
  LAYER VI3 ;
  RECT 951.120 5.940 951.320 6.140 ;
  LAYER VI3 ;
  RECT 950.720 6.340 950.920 6.540 ;
  LAYER VI3 ;
  RECT 950.720 5.940 950.920 6.140 ;
  LAYER VI3 ;
  RECT 950.320 6.340 950.520 6.540 ;
  LAYER VI3 ;
  RECT 950.320 5.940 950.520 6.140 ;
  LAYER VI3 ;
  RECT 949.920 6.340 950.120 6.540 ;
  LAYER VI3 ;
  RECT 949.920 5.940 950.120 6.140 ;
  LAYER VI3 ;
  RECT 949.520 6.340 949.720 6.540 ;
  LAYER VI3 ;
  RECT 949.520 5.940 949.720 6.140 ;
  LAYER VI3 ;
  RECT 969.360 5.880 977.360 6.740 ;
  LAYER VI3 ;
  RECT 976.960 6.340 977.160 6.540 ;
  LAYER VI3 ;
  RECT 976.960 5.940 977.160 6.140 ;
  LAYER VI3 ;
  RECT 976.560 6.340 976.760 6.540 ;
  LAYER VI3 ;
  RECT 976.560 5.940 976.760 6.140 ;
  LAYER VI3 ;
  RECT 976.160 6.340 976.360 6.540 ;
  LAYER VI3 ;
  RECT 976.160 5.940 976.360 6.140 ;
  LAYER VI3 ;
  RECT 975.760 6.340 975.960 6.540 ;
  LAYER VI3 ;
  RECT 975.760 5.940 975.960 6.140 ;
  LAYER VI3 ;
  RECT 975.360 6.340 975.560 6.540 ;
  LAYER VI3 ;
  RECT 975.360 5.940 975.560 6.140 ;
  LAYER VI3 ;
  RECT 974.960 6.340 975.160 6.540 ;
  LAYER VI3 ;
  RECT 974.960 5.940 975.160 6.140 ;
  LAYER VI3 ;
  RECT 974.560 6.340 974.760 6.540 ;
  LAYER VI3 ;
  RECT 974.560 5.940 974.760 6.140 ;
  LAYER VI3 ;
  RECT 974.160 6.340 974.360 6.540 ;
  LAYER VI3 ;
  RECT 974.160 5.940 974.360 6.140 ;
  LAYER VI3 ;
  RECT 973.760 6.340 973.960 6.540 ;
  LAYER VI3 ;
  RECT 973.760 5.940 973.960 6.140 ;
  LAYER VI3 ;
  RECT 973.360 6.340 973.560 6.540 ;
  LAYER VI3 ;
  RECT 973.360 5.940 973.560 6.140 ;
  LAYER VI3 ;
  RECT 972.960 6.340 973.160 6.540 ;
  LAYER VI3 ;
  RECT 972.960 5.940 973.160 6.140 ;
  LAYER VI3 ;
  RECT 972.560 6.340 972.760 6.540 ;
  LAYER VI3 ;
  RECT 972.560 5.940 972.760 6.140 ;
  LAYER VI3 ;
  RECT 972.160 6.340 972.360 6.540 ;
  LAYER VI3 ;
  RECT 972.160 5.940 972.360 6.140 ;
  LAYER VI3 ;
  RECT 971.760 6.340 971.960 6.540 ;
  LAYER VI3 ;
  RECT 971.760 5.940 971.960 6.140 ;
  LAYER VI3 ;
  RECT 971.360 6.340 971.560 6.540 ;
  LAYER VI3 ;
  RECT 971.360 5.940 971.560 6.140 ;
  LAYER VI3 ;
  RECT 970.960 6.340 971.160 6.540 ;
  LAYER VI3 ;
  RECT 970.960 5.940 971.160 6.140 ;
  LAYER VI3 ;
  RECT 970.560 6.340 970.760 6.540 ;
  LAYER VI3 ;
  RECT 970.560 5.940 970.760 6.140 ;
  LAYER VI3 ;
  RECT 970.160 6.340 970.360 6.540 ;
  LAYER VI3 ;
  RECT 970.160 5.940 970.360 6.140 ;
  LAYER VI3 ;
  RECT 969.760 6.340 969.960 6.540 ;
  LAYER VI3 ;
  RECT 969.760 5.940 969.960 6.140 ;
  LAYER VI3 ;
  RECT 969.360 6.340 969.560 6.540 ;
  LAYER VI3 ;
  RECT 969.360 5.940 969.560 6.140 ;
  LAYER VI3 ;
  RECT 990.440 5.880 998.440 6.740 ;
  LAYER VI3 ;
  RECT 998.040 6.340 998.240 6.540 ;
  LAYER VI3 ;
  RECT 998.040 5.940 998.240 6.140 ;
  LAYER VI3 ;
  RECT 997.640 6.340 997.840 6.540 ;
  LAYER VI3 ;
  RECT 997.640 5.940 997.840 6.140 ;
  LAYER VI3 ;
  RECT 997.240 6.340 997.440 6.540 ;
  LAYER VI3 ;
  RECT 997.240 5.940 997.440 6.140 ;
  LAYER VI3 ;
  RECT 996.840 6.340 997.040 6.540 ;
  LAYER VI3 ;
  RECT 996.840 5.940 997.040 6.140 ;
  LAYER VI3 ;
  RECT 996.440 6.340 996.640 6.540 ;
  LAYER VI3 ;
  RECT 996.440 5.940 996.640 6.140 ;
  LAYER VI3 ;
  RECT 996.040 6.340 996.240 6.540 ;
  LAYER VI3 ;
  RECT 996.040 5.940 996.240 6.140 ;
  LAYER VI3 ;
  RECT 995.640 6.340 995.840 6.540 ;
  LAYER VI3 ;
  RECT 995.640 5.940 995.840 6.140 ;
  LAYER VI3 ;
  RECT 995.240 6.340 995.440 6.540 ;
  LAYER VI3 ;
  RECT 995.240 5.940 995.440 6.140 ;
  LAYER VI3 ;
  RECT 994.840 6.340 995.040 6.540 ;
  LAYER VI3 ;
  RECT 994.840 5.940 995.040 6.140 ;
  LAYER VI3 ;
  RECT 994.440 6.340 994.640 6.540 ;
  LAYER VI3 ;
  RECT 994.440 5.940 994.640 6.140 ;
  LAYER VI3 ;
  RECT 994.040 6.340 994.240 6.540 ;
  LAYER VI3 ;
  RECT 994.040 5.940 994.240 6.140 ;
  LAYER VI3 ;
  RECT 993.640 6.340 993.840 6.540 ;
  LAYER VI3 ;
  RECT 993.640 5.940 993.840 6.140 ;
  LAYER VI3 ;
  RECT 993.240 6.340 993.440 6.540 ;
  LAYER VI3 ;
  RECT 993.240 5.940 993.440 6.140 ;
  LAYER VI3 ;
  RECT 992.840 6.340 993.040 6.540 ;
  LAYER VI3 ;
  RECT 992.840 5.940 993.040 6.140 ;
  LAYER VI3 ;
  RECT 992.440 6.340 992.640 6.540 ;
  LAYER VI3 ;
  RECT 992.440 5.940 992.640 6.140 ;
  LAYER VI3 ;
  RECT 992.040 6.340 992.240 6.540 ;
  LAYER VI3 ;
  RECT 992.040 5.940 992.240 6.140 ;
  LAYER VI3 ;
  RECT 991.640 6.340 991.840 6.540 ;
  LAYER VI3 ;
  RECT 991.640 5.940 991.840 6.140 ;
  LAYER VI3 ;
  RECT 991.240 6.340 991.440 6.540 ;
  LAYER VI3 ;
  RECT 991.240 5.940 991.440 6.140 ;
  LAYER VI3 ;
  RECT 990.840 6.340 991.040 6.540 ;
  LAYER VI3 ;
  RECT 990.840 5.940 991.040 6.140 ;
  LAYER VI3 ;
  RECT 990.440 6.340 990.640 6.540 ;
  LAYER VI3 ;
  RECT 990.440 5.940 990.640 6.140 ;
  LAYER VI3 ;
  RECT 1010.280 5.880 1018.280 6.740 ;
  LAYER VI3 ;
  RECT 1017.880 6.340 1018.080 6.540 ;
  LAYER VI3 ;
  RECT 1017.880 5.940 1018.080 6.140 ;
  LAYER VI3 ;
  RECT 1017.480 6.340 1017.680 6.540 ;
  LAYER VI3 ;
  RECT 1017.480 5.940 1017.680 6.140 ;
  LAYER VI3 ;
  RECT 1017.080 6.340 1017.280 6.540 ;
  LAYER VI3 ;
  RECT 1017.080 5.940 1017.280 6.140 ;
  LAYER VI3 ;
  RECT 1016.680 6.340 1016.880 6.540 ;
  LAYER VI3 ;
  RECT 1016.680 5.940 1016.880 6.140 ;
  LAYER VI3 ;
  RECT 1016.280 6.340 1016.480 6.540 ;
  LAYER VI3 ;
  RECT 1016.280 5.940 1016.480 6.140 ;
  LAYER VI3 ;
  RECT 1015.880 6.340 1016.080 6.540 ;
  LAYER VI3 ;
  RECT 1015.880 5.940 1016.080 6.140 ;
  LAYER VI3 ;
  RECT 1015.480 6.340 1015.680 6.540 ;
  LAYER VI3 ;
  RECT 1015.480 5.940 1015.680 6.140 ;
  LAYER VI3 ;
  RECT 1015.080 6.340 1015.280 6.540 ;
  LAYER VI3 ;
  RECT 1015.080 5.940 1015.280 6.140 ;
  LAYER VI3 ;
  RECT 1014.680 6.340 1014.880 6.540 ;
  LAYER VI3 ;
  RECT 1014.680 5.940 1014.880 6.140 ;
  LAYER VI3 ;
  RECT 1014.280 6.340 1014.480 6.540 ;
  LAYER VI3 ;
  RECT 1014.280 5.940 1014.480 6.140 ;
  LAYER VI3 ;
  RECT 1013.880 6.340 1014.080 6.540 ;
  LAYER VI3 ;
  RECT 1013.880 5.940 1014.080 6.140 ;
  LAYER VI3 ;
  RECT 1013.480 6.340 1013.680 6.540 ;
  LAYER VI3 ;
  RECT 1013.480 5.940 1013.680 6.140 ;
  LAYER VI3 ;
  RECT 1013.080 6.340 1013.280 6.540 ;
  LAYER VI3 ;
  RECT 1013.080 5.940 1013.280 6.140 ;
  LAYER VI3 ;
  RECT 1012.680 6.340 1012.880 6.540 ;
  LAYER VI3 ;
  RECT 1012.680 5.940 1012.880 6.140 ;
  LAYER VI3 ;
  RECT 1012.280 6.340 1012.480 6.540 ;
  LAYER VI3 ;
  RECT 1012.280 5.940 1012.480 6.140 ;
  LAYER VI3 ;
  RECT 1011.880 6.340 1012.080 6.540 ;
  LAYER VI3 ;
  RECT 1011.880 5.940 1012.080 6.140 ;
  LAYER VI3 ;
  RECT 1011.480 6.340 1011.680 6.540 ;
  LAYER VI3 ;
  RECT 1011.480 5.940 1011.680 6.140 ;
  LAYER VI3 ;
  RECT 1011.080 6.340 1011.280 6.540 ;
  LAYER VI3 ;
  RECT 1011.080 5.940 1011.280 6.140 ;
  LAYER VI3 ;
  RECT 1010.680 6.340 1010.880 6.540 ;
  LAYER VI3 ;
  RECT 1010.680 5.940 1010.880 6.140 ;
  LAYER VI3 ;
  RECT 1010.280 6.340 1010.480 6.540 ;
  LAYER VI3 ;
  RECT 1010.280 5.940 1010.480 6.140 ;
  LAYER VI3 ;
  RECT 1031.360 5.880 1039.360 6.740 ;
  LAYER VI3 ;
  RECT 1038.960 6.340 1039.160 6.540 ;
  LAYER VI3 ;
  RECT 1038.960 5.940 1039.160 6.140 ;
  LAYER VI3 ;
  RECT 1038.560 6.340 1038.760 6.540 ;
  LAYER VI3 ;
  RECT 1038.560 5.940 1038.760 6.140 ;
  LAYER VI3 ;
  RECT 1038.160 6.340 1038.360 6.540 ;
  LAYER VI3 ;
  RECT 1038.160 5.940 1038.360 6.140 ;
  LAYER VI3 ;
  RECT 1037.760 6.340 1037.960 6.540 ;
  LAYER VI3 ;
  RECT 1037.760 5.940 1037.960 6.140 ;
  LAYER VI3 ;
  RECT 1037.360 6.340 1037.560 6.540 ;
  LAYER VI3 ;
  RECT 1037.360 5.940 1037.560 6.140 ;
  LAYER VI3 ;
  RECT 1036.960 6.340 1037.160 6.540 ;
  LAYER VI3 ;
  RECT 1036.960 5.940 1037.160 6.140 ;
  LAYER VI3 ;
  RECT 1036.560 6.340 1036.760 6.540 ;
  LAYER VI3 ;
  RECT 1036.560 5.940 1036.760 6.140 ;
  LAYER VI3 ;
  RECT 1036.160 6.340 1036.360 6.540 ;
  LAYER VI3 ;
  RECT 1036.160 5.940 1036.360 6.140 ;
  LAYER VI3 ;
  RECT 1035.760 6.340 1035.960 6.540 ;
  LAYER VI3 ;
  RECT 1035.760 5.940 1035.960 6.140 ;
  LAYER VI3 ;
  RECT 1035.360 6.340 1035.560 6.540 ;
  LAYER VI3 ;
  RECT 1035.360 5.940 1035.560 6.140 ;
  LAYER VI3 ;
  RECT 1034.960 6.340 1035.160 6.540 ;
  LAYER VI3 ;
  RECT 1034.960 5.940 1035.160 6.140 ;
  LAYER VI3 ;
  RECT 1034.560 6.340 1034.760 6.540 ;
  LAYER VI3 ;
  RECT 1034.560 5.940 1034.760 6.140 ;
  LAYER VI3 ;
  RECT 1034.160 6.340 1034.360 6.540 ;
  LAYER VI3 ;
  RECT 1034.160 5.940 1034.360 6.140 ;
  LAYER VI3 ;
  RECT 1033.760 6.340 1033.960 6.540 ;
  LAYER VI3 ;
  RECT 1033.760 5.940 1033.960 6.140 ;
  LAYER VI3 ;
  RECT 1033.360 6.340 1033.560 6.540 ;
  LAYER VI3 ;
  RECT 1033.360 5.940 1033.560 6.140 ;
  LAYER VI3 ;
  RECT 1032.960 6.340 1033.160 6.540 ;
  LAYER VI3 ;
  RECT 1032.960 5.940 1033.160 6.140 ;
  LAYER VI3 ;
  RECT 1032.560 6.340 1032.760 6.540 ;
  LAYER VI3 ;
  RECT 1032.560 5.940 1032.760 6.140 ;
  LAYER VI3 ;
  RECT 1032.160 6.340 1032.360 6.540 ;
  LAYER VI3 ;
  RECT 1032.160 5.940 1032.360 6.140 ;
  LAYER VI3 ;
  RECT 1031.760 6.340 1031.960 6.540 ;
  LAYER VI3 ;
  RECT 1031.760 5.940 1031.960 6.140 ;
  LAYER VI3 ;
  RECT 1031.360 6.340 1031.560 6.540 ;
  LAYER VI3 ;
  RECT 1031.360 5.940 1031.560 6.140 ;
  LAYER VI3 ;
  RECT 1051.200 5.880 1059.200 6.740 ;
  LAYER VI3 ;
  RECT 1058.800 6.340 1059.000 6.540 ;
  LAYER VI3 ;
  RECT 1058.800 5.940 1059.000 6.140 ;
  LAYER VI3 ;
  RECT 1058.400 6.340 1058.600 6.540 ;
  LAYER VI3 ;
  RECT 1058.400 5.940 1058.600 6.140 ;
  LAYER VI3 ;
  RECT 1058.000 6.340 1058.200 6.540 ;
  LAYER VI3 ;
  RECT 1058.000 5.940 1058.200 6.140 ;
  LAYER VI3 ;
  RECT 1057.600 6.340 1057.800 6.540 ;
  LAYER VI3 ;
  RECT 1057.600 5.940 1057.800 6.140 ;
  LAYER VI3 ;
  RECT 1057.200 6.340 1057.400 6.540 ;
  LAYER VI3 ;
  RECT 1057.200 5.940 1057.400 6.140 ;
  LAYER VI3 ;
  RECT 1056.800 6.340 1057.000 6.540 ;
  LAYER VI3 ;
  RECT 1056.800 5.940 1057.000 6.140 ;
  LAYER VI3 ;
  RECT 1056.400 6.340 1056.600 6.540 ;
  LAYER VI3 ;
  RECT 1056.400 5.940 1056.600 6.140 ;
  LAYER VI3 ;
  RECT 1056.000 6.340 1056.200 6.540 ;
  LAYER VI3 ;
  RECT 1056.000 5.940 1056.200 6.140 ;
  LAYER VI3 ;
  RECT 1055.600 6.340 1055.800 6.540 ;
  LAYER VI3 ;
  RECT 1055.600 5.940 1055.800 6.140 ;
  LAYER VI3 ;
  RECT 1055.200 6.340 1055.400 6.540 ;
  LAYER VI3 ;
  RECT 1055.200 5.940 1055.400 6.140 ;
  LAYER VI3 ;
  RECT 1054.800 6.340 1055.000 6.540 ;
  LAYER VI3 ;
  RECT 1054.800 5.940 1055.000 6.140 ;
  LAYER VI3 ;
  RECT 1054.400 6.340 1054.600 6.540 ;
  LAYER VI3 ;
  RECT 1054.400 5.940 1054.600 6.140 ;
  LAYER VI3 ;
  RECT 1054.000 6.340 1054.200 6.540 ;
  LAYER VI3 ;
  RECT 1054.000 5.940 1054.200 6.140 ;
  LAYER VI3 ;
  RECT 1053.600 6.340 1053.800 6.540 ;
  LAYER VI3 ;
  RECT 1053.600 5.940 1053.800 6.140 ;
  LAYER VI3 ;
  RECT 1053.200 6.340 1053.400 6.540 ;
  LAYER VI3 ;
  RECT 1053.200 5.940 1053.400 6.140 ;
  LAYER VI3 ;
  RECT 1052.800 6.340 1053.000 6.540 ;
  LAYER VI3 ;
  RECT 1052.800 5.940 1053.000 6.140 ;
  LAYER VI3 ;
  RECT 1052.400 6.340 1052.600 6.540 ;
  LAYER VI3 ;
  RECT 1052.400 5.940 1052.600 6.140 ;
  LAYER VI3 ;
  RECT 1052.000 6.340 1052.200 6.540 ;
  LAYER VI3 ;
  RECT 1052.000 5.940 1052.200 6.140 ;
  LAYER VI3 ;
  RECT 1051.600 6.340 1051.800 6.540 ;
  LAYER VI3 ;
  RECT 1051.600 5.940 1051.800 6.140 ;
  LAYER VI3 ;
  RECT 1051.200 6.340 1051.400 6.540 ;
  LAYER VI3 ;
  RECT 1051.200 5.940 1051.400 6.140 ;
  LAYER VI3 ;
  RECT 1072.280 5.880 1080.280 6.740 ;
  LAYER VI3 ;
  RECT 1079.880 6.340 1080.080 6.540 ;
  LAYER VI3 ;
  RECT 1079.880 5.940 1080.080 6.140 ;
  LAYER VI3 ;
  RECT 1079.480 6.340 1079.680 6.540 ;
  LAYER VI3 ;
  RECT 1079.480 5.940 1079.680 6.140 ;
  LAYER VI3 ;
  RECT 1079.080 6.340 1079.280 6.540 ;
  LAYER VI3 ;
  RECT 1079.080 5.940 1079.280 6.140 ;
  LAYER VI3 ;
  RECT 1078.680 6.340 1078.880 6.540 ;
  LAYER VI3 ;
  RECT 1078.680 5.940 1078.880 6.140 ;
  LAYER VI3 ;
  RECT 1078.280 6.340 1078.480 6.540 ;
  LAYER VI3 ;
  RECT 1078.280 5.940 1078.480 6.140 ;
  LAYER VI3 ;
  RECT 1077.880 6.340 1078.080 6.540 ;
  LAYER VI3 ;
  RECT 1077.880 5.940 1078.080 6.140 ;
  LAYER VI3 ;
  RECT 1077.480 6.340 1077.680 6.540 ;
  LAYER VI3 ;
  RECT 1077.480 5.940 1077.680 6.140 ;
  LAYER VI3 ;
  RECT 1077.080 6.340 1077.280 6.540 ;
  LAYER VI3 ;
  RECT 1077.080 5.940 1077.280 6.140 ;
  LAYER VI3 ;
  RECT 1076.680 6.340 1076.880 6.540 ;
  LAYER VI3 ;
  RECT 1076.680 5.940 1076.880 6.140 ;
  LAYER VI3 ;
  RECT 1076.280 6.340 1076.480 6.540 ;
  LAYER VI3 ;
  RECT 1076.280 5.940 1076.480 6.140 ;
  LAYER VI3 ;
  RECT 1075.880 6.340 1076.080 6.540 ;
  LAYER VI3 ;
  RECT 1075.880 5.940 1076.080 6.140 ;
  LAYER VI3 ;
  RECT 1075.480 6.340 1075.680 6.540 ;
  LAYER VI3 ;
  RECT 1075.480 5.940 1075.680 6.140 ;
  LAYER VI3 ;
  RECT 1075.080 6.340 1075.280 6.540 ;
  LAYER VI3 ;
  RECT 1075.080 5.940 1075.280 6.140 ;
  LAYER VI3 ;
  RECT 1074.680 6.340 1074.880 6.540 ;
  LAYER VI3 ;
  RECT 1074.680 5.940 1074.880 6.140 ;
  LAYER VI3 ;
  RECT 1074.280 6.340 1074.480 6.540 ;
  LAYER VI3 ;
  RECT 1074.280 5.940 1074.480 6.140 ;
  LAYER VI3 ;
  RECT 1073.880 6.340 1074.080 6.540 ;
  LAYER VI3 ;
  RECT 1073.880 5.940 1074.080 6.140 ;
  LAYER VI3 ;
  RECT 1073.480 6.340 1073.680 6.540 ;
  LAYER VI3 ;
  RECT 1073.480 5.940 1073.680 6.140 ;
  LAYER VI3 ;
  RECT 1073.080 6.340 1073.280 6.540 ;
  LAYER VI3 ;
  RECT 1073.080 5.940 1073.280 6.140 ;
  LAYER VI3 ;
  RECT 1072.680 6.340 1072.880 6.540 ;
  LAYER VI3 ;
  RECT 1072.680 5.940 1072.880 6.140 ;
  LAYER VI3 ;
  RECT 1072.280 6.340 1072.480 6.540 ;
  LAYER VI3 ;
  RECT 1072.280 5.940 1072.480 6.140 ;
  LAYER VI3 ;
  RECT 1092.120 5.880 1100.120 6.740 ;
  LAYER VI3 ;
  RECT 1099.720 6.340 1099.920 6.540 ;
  LAYER VI3 ;
  RECT 1099.720 5.940 1099.920 6.140 ;
  LAYER VI3 ;
  RECT 1099.320 6.340 1099.520 6.540 ;
  LAYER VI3 ;
  RECT 1099.320 5.940 1099.520 6.140 ;
  LAYER VI3 ;
  RECT 1098.920 6.340 1099.120 6.540 ;
  LAYER VI3 ;
  RECT 1098.920 5.940 1099.120 6.140 ;
  LAYER VI3 ;
  RECT 1098.520 6.340 1098.720 6.540 ;
  LAYER VI3 ;
  RECT 1098.520 5.940 1098.720 6.140 ;
  LAYER VI3 ;
  RECT 1098.120 6.340 1098.320 6.540 ;
  LAYER VI3 ;
  RECT 1098.120 5.940 1098.320 6.140 ;
  LAYER VI3 ;
  RECT 1097.720 6.340 1097.920 6.540 ;
  LAYER VI3 ;
  RECT 1097.720 5.940 1097.920 6.140 ;
  LAYER VI3 ;
  RECT 1097.320 6.340 1097.520 6.540 ;
  LAYER VI3 ;
  RECT 1097.320 5.940 1097.520 6.140 ;
  LAYER VI3 ;
  RECT 1096.920 6.340 1097.120 6.540 ;
  LAYER VI3 ;
  RECT 1096.920 5.940 1097.120 6.140 ;
  LAYER VI3 ;
  RECT 1096.520 6.340 1096.720 6.540 ;
  LAYER VI3 ;
  RECT 1096.520 5.940 1096.720 6.140 ;
  LAYER VI3 ;
  RECT 1096.120 6.340 1096.320 6.540 ;
  LAYER VI3 ;
  RECT 1096.120 5.940 1096.320 6.140 ;
  LAYER VI3 ;
  RECT 1095.720 6.340 1095.920 6.540 ;
  LAYER VI3 ;
  RECT 1095.720 5.940 1095.920 6.140 ;
  LAYER VI3 ;
  RECT 1095.320 6.340 1095.520 6.540 ;
  LAYER VI3 ;
  RECT 1095.320 5.940 1095.520 6.140 ;
  LAYER VI3 ;
  RECT 1094.920 6.340 1095.120 6.540 ;
  LAYER VI3 ;
  RECT 1094.920 5.940 1095.120 6.140 ;
  LAYER VI3 ;
  RECT 1094.520 6.340 1094.720 6.540 ;
  LAYER VI3 ;
  RECT 1094.520 5.940 1094.720 6.140 ;
  LAYER VI3 ;
  RECT 1094.120 6.340 1094.320 6.540 ;
  LAYER VI3 ;
  RECT 1094.120 5.940 1094.320 6.140 ;
  LAYER VI3 ;
  RECT 1093.720 6.340 1093.920 6.540 ;
  LAYER VI3 ;
  RECT 1093.720 5.940 1093.920 6.140 ;
  LAYER VI3 ;
  RECT 1093.320 6.340 1093.520 6.540 ;
  LAYER VI3 ;
  RECT 1093.320 5.940 1093.520 6.140 ;
  LAYER VI3 ;
  RECT 1092.920 6.340 1093.120 6.540 ;
  LAYER VI3 ;
  RECT 1092.920 5.940 1093.120 6.140 ;
  LAYER VI3 ;
  RECT 1092.520 6.340 1092.720 6.540 ;
  LAYER VI3 ;
  RECT 1092.520 5.940 1092.720 6.140 ;
  LAYER VI3 ;
  RECT 1092.120 6.340 1092.320 6.540 ;
  LAYER VI3 ;
  RECT 1092.120 5.940 1092.320 6.140 ;
  LAYER VI3 ;
  RECT 1113.200 5.880 1121.200 6.740 ;
  LAYER VI3 ;
  RECT 1120.800 6.340 1121.000 6.540 ;
  LAYER VI3 ;
  RECT 1120.800 5.940 1121.000 6.140 ;
  LAYER VI3 ;
  RECT 1120.400 6.340 1120.600 6.540 ;
  LAYER VI3 ;
  RECT 1120.400 5.940 1120.600 6.140 ;
  LAYER VI3 ;
  RECT 1120.000 6.340 1120.200 6.540 ;
  LAYER VI3 ;
  RECT 1120.000 5.940 1120.200 6.140 ;
  LAYER VI3 ;
  RECT 1119.600 6.340 1119.800 6.540 ;
  LAYER VI3 ;
  RECT 1119.600 5.940 1119.800 6.140 ;
  LAYER VI3 ;
  RECT 1119.200 6.340 1119.400 6.540 ;
  LAYER VI3 ;
  RECT 1119.200 5.940 1119.400 6.140 ;
  LAYER VI3 ;
  RECT 1118.800 6.340 1119.000 6.540 ;
  LAYER VI3 ;
  RECT 1118.800 5.940 1119.000 6.140 ;
  LAYER VI3 ;
  RECT 1118.400 6.340 1118.600 6.540 ;
  LAYER VI3 ;
  RECT 1118.400 5.940 1118.600 6.140 ;
  LAYER VI3 ;
  RECT 1118.000 6.340 1118.200 6.540 ;
  LAYER VI3 ;
  RECT 1118.000 5.940 1118.200 6.140 ;
  LAYER VI3 ;
  RECT 1117.600 6.340 1117.800 6.540 ;
  LAYER VI3 ;
  RECT 1117.600 5.940 1117.800 6.140 ;
  LAYER VI3 ;
  RECT 1117.200 6.340 1117.400 6.540 ;
  LAYER VI3 ;
  RECT 1117.200 5.940 1117.400 6.140 ;
  LAYER VI3 ;
  RECT 1116.800 6.340 1117.000 6.540 ;
  LAYER VI3 ;
  RECT 1116.800 5.940 1117.000 6.140 ;
  LAYER VI3 ;
  RECT 1116.400 6.340 1116.600 6.540 ;
  LAYER VI3 ;
  RECT 1116.400 5.940 1116.600 6.140 ;
  LAYER VI3 ;
  RECT 1116.000 6.340 1116.200 6.540 ;
  LAYER VI3 ;
  RECT 1116.000 5.940 1116.200 6.140 ;
  LAYER VI3 ;
  RECT 1115.600 6.340 1115.800 6.540 ;
  LAYER VI3 ;
  RECT 1115.600 5.940 1115.800 6.140 ;
  LAYER VI3 ;
  RECT 1115.200 6.340 1115.400 6.540 ;
  LAYER VI3 ;
  RECT 1115.200 5.940 1115.400 6.140 ;
  LAYER VI3 ;
  RECT 1114.800 6.340 1115.000 6.540 ;
  LAYER VI3 ;
  RECT 1114.800 5.940 1115.000 6.140 ;
  LAYER VI3 ;
  RECT 1114.400 6.340 1114.600 6.540 ;
  LAYER VI3 ;
  RECT 1114.400 5.940 1114.600 6.140 ;
  LAYER VI3 ;
  RECT 1114.000 6.340 1114.200 6.540 ;
  LAYER VI3 ;
  RECT 1114.000 5.940 1114.200 6.140 ;
  LAYER VI3 ;
  RECT 1113.600 6.340 1113.800 6.540 ;
  LAYER VI3 ;
  RECT 1113.600 5.940 1113.800 6.140 ;
  LAYER VI3 ;
  RECT 1113.200 6.340 1113.400 6.540 ;
  LAYER VI3 ;
  RECT 1113.200 5.940 1113.400 6.140 ;
  LAYER VI3 ;
  RECT 1133.040 5.880 1141.040 6.740 ;
  LAYER VI3 ;
  RECT 1140.640 6.340 1140.840 6.540 ;
  LAYER VI3 ;
  RECT 1140.640 5.940 1140.840 6.140 ;
  LAYER VI3 ;
  RECT 1140.240 6.340 1140.440 6.540 ;
  LAYER VI3 ;
  RECT 1140.240 5.940 1140.440 6.140 ;
  LAYER VI3 ;
  RECT 1139.840 6.340 1140.040 6.540 ;
  LAYER VI3 ;
  RECT 1139.840 5.940 1140.040 6.140 ;
  LAYER VI3 ;
  RECT 1139.440 6.340 1139.640 6.540 ;
  LAYER VI3 ;
  RECT 1139.440 5.940 1139.640 6.140 ;
  LAYER VI3 ;
  RECT 1139.040 6.340 1139.240 6.540 ;
  LAYER VI3 ;
  RECT 1139.040 5.940 1139.240 6.140 ;
  LAYER VI3 ;
  RECT 1138.640 6.340 1138.840 6.540 ;
  LAYER VI3 ;
  RECT 1138.640 5.940 1138.840 6.140 ;
  LAYER VI3 ;
  RECT 1138.240 6.340 1138.440 6.540 ;
  LAYER VI3 ;
  RECT 1138.240 5.940 1138.440 6.140 ;
  LAYER VI3 ;
  RECT 1137.840 6.340 1138.040 6.540 ;
  LAYER VI3 ;
  RECT 1137.840 5.940 1138.040 6.140 ;
  LAYER VI3 ;
  RECT 1137.440 6.340 1137.640 6.540 ;
  LAYER VI3 ;
  RECT 1137.440 5.940 1137.640 6.140 ;
  LAYER VI3 ;
  RECT 1137.040 6.340 1137.240 6.540 ;
  LAYER VI3 ;
  RECT 1137.040 5.940 1137.240 6.140 ;
  LAYER VI3 ;
  RECT 1136.640 6.340 1136.840 6.540 ;
  LAYER VI3 ;
  RECT 1136.640 5.940 1136.840 6.140 ;
  LAYER VI3 ;
  RECT 1136.240 6.340 1136.440 6.540 ;
  LAYER VI3 ;
  RECT 1136.240 5.940 1136.440 6.140 ;
  LAYER VI3 ;
  RECT 1135.840 6.340 1136.040 6.540 ;
  LAYER VI3 ;
  RECT 1135.840 5.940 1136.040 6.140 ;
  LAYER VI3 ;
  RECT 1135.440 6.340 1135.640 6.540 ;
  LAYER VI3 ;
  RECT 1135.440 5.940 1135.640 6.140 ;
  LAYER VI3 ;
  RECT 1135.040 6.340 1135.240 6.540 ;
  LAYER VI3 ;
  RECT 1135.040 5.940 1135.240 6.140 ;
  LAYER VI3 ;
  RECT 1134.640 6.340 1134.840 6.540 ;
  LAYER VI3 ;
  RECT 1134.640 5.940 1134.840 6.140 ;
  LAYER VI3 ;
  RECT 1134.240 6.340 1134.440 6.540 ;
  LAYER VI3 ;
  RECT 1134.240 5.940 1134.440 6.140 ;
  LAYER VI3 ;
  RECT 1133.840 6.340 1134.040 6.540 ;
  LAYER VI3 ;
  RECT 1133.840 5.940 1134.040 6.140 ;
  LAYER VI3 ;
  RECT 1133.440 6.340 1133.640 6.540 ;
  LAYER VI3 ;
  RECT 1133.440 5.940 1133.640 6.140 ;
  LAYER VI3 ;
  RECT 1133.040 6.340 1133.240 6.540 ;
  LAYER VI3 ;
  RECT 1133.040 5.940 1133.240 6.140 ;
  LAYER VI3 ;
  RECT 1154.120 5.880 1162.120 6.740 ;
  LAYER VI3 ;
  RECT 1161.720 6.340 1161.920 6.540 ;
  LAYER VI3 ;
  RECT 1161.720 5.940 1161.920 6.140 ;
  LAYER VI3 ;
  RECT 1161.320 6.340 1161.520 6.540 ;
  LAYER VI3 ;
  RECT 1161.320 5.940 1161.520 6.140 ;
  LAYER VI3 ;
  RECT 1160.920 6.340 1161.120 6.540 ;
  LAYER VI3 ;
  RECT 1160.920 5.940 1161.120 6.140 ;
  LAYER VI3 ;
  RECT 1160.520 6.340 1160.720 6.540 ;
  LAYER VI3 ;
  RECT 1160.520 5.940 1160.720 6.140 ;
  LAYER VI3 ;
  RECT 1160.120 6.340 1160.320 6.540 ;
  LAYER VI3 ;
  RECT 1160.120 5.940 1160.320 6.140 ;
  LAYER VI3 ;
  RECT 1159.720 6.340 1159.920 6.540 ;
  LAYER VI3 ;
  RECT 1159.720 5.940 1159.920 6.140 ;
  LAYER VI3 ;
  RECT 1159.320 6.340 1159.520 6.540 ;
  LAYER VI3 ;
  RECT 1159.320 5.940 1159.520 6.140 ;
  LAYER VI3 ;
  RECT 1158.920 6.340 1159.120 6.540 ;
  LAYER VI3 ;
  RECT 1158.920 5.940 1159.120 6.140 ;
  LAYER VI3 ;
  RECT 1158.520 6.340 1158.720 6.540 ;
  LAYER VI3 ;
  RECT 1158.520 5.940 1158.720 6.140 ;
  LAYER VI3 ;
  RECT 1158.120 6.340 1158.320 6.540 ;
  LAYER VI3 ;
  RECT 1158.120 5.940 1158.320 6.140 ;
  LAYER VI3 ;
  RECT 1157.720 6.340 1157.920 6.540 ;
  LAYER VI3 ;
  RECT 1157.720 5.940 1157.920 6.140 ;
  LAYER VI3 ;
  RECT 1157.320 6.340 1157.520 6.540 ;
  LAYER VI3 ;
  RECT 1157.320 5.940 1157.520 6.140 ;
  LAYER VI3 ;
  RECT 1156.920 6.340 1157.120 6.540 ;
  LAYER VI3 ;
  RECT 1156.920 5.940 1157.120 6.140 ;
  LAYER VI3 ;
  RECT 1156.520 6.340 1156.720 6.540 ;
  LAYER VI3 ;
  RECT 1156.520 5.940 1156.720 6.140 ;
  LAYER VI3 ;
  RECT 1156.120 6.340 1156.320 6.540 ;
  LAYER VI3 ;
  RECT 1156.120 5.940 1156.320 6.140 ;
  LAYER VI3 ;
  RECT 1155.720 6.340 1155.920 6.540 ;
  LAYER VI3 ;
  RECT 1155.720 5.940 1155.920 6.140 ;
  LAYER VI3 ;
  RECT 1155.320 6.340 1155.520 6.540 ;
  LAYER VI3 ;
  RECT 1155.320 5.940 1155.520 6.140 ;
  LAYER VI3 ;
  RECT 1154.920 6.340 1155.120 6.540 ;
  LAYER VI3 ;
  RECT 1154.920 5.940 1155.120 6.140 ;
  LAYER VI3 ;
  RECT 1154.520 6.340 1154.720 6.540 ;
  LAYER VI3 ;
  RECT 1154.520 5.940 1154.720 6.140 ;
  LAYER VI3 ;
  RECT 1154.120 6.340 1154.320 6.540 ;
  LAYER VI3 ;
  RECT 1154.120 5.940 1154.320 6.140 ;
  LAYER VI3 ;
  RECT 1173.960 5.880 1181.960 6.740 ;
  LAYER VI3 ;
  RECT 1181.560 6.340 1181.760 6.540 ;
  LAYER VI3 ;
  RECT 1181.560 5.940 1181.760 6.140 ;
  LAYER VI3 ;
  RECT 1181.160 6.340 1181.360 6.540 ;
  LAYER VI3 ;
  RECT 1181.160 5.940 1181.360 6.140 ;
  LAYER VI3 ;
  RECT 1180.760 6.340 1180.960 6.540 ;
  LAYER VI3 ;
  RECT 1180.760 5.940 1180.960 6.140 ;
  LAYER VI3 ;
  RECT 1180.360 6.340 1180.560 6.540 ;
  LAYER VI3 ;
  RECT 1180.360 5.940 1180.560 6.140 ;
  LAYER VI3 ;
  RECT 1179.960 6.340 1180.160 6.540 ;
  LAYER VI3 ;
  RECT 1179.960 5.940 1180.160 6.140 ;
  LAYER VI3 ;
  RECT 1179.560 6.340 1179.760 6.540 ;
  LAYER VI3 ;
  RECT 1179.560 5.940 1179.760 6.140 ;
  LAYER VI3 ;
  RECT 1179.160 6.340 1179.360 6.540 ;
  LAYER VI3 ;
  RECT 1179.160 5.940 1179.360 6.140 ;
  LAYER VI3 ;
  RECT 1178.760 6.340 1178.960 6.540 ;
  LAYER VI3 ;
  RECT 1178.760 5.940 1178.960 6.140 ;
  LAYER VI3 ;
  RECT 1178.360 6.340 1178.560 6.540 ;
  LAYER VI3 ;
  RECT 1178.360 5.940 1178.560 6.140 ;
  LAYER VI3 ;
  RECT 1177.960 6.340 1178.160 6.540 ;
  LAYER VI3 ;
  RECT 1177.960 5.940 1178.160 6.140 ;
  LAYER VI3 ;
  RECT 1177.560 6.340 1177.760 6.540 ;
  LAYER VI3 ;
  RECT 1177.560 5.940 1177.760 6.140 ;
  LAYER VI3 ;
  RECT 1177.160 6.340 1177.360 6.540 ;
  LAYER VI3 ;
  RECT 1177.160 5.940 1177.360 6.140 ;
  LAYER VI3 ;
  RECT 1176.760 6.340 1176.960 6.540 ;
  LAYER VI3 ;
  RECT 1176.760 5.940 1176.960 6.140 ;
  LAYER VI3 ;
  RECT 1176.360 6.340 1176.560 6.540 ;
  LAYER VI3 ;
  RECT 1176.360 5.940 1176.560 6.140 ;
  LAYER VI3 ;
  RECT 1175.960 6.340 1176.160 6.540 ;
  LAYER VI3 ;
  RECT 1175.960 5.940 1176.160 6.140 ;
  LAYER VI3 ;
  RECT 1175.560 6.340 1175.760 6.540 ;
  LAYER VI3 ;
  RECT 1175.560 5.940 1175.760 6.140 ;
  LAYER VI3 ;
  RECT 1175.160 6.340 1175.360 6.540 ;
  LAYER VI3 ;
  RECT 1175.160 5.940 1175.360 6.140 ;
  LAYER VI3 ;
  RECT 1174.760 6.340 1174.960 6.540 ;
  LAYER VI3 ;
  RECT 1174.760 5.940 1174.960 6.140 ;
  LAYER VI3 ;
  RECT 1174.360 6.340 1174.560 6.540 ;
  LAYER VI3 ;
  RECT 1174.360 5.940 1174.560 6.140 ;
  LAYER VI3 ;
  RECT 1173.960 6.340 1174.160 6.540 ;
  LAYER VI3 ;
  RECT 1173.960 5.940 1174.160 6.140 ;
  LAYER VI3 ;
  RECT 1195.040 5.880 1203.040 6.740 ;
  LAYER VI3 ;
  RECT 1202.640 6.340 1202.840 6.540 ;
  LAYER VI3 ;
  RECT 1202.640 5.940 1202.840 6.140 ;
  LAYER VI3 ;
  RECT 1202.240 6.340 1202.440 6.540 ;
  LAYER VI3 ;
  RECT 1202.240 5.940 1202.440 6.140 ;
  LAYER VI3 ;
  RECT 1201.840 6.340 1202.040 6.540 ;
  LAYER VI3 ;
  RECT 1201.840 5.940 1202.040 6.140 ;
  LAYER VI3 ;
  RECT 1201.440 6.340 1201.640 6.540 ;
  LAYER VI3 ;
  RECT 1201.440 5.940 1201.640 6.140 ;
  LAYER VI3 ;
  RECT 1201.040 6.340 1201.240 6.540 ;
  LAYER VI3 ;
  RECT 1201.040 5.940 1201.240 6.140 ;
  LAYER VI3 ;
  RECT 1200.640 6.340 1200.840 6.540 ;
  LAYER VI3 ;
  RECT 1200.640 5.940 1200.840 6.140 ;
  LAYER VI3 ;
  RECT 1200.240 6.340 1200.440 6.540 ;
  LAYER VI3 ;
  RECT 1200.240 5.940 1200.440 6.140 ;
  LAYER VI3 ;
  RECT 1199.840 6.340 1200.040 6.540 ;
  LAYER VI3 ;
  RECT 1199.840 5.940 1200.040 6.140 ;
  LAYER VI3 ;
  RECT 1199.440 6.340 1199.640 6.540 ;
  LAYER VI3 ;
  RECT 1199.440 5.940 1199.640 6.140 ;
  LAYER VI3 ;
  RECT 1199.040 6.340 1199.240 6.540 ;
  LAYER VI3 ;
  RECT 1199.040 5.940 1199.240 6.140 ;
  LAYER VI3 ;
  RECT 1198.640 6.340 1198.840 6.540 ;
  LAYER VI3 ;
  RECT 1198.640 5.940 1198.840 6.140 ;
  LAYER VI3 ;
  RECT 1198.240 6.340 1198.440 6.540 ;
  LAYER VI3 ;
  RECT 1198.240 5.940 1198.440 6.140 ;
  LAYER VI3 ;
  RECT 1197.840 6.340 1198.040 6.540 ;
  LAYER VI3 ;
  RECT 1197.840 5.940 1198.040 6.140 ;
  LAYER VI3 ;
  RECT 1197.440 6.340 1197.640 6.540 ;
  LAYER VI3 ;
  RECT 1197.440 5.940 1197.640 6.140 ;
  LAYER VI3 ;
  RECT 1197.040 6.340 1197.240 6.540 ;
  LAYER VI3 ;
  RECT 1197.040 5.940 1197.240 6.140 ;
  LAYER VI3 ;
  RECT 1196.640 6.340 1196.840 6.540 ;
  LAYER VI3 ;
  RECT 1196.640 5.940 1196.840 6.140 ;
  LAYER VI3 ;
  RECT 1196.240 6.340 1196.440 6.540 ;
  LAYER VI3 ;
  RECT 1196.240 5.940 1196.440 6.140 ;
  LAYER VI3 ;
  RECT 1195.840 6.340 1196.040 6.540 ;
  LAYER VI3 ;
  RECT 1195.840 5.940 1196.040 6.140 ;
  LAYER VI3 ;
  RECT 1195.440 6.340 1195.640 6.540 ;
  LAYER VI3 ;
  RECT 1195.440 5.940 1195.640 6.140 ;
  LAYER VI3 ;
  RECT 1195.040 6.340 1195.240 6.540 ;
  LAYER VI3 ;
  RECT 1195.040 5.940 1195.240 6.140 ;
  LAYER VI3 ;
  RECT 1214.880 5.880 1222.880 6.740 ;
  LAYER VI3 ;
  RECT 1222.480 6.340 1222.680 6.540 ;
  LAYER VI3 ;
  RECT 1222.480 5.940 1222.680 6.140 ;
  LAYER VI3 ;
  RECT 1222.080 6.340 1222.280 6.540 ;
  LAYER VI3 ;
  RECT 1222.080 5.940 1222.280 6.140 ;
  LAYER VI3 ;
  RECT 1221.680 6.340 1221.880 6.540 ;
  LAYER VI3 ;
  RECT 1221.680 5.940 1221.880 6.140 ;
  LAYER VI3 ;
  RECT 1221.280 6.340 1221.480 6.540 ;
  LAYER VI3 ;
  RECT 1221.280 5.940 1221.480 6.140 ;
  LAYER VI3 ;
  RECT 1220.880 6.340 1221.080 6.540 ;
  LAYER VI3 ;
  RECT 1220.880 5.940 1221.080 6.140 ;
  LAYER VI3 ;
  RECT 1220.480 6.340 1220.680 6.540 ;
  LAYER VI3 ;
  RECT 1220.480 5.940 1220.680 6.140 ;
  LAYER VI3 ;
  RECT 1220.080 6.340 1220.280 6.540 ;
  LAYER VI3 ;
  RECT 1220.080 5.940 1220.280 6.140 ;
  LAYER VI3 ;
  RECT 1219.680 6.340 1219.880 6.540 ;
  LAYER VI3 ;
  RECT 1219.680 5.940 1219.880 6.140 ;
  LAYER VI3 ;
  RECT 1219.280 6.340 1219.480 6.540 ;
  LAYER VI3 ;
  RECT 1219.280 5.940 1219.480 6.140 ;
  LAYER VI3 ;
  RECT 1218.880 6.340 1219.080 6.540 ;
  LAYER VI3 ;
  RECT 1218.880 5.940 1219.080 6.140 ;
  LAYER VI3 ;
  RECT 1218.480 6.340 1218.680 6.540 ;
  LAYER VI3 ;
  RECT 1218.480 5.940 1218.680 6.140 ;
  LAYER VI3 ;
  RECT 1218.080 6.340 1218.280 6.540 ;
  LAYER VI3 ;
  RECT 1218.080 5.940 1218.280 6.140 ;
  LAYER VI3 ;
  RECT 1217.680 6.340 1217.880 6.540 ;
  LAYER VI3 ;
  RECT 1217.680 5.940 1217.880 6.140 ;
  LAYER VI3 ;
  RECT 1217.280 6.340 1217.480 6.540 ;
  LAYER VI3 ;
  RECT 1217.280 5.940 1217.480 6.140 ;
  LAYER VI3 ;
  RECT 1216.880 6.340 1217.080 6.540 ;
  LAYER VI3 ;
  RECT 1216.880 5.940 1217.080 6.140 ;
  LAYER VI3 ;
  RECT 1216.480 6.340 1216.680 6.540 ;
  LAYER VI3 ;
  RECT 1216.480 5.940 1216.680 6.140 ;
  LAYER VI3 ;
  RECT 1216.080 6.340 1216.280 6.540 ;
  LAYER VI3 ;
  RECT 1216.080 5.940 1216.280 6.140 ;
  LAYER VI3 ;
  RECT 1215.680 6.340 1215.880 6.540 ;
  LAYER VI3 ;
  RECT 1215.680 5.940 1215.880 6.140 ;
  LAYER VI3 ;
  RECT 1215.280 6.340 1215.480 6.540 ;
  LAYER VI3 ;
  RECT 1215.280 5.940 1215.480 6.140 ;
  LAYER VI3 ;
  RECT 1214.880 6.340 1215.080 6.540 ;
  LAYER VI3 ;
  RECT 1214.880 5.940 1215.080 6.140 ;
  LAYER VI3 ;
  RECT 1235.960 5.880 1243.960 6.740 ;
  LAYER VI3 ;
  RECT 1243.560 6.340 1243.760 6.540 ;
  LAYER VI3 ;
  RECT 1243.560 5.940 1243.760 6.140 ;
  LAYER VI3 ;
  RECT 1243.160 6.340 1243.360 6.540 ;
  LAYER VI3 ;
  RECT 1243.160 5.940 1243.360 6.140 ;
  LAYER VI3 ;
  RECT 1242.760 6.340 1242.960 6.540 ;
  LAYER VI3 ;
  RECT 1242.760 5.940 1242.960 6.140 ;
  LAYER VI3 ;
  RECT 1242.360 6.340 1242.560 6.540 ;
  LAYER VI3 ;
  RECT 1242.360 5.940 1242.560 6.140 ;
  LAYER VI3 ;
  RECT 1241.960 6.340 1242.160 6.540 ;
  LAYER VI3 ;
  RECT 1241.960 5.940 1242.160 6.140 ;
  LAYER VI3 ;
  RECT 1241.560 6.340 1241.760 6.540 ;
  LAYER VI3 ;
  RECT 1241.560 5.940 1241.760 6.140 ;
  LAYER VI3 ;
  RECT 1241.160 6.340 1241.360 6.540 ;
  LAYER VI3 ;
  RECT 1241.160 5.940 1241.360 6.140 ;
  LAYER VI3 ;
  RECT 1240.760 6.340 1240.960 6.540 ;
  LAYER VI3 ;
  RECT 1240.760 5.940 1240.960 6.140 ;
  LAYER VI3 ;
  RECT 1240.360 6.340 1240.560 6.540 ;
  LAYER VI3 ;
  RECT 1240.360 5.940 1240.560 6.140 ;
  LAYER VI3 ;
  RECT 1239.960 6.340 1240.160 6.540 ;
  LAYER VI3 ;
  RECT 1239.960 5.940 1240.160 6.140 ;
  LAYER VI3 ;
  RECT 1239.560 6.340 1239.760 6.540 ;
  LAYER VI3 ;
  RECT 1239.560 5.940 1239.760 6.140 ;
  LAYER VI3 ;
  RECT 1239.160 6.340 1239.360 6.540 ;
  LAYER VI3 ;
  RECT 1239.160 5.940 1239.360 6.140 ;
  LAYER VI3 ;
  RECT 1238.760 6.340 1238.960 6.540 ;
  LAYER VI3 ;
  RECT 1238.760 5.940 1238.960 6.140 ;
  LAYER VI3 ;
  RECT 1238.360 6.340 1238.560 6.540 ;
  LAYER VI3 ;
  RECT 1238.360 5.940 1238.560 6.140 ;
  LAYER VI3 ;
  RECT 1237.960 6.340 1238.160 6.540 ;
  LAYER VI3 ;
  RECT 1237.960 5.940 1238.160 6.140 ;
  LAYER VI3 ;
  RECT 1237.560 6.340 1237.760 6.540 ;
  LAYER VI3 ;
  RECT 1237.560 5.940 1237.760 6.140 ;
  LAYER VI3 ;
  RECT 1237.160 6.340 1237.360 6.540 ;
  LAYER VI3 ;
  RECT 1237.160 5.940 1237.360 6.140 ;
  LAYER VI3 ;
  RECT 1236.760 6.340 1236.960 6.540 ;
  LAYER VI3 ;
  RECT 1236.760 5.940 1236.960 6.140 ;
  LAYER VI3 ;
  RECT 1236.360 6.340 1236.560 6.540 ;
  LAYER VI3 ;
  RECT 1236.360 5.940 1236.560 6.140 ;
  LAYER VI3 ;
  RECT 1235.960 6.340 1236.160 6.540 ;
  LAYER VI3 ;
  RECT 1235.960 5.940 1236.160 6.140 ;
  LAYER VI3 ;
  RECT 1255.800 5.880 1263.800 6.740 ;
  LAYER VI3 ;
  RECT 1263.400 6.340 1263.600 6.540 ;
  LAYER VI3 ;
  RECT 1263.400 5.940 1263.600 6.140 ;
  LAYER VI3 ;
  RECT 1263.000 6.340 1263.200 6.540 ;
  LAYER VI3 ;
  RECT 1263.000 5.940 1263.200 6.140 ;
  LAYER VI3 ;
  RECT 1262.600 6.340 1262.800 6.540 ;
  LAYER VI3 ;
  RECT 1262.600 5.940 1262.800 6.140 ;
  LAYER VI3 ;
  RECT 1262.200 6.340 1262.400 6.540 ;
  LAYER VI3 ;
  RECT 1262.200 5.940 1262.400 6.140 ;
  LAYER VI3 ;
  RECT 1261.800 6.340 1262.000 6.540 ;
  LAYER VI3 ;
  RECT 1261.800 5.940 1262.000 6.140 ;
  LAYER VI3 ;
  RECT 1261.400 6.340 1261.600 6.540 ;
  LAYER VI3 ;
  RECT 1261.400 5.940 1261.600 6.140 ;
  LAYER VI3 ;
  RECT 1261.000 6.340 1261.200 6.540 ;
  LAYER VI3 ;
  RECT 1261.000 5.940 1261.200 6.140 ;
  LAYER VI3 ;
  RECT 1260.600 6.340 1260.800 6.540 ;
  LAYER VI3 ;
  RECT 1260.600 5.940 1260.800 6.140 ;
  LAYER VI3 ;
  RECT 1260.200 6.340 1260.400 6.540 ;
  LAYER VI3 ;
  RECT 1260.200 5.940 1260.400 6.140 ;
  LAYER VI3 ;
  RECT 1259.800 6.340 1260.000 6.540 ;
  LAYER VI3 ;
  RECT 1259.800 5.940 1260.000 6.140 ;
  LAYER VI3 ;
  RECT 1259.400 6.340 1259.600 6.540 ;
  LAYER VI3 ;
  RECT 1259.400 5.940 1259.600 6.140 ;
  LAYER VI3 ;
  RECT 1259.000 6.340 1259.200 6.540 ;
  LAYER VI3 ;
  RECT 1259.000 5.940 1259.200 6.140 ;
  LAYER VI3 ;
  RECT 1258.600 6.340 1258.800 6.540 ;
  LAYER VI3 ;
  RECT 1258.600 5.940 1258.800 6.140 ;
  LAYER VI3 ;
  RECT 1258.200 6.340 1258.400 6.540 ;
  LAYER VI3 ;
  RECT 1258.200 5.940 1258.400 6.140 ;
  LAYER VI3 ;
  RECT 1257.800 6.340 1258.000 6.540 ;
  LAYER VI3 ;
  RECT 1257.800 5.940 1258.000 6.140 ;
  LAYER VI3 ;
  RECT 1257.400 6.340 1257.600 6.540 ;
  LAYER VI3 ;
  RECT 1257.400 5.940 1257.600 6.140 ;
  LAYER VI3 ;
  RECT 1257.000 6.340 1257.200 6.540 ;
  LAYER VI3 ;
  RECT 1257.000 5.940 1257.200 6.140 ;
  LAYER VI3 ;
  RECT 1256.600 6.340 1256.800 6.540 ;
  LAYER VI3 ;
  RECT 1256.600 5.940 1256.800 6.140 ;
  LAYER VI3 ;
  RECT 1256.200 6.340 1256.400 6.540 ;
  LAYER VI3 ;
  RECT 1256.200 5.940 1256.400 6.140 ;
  LAYER VI3 ;
  RECT 1255.800 6.340 1256.000 6.540 ;
  LAYER VI3 ;
  RECT 1255.800 5.940 1256.000 6.140 ;
  LAYER VI3 ;
  RECT 1276.880 5.880 1284.880 6.740 ;
  LAYER VI3 ;
  RECT 1284.480 6.340 1284.680 6.540 ;
  LAYER VI3 ;
  RECT 1284.480 5.940 1284.680 6.140 ;
  LAYER VI3 ;
  RECT 1284.080 6.340 1284.280 6.540 ;
  LAYER VI3 ;
  RECT 1284.080 5.940 1284.280 6.140 ;
  LAYER VI3 ;
  RECT 1283.680 6.340 1283.880 6.540 ;
  LAYER VI3 ;
  RECT 1283.680 5.940 1283.880 6.140 ;
  LAYER VI3 ;
  RECT 1283.280 6.340 1283.480 6.540 ;
  LAYER VI3 ;
  RECT 1283.280 5.940 1283.480 6.140 ;
  LAYER VI3 ;
  RECT 1282.880 6.340 1283.080 6.540 ;
  LAYER VI3 ;
  RECT 1282.880 5.940 1283.080 6.140 ;
  LAYER VI3 ;
  RECT 1282.480 6.340 1282.680 6.540 ;
  LAYER VI3 ;
  RECT 1282.480 5.940 1282.680 6.140 ;
  LAYER VI3 ;
  RECT 1282.080 6.340 1282.280 6.540 ;
  LAYER VI3 ;
  RECT 1282.080 5.940 1282.280 6.140 ;
  LAYER VI3 ;
  RECT 1281.680 6.340 1281.880 6.540 ;
  LAYER VI3 ;
  RECT 1281.680 5.940 1281.880 6.140 ;
  LAYER VI3 ;
  RECT 1281.280 6.340 1281.480 6.540 ;
  LAYER VI3 ;
  RECT 1281.280 5.940 1281.480 6.140 ;
  LAYER VI3 ;
  RECT 1280.880 6.340 1281.080 6.540 ;
  LAYER VI3 ;
  RECT 1280.880 5.940 1281.080 6.140 ;
  LAYER VI3 ;
  RECT 1280.480 6.340 1280.680 6.540 ;
  LAYER VI3 ;
  RECT 1280.480 5.940 1280.680 6.140 ;
  LAYER VI3 ;
  RECT 1280.080 6.340 1280.280 6.540 ;
  LAYER VI3 ;
  RECT 1280.080 5.940 1280.280 6.140 ;
  LAYER VI3 ;
  RECT 1279.680 6.340 1279.880 6.540 ;
  LAYER VI3 ;
  RECT 1279.680 5.940 1279.880 6.140 ;
  LAYER VI3 ;
  RECT 1279.280 6.340 1279.480 6.540 ;
  LAYER VI3 ;
  RECT 1279.280 5.940 1279.480 6.140 ;
  LAYER VI3 ;
  RECT 1278.880 6.340 1279.080 6.540 ;
  LAYER VI3 ;
  RECT 1278.880 5.940 1279.080 6.140 ;
  LAYER VI3 ;
  RECT 1278.480 6.340 1278.680 6.540 ;
  LAYER VI3 ;
  RECT 1278.480 5.940 1278.680 6.140 ;
  LAYER VI3 ;
  RECT 1278.080 6.340 1278.280 6.540 ;
  LAYER VI3 ;
  RECT 1278.080 5.940 1278.280 6.140 ;
  LAYER VI3 ;
  RECT 1277.680 6.340 1277.880 6.540 ;
  LAYER VI3 ;
  RECT 1277.680 5.940 1277.880 6.140 ;
  LAYER VI3 ;
  RECT 1277.280 6.340 1277.480 6.540 ;
  LAYER VI3 ;
  RECT 1277.280 5.940 1277.480 6.140 ;
  LAYER VI3 ;
  RECT 1276.880 6.340 1277.080 6.540 ;
  LAYER VI3 ;
  RECT 1276.880 5.940 1277.080 6.140 ;
  LAYER VI3 ;
  RECT 1296.720 5.880 1304.720 6.740 ;
  LAYER VI3 ;
  RECT 1304.320 6.340 1304.520 6.540 ;
  LAYER VI3 ;
  RECT 1304.320 5.940 1304.520 6.140 ;
  LAYER VI3 ;
  RECT 1303.920 6.340 1304.120 6.540 ;
  LAYER VI3 ;
  RECT 1303.920 5.940 1304.120 6.140 ;
  LAYER VI3 ;
  RECT 1303.520 6.340 1303.720 6.540 ;
  LAYER VI3 ;
  RECT 1303.520 5.940 1303.720 6.140 ;
  LAYER VI3 ;
  RECT 1303.120 6.340 1303.320 6.540 ;
  LAYER VI3 ;
  RECT 1303.120 5.940 1303.320 6.140 ;
  LAYER VI3 ;
  RECT 1302.720 6.340 1302.920 6.540 ;
  LAYER VI3 ;
  RECT 1302.720 5.940 1302.920 6.140 ;
  LAYER VI3 ;
  RECT 1302.320 6.340 1302.520 6.540 ;
  LAYER VI3 ;
  RECT 1302.320 5.940 1302.520 6.140 ;
  LAYER VI3 ;
  RECT 1301.920 6.340 1302.120 6.540 ;
  LAYER VI3 ;
  RECT 1301.920 5.940 1302.120 6.140 ;
  LAYER VI3 ;
  RECT 1301.520 6.340 1301.720 6.540 ;
  LAYER VI3 ;
  RECT 1301.520 5.940 1301.720 6.140 ;
  LAYER VI3 ;
  RECT 1301.120 6.340 1301.320 6.540 ;
  LAYER VI3 ;
  RECT 1301.120 5.940 1301.320 6.140 ;
  LAYER VI3 ;
  RECT 1300.720 6.340 1300.920 6.540 ;
  LAYER VI3 ;
  RECT 1300.720 5.940 1300.920 6.140 ;
  LAYER VI3 ;
  RECT 1300.320 6.340 1300.520 6.540 ;
  LAYER VI3 ;
  RECT 1300.320 5.940 1300.520 6.140 ;
  LAYER VI3 ;
  RECT 1299.920 6.340 1300.120 6.540 ;
  LAYER VI3 ;
  RECT 1299.920 5.940 1300.120 6.140 ;
  LAYER VI3 ;
  RECT 1299.520 6.340 1299.720 6.540 ;
  LAYER VI3 ;
  RECT 1299.520 5.940 1299.720 6.140 ;
  LAYER VI3 ;
  RECT 1299.120 6.340 1299.320 6.540 ;
  LAYER VI3 ;
  RECT 1299.120 5.940 1299.320 6.140 ;
  LAYER VI3 ;
  RECT 1298.720 6.340 1298.920 6.540 ;
  LAYER VI3 ;
  RECT 1298.720 5.940 1298.920 6.140 ;
  LAYER VI3 ;
  RECT 1298.320 6.340 1298.520 6.540 ;
  LAYER VI3 ;
  RECT 1298.320 5.940 1298.520 6.140 ;
  LAYER VI3 ;
  RECT 1297.920 6.340 1298.120 6.540 ;
  LAYER VI3 ;
  RECT 1297.920 5.940 1298.120 6.140 ;
  LAYER VI3 ;
  RECT 1297.520 6.340 1297.720 6.540 ;
  LAYER VI3 ;
  RECT 1297.520 5.940 1297.720 6.140 ;
  LAYER VI3 ;
  RECT 1297.120 6.340 1297.320 6.540 ;
  LAYER VI3 ;
  RECT 1297.120 5.940 1297.320 6.140 ;
  LAYER VI3 ;
  RECT 1296.720 6.340 1296.920 6.540 ;
  LAYER VI3 ;
  RECT 1296.720 5.940 1296.920 6.140 ;
  LAYER VI3 ;
  RECT 2679.800 191.940 2680.660 192.320 ;
  LAYER VI3 ;
  RECT 2680.200 192.000 2680.400 192.200 ;
  LAYER VI3 ;
  RECT 2679.800 192.000 2680.000 192.200 ;
  LAYER VI2 ;
  RECT 2679.800 191.940 2680.660 192.320 ;
  LAYER VI2 ;
  RECT 2680.200 192.000 2680.400 192.200 ;
  LAYER VI2 ;
  RECT 2679.800 192.000 2680.000 192.200 ;
  LAYER VI3 ;
  RECT 2679.800 184.020 2680.660 184.300 ;
  LAYER VI3 ;
  RECT 2680.260 184.020 2680.460 184.220 ;
  LAYER VI3 ;
  RECT 2679.860 184.020 2680.060 184.220 ;
  LAYER VI2 ;
  RECT 2679.800 184.020 2680.660 184.300 ;
  LAYER VI2 ;
  RECT 2680.260 184.020 2680.460 184.220 ;
  LAYER VI2 ;
  RECT 2679.860 184.020 2680.060 184.220 ;
  LAYER VI3 ;
  RECT 2679.800 180.340 2680.660 180.620 ;
  LAYER VI3 ;
  RECT 2680.260 180.340 2680.460 180.540 ;
  LAYER VI3 ;
  RECT 2679.860 180.340 2680.060 180.540 ;
  LAYER VI2 ;
  RECT 2679.800 180.340 2680.660 180.620 ;
  LAYER VI2 ;
  RECT 2680.260 180.340 2680.460 180.540 ;
  LAYER VI2 ;
  RECT 2679.860 180.340 2680.060 180.540 ;
  LAYER VI3 ;
  RECT 2679.800 176.660 2680.660 176.940 ;
  LAYER VI3 ;
  RECT 2680.260 176.660 2680.460 176.860 ;
  LAYER VI3 ;
  RECT 2679.860 176.660 2680.060 176.860 ;
  LAYER VI2 ;
  RECT 2679.800 176.660 2680.660 176.940 ;
  LAYER VI2 ;
  RECT 2680.260 176.660 2680.460 176.860 ;
  LAYER VI2 ;
  RECT 2679.860 176.660 2680.060 176.860 ;
  LAYER VI3 ;
  RECT 2679.800 172.980 2680.660 173.260 ;
  LAYER VI3 ;
  RECT 2680.260 172.980 2680.460 173.180 ;
  LAYER VI3 ;
  RECT 2679.860 172.980 2680.060 173.180 ;
  LAYER VI2 ;
  RECT 2679.800 172.980 2680.660 173.260 ;
  LAYER VI2 ;
  RECT 2680.260 172.980 2680.460 173.180 ;
  LAYER VI2 ;
  RECT 2679.860 172.980 2680.060 173.180 ;
  LAYER VI3 ;
  RECT 2679.800 169.300 2680.660 169.580 ;
  LAYER VI3 ;
  RECT 2680.260 169.300 2680.460 169.500 ;
  LAYER VI3 ;
  RECT 2679.860 169.300 2680.060 169.500 ;
  LAYER VI2 ;
  RECT 2679.800 169.300 2680.660 169.580 ;
  LAYER VI2 ;
  RECT 2680.260 169.300 2680.460 169.500 ;
  LAYER VI2 ;
  RECT 2679.860 169.300 2680.060 169.500 ;
  LAYER VI3 ;
  RECT 2679.800 165.620 2680.660 165.900 ;
  LAYER VI3 ;
  RECT 2680.260 165.620 2680.460 165.820 ;
  LAYER VI3 ;
  RECT 2679.860 165.620 2680.060 165.820 ;
  LAYER VI2 ;
  RECT 2679.800 165.620 2680.660 165.900 ;
  LAYER VI2 ;
  RECT 2680.260 165.620 2680.460 165.820 ;
  LAYER VI2 ;
  RECT 2679.860 165.620 2680.060 165.820 ;
  LAYER VI3 ;
  RECT 2679.800 161.940 2680.660 162.220 ;
  LAYER VI3 ;
  RECT 2680.260 161.940 2680.460 162.140 ;
  LAYER VI3 ;
  RECT 2679.860 161.940 2680.060 162.140 ;
  LAYER VI2 ;
  RECT 2679.800 161.940 2680.660 162.220 ;
  LAYER VI2 ;
  RECT 2680.260 161.940 2680.460 162.140 ;
  LAYER VI2 ;
  RECT 2679.860 161.940 2680.060 162.140 ;
  LAYER VI3 ;
  RECT 2679.800 158.260 2680.660 158.540 ;
  LAYER VI3 ;
  RECT 2680.260 158.260 2680.460 158.460 ;
  LAYER VI3 ;
  RECT 2679.860 158.260 2680.060 158.460 ;
  LAYER VI2 ;
  RECT 2679.800 158.260 2680.660 158.540 ;
  LAYER VI2 ;
  RECT 2680.260 158.260 2680.460 158.460 ;
  LAYER VI2 ;
  RECT 2679.860 158.260 2680.060 158.460 ;
  LAYER VI3 ;
  RECT 2679.800 154.580 2680.660 154.860 ;
  LAYER VI3 ;
  RECT 2680.260 154.580 2680.460 154.780 ;
  LAYER VI3 ;
  RECT 2679.860 154.580 2680.060 154.780 ;
  LAYER VI2 ;
  RECT 2679.800 154.580 2680.660 154.860 ;
  LAYER VI2 ;
  RECT 2680.260 154.580 2680.460 154.780 ;
  LAYER VI2 ;
  RECT 2679.860 154.580 2680.060 154.780 ;
  LAYER VI3 ;
  RECT 2679.800 150.900 2680.660 151.180 ;
  LAYER VI3 ;
  RECT 2680.260 150.900 2680.460 151.100 ;
  LAYER VI3 ;
  RECT 2679.860 150.900 2680.060 151.100 ;
  LAYER VI2 ;
  RECT 2679.800 150.900 2680.660 151.180 ;
  LAYER VI2 ;
  RECT 2680.260 150.900 2680.460 151.100 ;
  LAYER VI2 ;
  RECT 2679.860 150.900 2680.060 151.100 ;
  LAYER VI3 ;
  RECT 2679.800 147.220 2680.660 147.500 ;
  LAYER VI3 ;
  RECT 2680.260 147.220 2680.460 147.420 ;
  LAYER VI3 ;
  RECT 2679.860 147.220 2680.060 147.420 ;
  LAYER VI2 ;
  RECT 2679.800 147.220 2680.660 147.500 ;
  LAYER VI2 ;
  RECT 2680.260 147.220 2680.460 147.420 ;
  LAYER VI2 ;
  RECT 2679.860 147.220 2680.060 147.420 ;
  LAYER VI3 ;
  RECT 2679.800 143.540 2680.660 143.820 ;
  LAYER VI3 ;
  RECT 2680.260 143.540 2680.460 143.740 ;
  LAYER VI3 ;
  RECT 2679.860 143.540 2680.060 143.740 ;
  LAYER VI2 ;
  RECT 2679.800 143.540 2680.660 143.820 ;
  LAYER VI2 ;
  RECT 2680.260 143.540 2680.460 143.740 ;
  LAYER VI2 ;
  RECT 2679.860 143.540 2680.060 143.740 ;
  LAYER VI3 ;
  RECT 2679.800 139.860 2680.660 140.140 ;
  LAYER VI3 ;
  RECT 2680.260 139.860 2680.460 140.060 ;
  LAYER VI3 ;
  RECT 2679.860 139.860 2680.060 140.060 ;
  LAYER VI2 ;
  RECT 2679.800 139.860 2680.660 140.140 ;
  LAYER VI2 ;
  RECT 2680.260 139.860 2680.460 140.060 ;
  LAYER VI2 ;
  RECT 2679.860 139.860 2680.060 140.060 ;
  LAYER VI3 ;
  RECT 2679.800 136.180 2680.660 136.460 ;
  LAYER VI3 ;
  RECT 2680.260 136.180 2680.460 136.380 ;
  LAYER VI3 ;
  RECT 2679.860 136.180 2680.060 136.380 ;
  LAYER VI2 ;
  RECT 2679.800 136.180 2680.660 136.460 ;
  LAYER VI2 ;
  RECT 2680.260 136.180 2680.460 136.380 ;
  LAYER VI2 ;
  RECT 2679.860 136.180 2680.060 136.380 ;
  LAYER VI3 ;
  RECT 2679.800 132.500 2680.660 132.780 ;
  LAYER VI3 ;
  RECT 2680.260 132.500 2680.460 132.700 ;
  LAYER VI3 ;
  RECT 2679.860 132.500 2680.060 132.700 ;
  LAYER VI2 ;
  RECT 2679.800 132.500 2680.660 132.780 ;
  LAYER VI2 ;
  RECT 2680.260 132.500 2680.460 132.700 ;
  LAYER VI2 ;
  RECT 2679.860 132.500 2680.060 132.700 ;
  LAYER VI3 ;
  RECT 2679.800 128.820 2680.660 129.100 ;
  LAYER VI3 ;
  RECT 2680.260 128.820 2680.460 129.020 ;
  LAYER VI3 ;
  RECT 2679.860 128.820 2680.060 129.020 ;
  LAYER VI2 ;
  RECT 2679.800 128.820 2680.660 129.100 ;
  LAYER VI2 ;
  RECT 2680.260 128.820 2680.460 129.020 ;
  LAYER VI2 ;
  RECT 2679.860 128.820 2680.060 129.020 ;
  LAYER VI3 ;
  RECT 2679.800 125.140 2680.660 125.420 ;
  LAYER VI3 ;
  RECT 2680.260 125.140 2680.460 125.340 ;
  LAYER VI3 ;
  RECT 2679.860 125.140 2680.060 125.340 ;
  LAYER VI2 ;
  RECT 2679.800 125.140 2680.660 125.420 ;
  LAYER VI2 ;
  RECT 2680.260 125.140 2680.460 125.340 ;
  LAYER VI2 ;
  RECT 2679.860 125.140 2680.060 125.340 ;
  LAYER VI3 ;
  RECT 2679.800 121.460 2680.660 121.740 ;
  LAYER VI3 ;
  RECT 2680.260 121.460 2680.460 121.660 ;
  LAYER VI3 ;
  RECT 2679.860 121.460 2680.060 121.660 ;
  LAYER VI2 ;
  RECT 2679.800 121.460 2680.660 121.740 ;
  LAYER VI2 ;
  RECT 2680.260 121.460 2680.460 121.660 ;
  LAYER VI2 ;
  RECT 2679.860 121.460 2680.060 121.660 ;
  LAYER VI3 ;
  RECT 2679.800 117.780 2680.660 118.060 ;
  LAYER VI3 ;
  RECT 2680.260 117.780 2680.460 117.980 ;
  LAYER VI3 ;
  RECT 2679.860 117.780 2680.060 117.980 ;
  LAYER VI2 ;
  RECT 2679.800 117.780 2680.660 118.060 ;
  LAYER VI2 ;
  RECT 2680.260 117.780 2680.460 117.980 ;
  LAYER VI2 ;
  RECT 2679.860 117.780 2680.060 117.980 ;
  LAYER VI3 ;
  RECT 2679.800 114.100 2680.660 114.380 ;
  LAYER VI3 ;
  RECT 2680.260 114.100 2680.460 114.300 ;
  LAYER VI3 ;
  RECT 2679.860 114.100 2680.060 114.300 ;
  LAYER VI2 ;
  RECT 2679.800 114.100 2680.660 114.380 ;
  LAYER VI2 ;
  RECT 2680.260 114.100 2680.460 114.300 ;
  LAYER VI2 ;
  RECT 2679.860 114.100 2680.060 114.300 ;
  LAYER VI3 ;
  RECT 2679.800 110.420 2680.660 110.700 ;
  LAYER VI3 ;
  RECT 2680.260 110.420 2680.460 110.620 ;
  LAYER VI3 ;
  RECT 2679.860 110.420 2680.060 110.620 ;
  LAYER VI2 ;
  RECT 2679.800 110.420 2680.660 110.700 ;
  LAYER VI2 ;
  RECT 2680.260 110.420 2680.460 110.620 ;
  LAYER VI2 ;
  RECT 2679.860 110.420 2680.060 110.620 ;
  LAYER VI3 ;
  RECT 2679.800 106.740 2680.660 107.020 ;
  LAYER VI3 ;
  RECT 2680.260 106.740 2680.460 106.940 ;
  LAYER VI3 ;
  RECT 2679.860 106.740 2680.060 106.940 ;
  LAYER VI2 ;
  RECT 2679.800 106.740 2680.660 107.020 ;
  LAYER VI2 ;
  RECT 2680.260 106.740 2680.460 106.940 ;
  LAYER VI2 ;
  RECT 2679.860 106.740 2680.060 106.940 ;
  LAYER VI3 ;
  RECT 2679.800 103.060 2680.660 103.340 ;
  LAYER VI3 ;
  RECT 2680.260 103.060 2680.460 103.260 ;
  LAYER VI3 ;
  RECT 2679.860 103.060 2680.060 103.260 ;
  LAYER VI2 ;
  RECT 2679.800 103.060 2680.660 103.340 ;
  LAYER VI2 ;
  RECT 2680.260 103.060 2680.460 103.260 ;
  LAYER VI2 ;
  RECT 2679.860 103.060 2680.060 103.260 ;
  LAYER VI3 ;
  RECT 2679.800 99.380 2680.660 99.660 ;
  LAYER VI3 ;
  RECT 2680.260 99.380 2680.460 99.580 ;
  LAYER VI3 ;
  RECT 2679.860 99.380 2680.060 99.580 ;
  LAYER VI2 ;
  RECT 2679.800 99.380 2680.660 99.660 ;
  LAYER VI2 ;
  RECT 2680.260 99.380 2680.460 99.580 ;
  LAYER VI2 ;
  RECT 2679.860 99.380 2680.060 99.580 ;
  LAYER VI3 ;
  RECT 2679.800 95.700 2680.660 95.980 ;
  LAYER VI3 ;
  RECT 2680.260 95.700 2680.460 95.900 ;
  LAYER VI3 ;
  RECT 2679.860 95.700 2680.060 95.900 ;
  LAYER VI2 ;
  RECT 2679.800 95.700 2680.660 95.980 ;
  LAYER VI2 ;
  RECT 2680.260 95.700 2680.460 95.900 ;
  LAYER VI2 ;
  RECT 2679.860 95.700 2680.060 95.900 ;
  LAYER VI3 ;
  RECT 2679.800 92.020 2680.660 92.300 ;
  LAYER VI3 ;
  RECT 2680.260 92.020 2680.460 92.220 ;
  LAYER VI3 ;
  RECT 2679.860 92.020 2680.060 92.220 ;
  LAYER VI2 ;
  RECT 2679.800 92.020 2680.660 92.300 ;
  LAYER VI2 ;
  RECT 2680.260 92.020 2680.460 92.220 ;
  LAYER VI2 ;
  RECT 2679.860 92.020 2680.060 92.220 ;
  LAYER VI3 ;
  RECT 2679.800 88.340 2680.660 88.620 ;
  LAYER VI3 ;
  RECT 2680.260 88.340 2680.460 88.540 ;
  LAYER VI3 ;
  RECT 2679.860 88.340 2680.060 88.540 ;
  LAYER VI2 ;
  RECT 2679.800 88.340 2680.660 88.620 ;
  LAYER VI2 ;
  RECT 2680.260 88.340 2680.460 88.540 ;
  LAYER VI2 ;
  RECT 2679.860 88.340 2680.060 88.540 ;
  LAYER VI3 ;
  RECT 2679.800 84.660 2680.660 84.940 ;
  LAYER VI3 ;
  RECT 2680.260 84.660 2680.460 84.860 ;
  LAYER VI3 ;
  RECT 2679.860 84.660 2680.060 84.860 ;
  LAYER VI2 ;
  RECT 2679.800 84.660 2680.660 84.940 ;
  LAYER VI2 ;
  RECT 2680.260 84.660 2680.460 84.860 ;
  LAYER VI2 ;
  RECT 2679.860 84.660 2680.060 84.860 ;
  LAYER VI3 ;
  RECT 2679.800 80.980 2680.660 81.260 ;
  LAYER VI3 ;
  RECT 2680.260 80.980 2680.460 81.180 ;
  LAYER VI3 ;
  RECT 2679.860 80.980 2680.060 81.180 ;
  LAYER VI2 ;
  RECT 2679.800 80.980 2680.660 81.260 ;
  LAYER VI2 ;
  RECT 2680.260 80.980 2680.460 81.180 ;
  LAYER VI2 ;
  RECT 2679.860 80.980 2680.060 81.180 ;
  LAYER VI3 ;
  RECT 2679.800 77.300 2680.660 77.580 ;
  LAYER VI3 ;
  RECT 2680.260 77.300 2680.460 77.500 ;
  LAYER VI3 ;
  RECT 2679.860 77.300 2680.060 77.500 ;
  LAYER VI2 ;
  RECT 2679.800 77.300 2680.660 77.580 ;
  LAYER VI2 ;
  RECT 2680.260 77.300 2680.460 77.500 ;
  LAYER VI2 ;
  RECT 2679.860 77.300 2680.060 77.500 ;
  LAYER VI3 ;
  RECT 2679.800 73.620 2680.660 73.900 ;
  LAYER VI3 ;
  RECT 2680.260 73.620 2680.460 73.820 ;
  LAYER VI3 ;
  RECT 2679.860 73.620 2680.060 73.820 ;
  LAYER VI2 ;
  RECT 2679.800 73.620 2680.660 73.900 ;
  LAYER VI2 ;
  RECT 2680.260 73.620 2680.460 73.820 ;
  LAYER VI2 ;
  RECT 2679.860 73.620 2680.060 73.820 ;
  LAYER VI3 ;
  RECT 2679.800 69.940 2680.660 70.220 ;
  LAYER VI3 ;
  RECT 2680.260 69.940 2680.460 70.140 ;
  LAYER VI3 ;
  RECT 2679.860 69.940 2680.060 70.140 ;
  LAYER VI2 ;
  RECT 2679.800 69.940 2680.660 70.220 ;
  LAYER VI2 ;
  RECT 2680.260 69.940 2680.460 70.140 ;
  LAYER VI2 ;
  RECT 2679.860 69.940 2680.060 70.140 ;
  LAYER VI3 ;
  RECT 2679.800 65.600 2680.660 65.980 ;
  LAYER VI3 ;
  RECT 2680.200 65.660 2680.400 65.860 ;
  LAYER VI3 ;
  RECT 2679.800 65.660 2680.000 65.860 ;
  LAYER VI2 ;
  RECT 2679.800 65.600 2680.660 65.980 ;
  LAYER VI2 ;
  RECT 2680.200 65.660 2680.400 65.860 ;
  LAYER VI2 ;
  RECT 2679.800 65.660 2680.000 65.860 ;
  LAYER VI3 ;
  RECT 1368.820 192.790 1369.070 193.650 ;
  LAYER VI3 ;
  RECT 1368.820 193.250 1369.020 193.450 ;
  LAYER VI3 ;
  RECT 1368.820 192.850 1369.020 193.050 ;
  LAYER VI2 ;
  RECT 1368.820 192.790 1369.070 193.650 ;
  LAYER VI2 ;
  RECT 1368.820 193.250 1369.020 193.450 ;
  LAYER VI2 ;
  RECT 1368.820 192.850 1369.020 193.050 ;
  LAYER VI3 ;
  RECT 1409.740 192.790 1409.990 193.650 ;
  LAYER VI3 ;
  RECT 1409.740 193.250 1409.940 193.450 ;
  LAYER VI3 ;
  RECT 1409.740 192.850 1409.940 193.050 ;
  LAYER VI2 ;
  RECT 1409.740 192.790 1409.990 193.650 ;
  LAYER VI2 ;
  RECT 1409.740 193.250 1409.940 193.450 ;
  LAYER VI2 ;
  RECT 1409.740 192.850 1409.940 193.050 ;
  LAYER VI3 ;
  RECT 1450.660 192.790 1450.910 193.650 ;
  LAYER VI3 ;
  RECT 1450.660 193.250 1450.860 193.450 ;
  LAYER VI3 ;
  RECT 1450.660 192.850 1450.860 193.050 ;
  LAYER VI2 ;
  RECT 1450.660 192.790 1450.910 193.650 ;
  LAYER VI2 ;
  RECT 1450.660 193.250 1450.860 193.450 ;
  LAYER VI2 ;
  RECT 1450.660 192.850 1450.860 193.050 ;
  LAYER VI3 ;
  RECT 1491.580 192.790 1491.830 193.650 ;
  LAYER VI3 ;
  RECT 1491.580 193.250 1491.780 193.450 ;
  LAYER VI3 ;
  RECT 1491.580 192.850 1491.780 193.050 ;
  LAYER VI2 ;
  RECT 1491.580 192.790 1491.830 193.650 ;
  LAYER VI2 ;
  RECT 1491.580 193.250 1491.780 193.450 ;
  LAYER VI2 ;
  RECT 1491.580 192.850 1491.780 193.050 ;
  LAYER VI3 ;
  RECT 1532.500 192.790 1532.750 193.650 ;
  LAYER VI3 ;
  RECT 1532.500 193.250 1532.700 193.450 ;
  LAYER VI3 ;
  RECT 1532.500 192.850 1532.700 193.050 ;
  LAYER VI2 ;
  RECT 1532.500 192.790 1532.750 193.650 ;
  LAYER VI2 ;
  RECT 1532.500 193.250 1532.700 193.450 ;
  LAYER VI2 ;
  RECT 1532.500 192.850 1532.700 193.050 ;
  LAYER VI3 ;
  RECT 1573.420 192.790 1573.670 193.650 ;
  LAYER VI3 ;
  RECT 1573.420 193.250 1573.620 193.450 ;
  LAYER VI3 ;
  RECT 1573.420 192.850 1573.620 193.050 ;
  LAYER VI2 ;
  RECT 1573.420 192.790 1573.670 193.650 ;
  LAYER VI2 ;
  RECT 1573.420 193.250 1573.620 193.450 ;
  LAYER VI2 ;
  RECT 1573.420 192.850 1573.620 193.050 ;
  LAYER VI3 ;
  RECT 1614.340 192.790 1614.590 193.650 ;
  LAYER VI3 ;
  RECT 1614.340 193.250 1614.540 193.450 ;
  LAYER VI3 ;
  RECT 1614.340 192.850 1614.540 193.050 ;
  LAYER VI2 ;
  RECT 1614.340 192.790 1614.590 193.650 ;
  LAYER VI2 ;
  RECT 1614.340 193.250 1614.540 193.450 ;
  LAYER VI2 ;
  RECT 1614.340 192.850 1614.540 193.050 ;
  LAYER VI3 ;
  RECT 1655.260 192.790 1655.510 193.650 ;
  LAYER VI3 ;
  RECT 1655.260 193.250 1655.460 193.450 ;
  LAYER VI3 ;
  RECT 1655.260 192.850 1655.460 193.050 ;
  LAYER VI2 ;
  RECT 1655.260 192.790 1655.510 193.650 ;
  LAYER VI2 ;
  RECT 1655.260 193.250 1655.460 193.450 ;
  LAYER VI2 ;
  RECT 1655.260 192.850 1655.460 193.050 ;
  LAYER VI3 ;
  RECT 1696.180 192.790 1696.430 193.650 ;
  LAYER VI3 ;
  RECT 1696.180 193.250 1696.380 193.450 ;
  LAYER VI3 ;
  RECT 1696.180 192.850 1696.380 193.050 ;
  LAYER VI2 ;
  RECT 1696.180 192.790 1696.430 193.650 ;
  LAYER VI2 ;
  RECT 1696.180 193.250 1696.380 193.450 ;
  LAYER VI2 ;
  RECT 1696.180 192.850 1696.380 193.050 ;
  LAYER VI3 ;
  RECT 1737.100 192.790 1737.350 193.650 ;
  LAYER VI3 ;
  RECT 1737.100 193.250 1737.300 193.450 ;
  LAYER VI3 ;
  RECT 1737.100 192.850 1737.300 193.050 ;
  LAYER VI2 ;
  RECT 1737.100 192.790 1737.350 193.650 ;
  LAYER VI2 ;
  RECT 1737.100 193.250 1737.300 193.450 ;
  LAYER VI2 ;
  RECT 1737.100 192.850 1737.300 193.050 ;
  LAYER VI3 ;
  RECT 1778.020 192.790 1778.270 193.650 ;
  LAYER VI3 ;
  RECT 1778.020 193.250 1778.220 193.450 ;
  LAYER VI3 ;
  RECT 1778.020 192.850 1778.220 193.050 ;
  LAYER VI2 ;
  RECT 1778.020 192.790 1778.270 193.650 ;
  LAYER VI2 ;
  RECT 1778.020 193.250 1778.220 193.450 ;
  LAYER VI2 ;
  RECT 1778.020 192.850 1778.220 193.050 ;
  LAYER VI3 ;
  RECT 1818.940 192.790 1819.190 193.650 ;
  LAYER VI3 ;
  RECT 1818.940 193.250 1819.140 193.450 ;
  LAYER VI3 ;
  RECT 1818.940 192.850 1819.140 193.050 ;
  LAYER VI2 ;
  RECT 1818.940 192.790 1819.190 193.650 ;
  LAYER VI2 ;
  RECT 1818.940 193.250 1819.140 193.450 ;
  LAYER VI2 ;
  RECT 1818.940 192.850 1819.140 193.050 ;
  LAYER VI3 ;
  RECT 1859.860 192.790 1860.110 193.650 ;
  LAYER VI3 ;
  RECT 1859.860 193.250 1860.060 193.450 ;
  LAYER VI3 ;
  RECT 1859.860 192.850 1860.060 193.050 ;
  LAYER VI2 ;
  RECT 1859.860 192.790 1860.110 193.650 ;
  LAYER VI2 ;
  RECT 1859.860 193.250 1860.060 193.450 ;
  LAYER VI2 ;
  RECT 1859.860 192.850 1860.060 193.050 ;
  LAYER VI3 ;
  RECT 1900.780 192.790 1901.030 193.650 ;
  LAYER VI3 ;
  RECT 1900.780 193.250 1900.980 193.450 ;
  LAYER VI3 ;
  RECT 1900.780 192.850 1900.980 193.050 ;
  LAYER VI2 ;
  RECT 1900.780 192.790 1901.030 193.650 ;
  LAYER VI2 ;
  RECT 1900.780 193.250 1900.980 193.450 ;
  LAYER VI2 ;
  RECT 1900.780 192.850 1900.980 193.050 ;
  LAYER VI3 ;
  RECT 1941.700 192.790 1941.950 193.650 ;
  LAYER VI3 ;
  RECT 1941.700 193.250 1941.900 193.450 ;
  LAYER VI3 ;
  RECT 1941.700 192.850 1941.900 193.050 ;
  LAYER VI2 ;
  RECT 1941.700 192.790 1941.950 193.650 ;
  LAYER VI2 ;
  RECT 1941.700 193.250 1941.900 193.450 ;
  LAYER VI2 ;
  RECT 1941.700 192.850 1941.900 193.050 ;
  LAYER VI3 ;
  RECT 1982.620 192.790 1982.870 193.650 ;
  LAYER VI3 ;
  RECT 1982.620 193.250 1982.820 193.450 ;
  LAYER VI3 ;
  RECT 1982.620 192.850 1982.820 193.050 ;
  LAYER VI2 ;
  RECT 1982.620 192.790 1982.870 193.650 ;
  LAYER VI2 ;
  RECT 1982.620 193.250 1982.820 193.450 ;
  LAYER VI2 ;
  RECT 1982.620 192.850 1982.820 193.050 ;
  LAYER VI3 ;
  RECT 2023.540 192.790 2023.790 193.650 ;
  LAYER VI3 ;
  RECT 2023.540 193.250 2023.740 193.450 ;
  LAYER VI3 ;
  RECT 2023.540 192.850 2023.740 193.050 ;
  LAYER VI2 ;
  RECT 2023.540 192.790 2023.790 193.650 ;
  LAYER VI2 ;
  RECT 2023.540 193.250 2023.740 193.450 ;
  LAYER VI2 ;
  RECT 2023.540 192.850 2023.740 193.050 ;
  LAYER VI3 ;
  RECT 2064.460 192.790 2064.710 193.650 ;
  LAYER VI3 ;
  RECT 2064.460 193.250 2064.660 193.450 ;
  LAYER VI3 ;
  RECT 2064.460 192.850 2064.660 193.050 ;
  LAYER VI2 ;
  RECT 2064.460 192.790 2064.710 193.650 ;
  LAYER VI2 ;
  RECT 2064.460 193.250 2064.660 193.450 ;
  LAYER VI2 ;
  RECT 2064.460 192.850 2064.660 193.050 ;
  LAYER VI3 ;
  RECT 2105.380 192.790 2105.630 193.650 ;
  LAYER VI3 ;
  RECT 2105.380 193.250 2105.580 193.450 ;
  LAYER VI3 ;
  RECT 2105.380 192.850 2105.580 193.050 ;
  LAYER VI2 ;
  RECT 2105.380 192.790 2105.630 193.650 ;
  LAYER VI2 ;
  RECT 2105.380 193.250 2105.580 193.450 ;
  LAYER VI2 ;
  RECT 2105.380 192.850 2105.580 193.050 ;
  LAYER VI3 ;
  RECT 2146.300 192.790 2146.550 193.650 ;
  LAYER VI3 ;
  RECT 2146.300 193.250 2146.500 193.450 ;
  LAYER VI3 ;
  RECT 2146.300 192.850 2146.500 193.050 ;
  LAYER VI2 ;
  RECT 2146.300 192.790 2146.550 193.650 ;
  LAYER VI2 ;
  RECT 2146.300 193.250 2146.500 193.450 ;
  LAYER VI2 ;
  RECT 2146.300 192.850 2146.500 193.050 ;
  LAYER VI3 ;
  RECT 2187.220 192.790 2187.470 193.650 ;
  LAYER VI3 ;
  RECT 2187.220 193.250 2187.420 193.450 ;
  LAYER VI3 ;
  RECT 2187.220 192.850 2187.420 193.050 ;
  LAYER VI2 ;
  RECT 2187.220 192.790 2187.470 193.650 ;
  LAYER VI2 ;
  RECT 2187.220 193.250 2187.420 193.450 ;
  LAYER VI2 ;
  RECT 2187.220 192.850 2187.420 193.050 ;
  LAYER VI3 ;
  RECT 2228.140 192.790 2228.390 193.650 ;
  LAYER VI3 ;
  RECT 2228.140 193.250 2228.340 193.450 ;
  LAYER VI3 ;
  RECT 2228.140 192.850 2228.340 193.050 ;
  LAYER VI2 ;
  RECT 2228.140 192.790 2228.390 193.650 ;
  LAYER VI2 ;
  RECT 2228.140 193.250 2228.340 193.450 ;
  LAYER VI2 ;
  RECT 2228.140 192.850 2228.340 193.050 ;
  LAYER VI3 ;
  RECT 2269.060 192.790 2269.310 193.650 ;
  LAYER VI3 ;
  RECT 2269.060 193.250 2269.260 193.450 ;
  LAYER VI3 ;
  RECT 2269.060 192.850 2269.260 193.050 ;
  LAYER VI2 ;
  RECT 2269.060 192.790 2269.310 193.650 ;
  LAYER VI2 ;
  RECT 2269.060 193.250 2269.260 193.450 ;
  LAYER VI2 ;
  RECT 2269.060 192.850 2269.260 193.050 ;
  LAYER VI3 ;
  RECT 2309.980 192.790 2310.230 193.650 ;
  LAYER VI3 ;
  RECT 2309.980 193.250 2310.180 193.450 ;
  LAYER VI3 ;
  RECT 2309.980 192.850 2310.180 193.050 ;
  LAYER VI2 ;
  RECT 2309.980 192.790 2310.230 193.650 ;
  LAYER VI2 ;
  RECT 2309.980 193.250 2310.180 193.450 ;
  LAYER VI2 ;
  RECT 2309.980 192.850 2310.180 193.050 ;
  LAYER VI3 ;
  RECT 2350.900 192.790 2351.150 193.650 ;
  LAYER VI3 ;
  RECT 2350.900 193.250 2351.100 193.450 ;
  LAYER VI3 ;
  RECT 2350.900 192.850 2351.100 193.050 ;
  LAYER VI2 ;
  RECT 2350.900 192.790 2351.150 193.650 ;
  LAYER VI2 ;
  RECT 2350.900 193.250 2351.100 193.450 ;
  LAYER VI2 ;
  RECT 2350.900 192.850 2351.100 193.050 ;
  LAYER VI3 ;
  RECT 2391.820 192.790 2392.070 193.650 ;
  LAYER VI3 ;
  RECT 2391.820 193.250 2392.020 193.450 ;
  LAYER VI3 ;
  RECT 2391.820 192.850 2392.020 193.050 ;
  LAYER VI2 ;
  RECT 2391.820 192.790 2392.070 193.650 ;
  LAYER VI2 ;
  RECT 2391.820 193.250 2392.020 193.450 ;
  LAYER VI2 ;
  RECT 2391.820 192.850 2392.020 193.050 ;
  LAYER VI3 ;
  RECT 2432.740 192.790 2432.990 193.650 ;
  LAYER VI3 ;
  RECT 2432.740 193.250 2432.940 193.450 ;
  LAYER VI3 ;
  RECT 2432.740 192.850 2432.940 193.050 ;
  LAYER VI2 ;
  RECT 2432.740 192.790 2432.990 193.650 ;
  LAYER VI2 ;
  RECT 2432.740 193.250 2432.940 193.450 ;
  LAYER VI2 ;
  RECT 2432.740 192.850 2432.940 193.050 ;
  LAYER VI3 ;
  RECT 2473.660 192.790 2473.910 193.650 ;
  LAYER VI3 ;
  RECT 2473.660 193.250 2473.860 193.450 ;
  LAYER VI3 ;
  RECT 2473.660 192.850 2473.860 193.050 ;
  LAYER VI2 ;
  RECT 2473.660 192.790 2473.910 193.650 ;
  LAYER VI2 ;
  RECT 2473.660 193.250 2473.860 193.450 ;
  LAYER VI2 ;
  RECT 2473.660 192.850 2473.860 193.050 ;
  LAYER VI3 ;
  RECT 2514.580 192.790 2514.830 193.650 ;
  LAYER VI3 ;
  RECT 2514.580 193.250 2514.780 193.450 ;
  LAYER VI3 ;
  RECT 2514.580 192.850 2514.780 193.050 ;
  LAYER VI2 ;
  RECT 2514.580 192.790 2514.830 193.650 ;
  LAYER VI2 ;
  RECT 2514.580 193.250 2514.780 193.450 ;
  LAYER VI2 ;
  RECT 2514.580 192.850 2514.780 193.050 ;
  LAYER VI3 ;
  RECT 2555.500 192.790 2555.750 193.650 ;
  LAYER VI3 ;
  RECT 2555.500 193.250 2555.700 193.450 ;
  LAYER VI3 ;
  RECT 2555.500 192.850 2555.700 193.050 ;
  LAYER VI2 ;
  RECT 2555.500 192.790 2555.750 193.650 ;
  LAYER VI2 ;
  RECT 2555.500 193.250 2555.700 193.450 ;
  LAYER VI2 ;
  RECT 2555.500 192.850 2555.700 193.050 ;
  LAYER VI3 ;
  RECT 2596.420 192.790 2596.670 193.650 ;
  LAYER VI3 ;
  RECT 2596.420 193.250 2596.620 193.450 ;
  LAYER VI3 ;
  RECT 2596.420 192.850 2596.620 193.050 ;
  LAYER VI2 ;
  RECT 2596.420 192.790 2596.670 193.650 ;
  LAYER VI2 ;
  RECT 2596.420 193.250 2596.620 193.450 ;
  LAYER VI2 ;
  RECT 2596.420 192.850 2596.620 193.050 ;
  LAYER VI3 ;
  RECT 2637.340 192.790 2637.590 193.650 ;
  LAYER VI3 ;
  RECT 2637.340 193.250 2637.540 193.450 ;
  LAYER VI3 ;
  RECT 2637.340 192.850 2637.540 193.050 ;
  LAYER VI2 ;
  RECT 2637.340 192.790 2637.590 193.650 ;
  LAYER VI2 ;
  RECT 2637.340 193.250 2637.540 193.450 ;
  LAYER VI2 ;
  RECT 2637.340 192.850 2637.540 193.050 ;
  LAYER VI3 ;
  RECT 1351.810 192.790 1354.320 193.650 ;
  LAYER VI3 ;
  RECT 1353.810 193.250 1354.010 193.450 ;
  LAYER VI3 ;
  RECT 1353.810 192.850 1354.010 193.050 ;
  LAYER VI3 ;
  RECT 1353.410 193.250 1353.610 193.450 ;
  LAYER VI3 ;
  RECT 1353.410 192.850 1353.610 193.050 ;
  LAYER VI3 ;
  RECT 1353.010 193.250 1353.210 193.450 ;
  LAYER VI3 ;
  RECT 1353.010 192.850 1353.210 193.050 ;
  LAYER VI3 ;
  RECT 1352.610 193.250 1352.810 193.450 ;
  LAYER VI3 ;
  RECT 1352.610 192.850 1352.810 193.050 ;
  LAYER VI3 ;
  RECT 1352.210 193.250 1352.410 193.450 ;
  LAYER VI3 ;
  RECT 1352.210 192.850 1352.410 193.050 ;
  LAYER VI3 ;
  RECT 1351.810 193.250 1352.010 193.450 ;
  LAYER VI3 ;
  RECT 1351.810 192.850 1352.010 193.050 ;
  LAYER VI2 ;
  RECT 1351.810 192.790 1354.320 193.650 ;
  LAYER VI2 ;
  RECT 1353.810 193.250 1354.010 193.450 ;
  LAYER VI2 ;
  RECT 1353.810 192.850 1354.010 193.050 ;
  LAYER VI2 ;
  RECT 1353.410 193.250 1353.610 193.450 ;
  LAYER VI2 ;
  RECT 1353.410 192.850 1353.610 193.050 ;
  LAYER VI2 ;
  RECT 1353.010 193.250 1353.210 193.450 ;
  LAYER VI2 ;
  RECT 1353.010 192.850 1353.210 193.050 ;
  LAYER VI2 ;
  RECT 1352.610 193.250 1352.810 193.450 ;
  LAYER VI2 ;
  RECT 1352.610 192.850 1352.810 193.050 ;
  LAYER VI2 ;
  RECT 1352.210 193.250 1352.410 193.450 ;
  LAYER VI2 ;
  RECT 1352.210 192.850 1352.410 193.050 ;
  LAYER VI2 ;
  RECT 1351.810 193.250 1352.010 193.450 ;
  LAYER VI2 ;
  RECT 1351.810 192.850 1352.010 193.050 ;
  LAYER VI3 ;
  RECT 1339.390 192.790 1341.780 193.650 ;
  LAYER VI3 ;
  RECT 1341.390 193.250 1341.590 193.450 ;
  LAYER VI3 ;
  RECT 1341.390 192.850 1341.590 193.050 ;
  LAYER VI3 ;
  RECT 1340.990 193.250 1341.190 193.450 ;
  LAYER VI3 ;
  RECT 1340.990 192.850 1341.190 193.050 ;
  LAYER VI3 ;
  RECT 1340.590 193.250 1340.790 193.450 ;
  LAYER VI3 ;
  RECT 1340.590 192.850 1340.790 193.050 ;
  LAYER VI3 ;
  RECT 1340.190 193.250 1340.390 193.450 ;
  LAYER VI3 ;
  RECT 1340.190 192.850 1340.390 193.050 ;
  LAYER VI3 ;
  RECT 1339.790 193.250 1339.990 193.450 ;
  LAYER VI3 ;
  RECT 1339.790 192.850 1339.990 193.050 ;
  LAYER VI3 ;
  RECT 1339.390 193.250 1339.590 193.450 ;
  LAYER VI3 ;
  RECT 1339.390 192.850 1339.590 193.050 ;
  LAYER VI2 ;
  RECT 1339.390 192.790 1341.780 193.650 ;
  LAYER VI2 ;
  RECT 1341.390 193.250 1341.590 193.450 ;
  LAYER VI2 ;
  RECT 1341.390 192.850 1341.590 193.050 ;
  LAYER VI2 ;
  RECT 1340.990 193.250 1341.190 193.450 ;
  LAYER VI2 ;
  RECT 1340.990 192.850 1341.190 193.050 ;
  LAYER VI2 ;
  RECT 1340.590 193.250 1340.790 193.450 ;
  LAYER VI2 ;
  RECT 1340.590 192.850 1340.790 193.050 ;
  LAYER VI2 ;
  RECT 1340.190 193.250 1340.390 193.450 ;
  LAYER VI2 ;
  RECT 1340.190 192.850 1340.390 193.050 ;
  LAYER VI2 ;
  RECT 1339.790 193.250 1339.990 193.450 ;
  LAYER VI2 ;
  RECT 1339.790 192.850 1339.990 193.050 ;
  LAYER VI2 ;
  RECT 1339.390 193.250 1339.590 193.450 ;
  LAYER VI2 ;
  RECT 1339.390 192.850 1339.590 193.050 ;
  LAYER VI3 ;
  RECT 1331.880 192.790 1334.940 193.650 ;
  LAYER VI3 ;
  RECT 1334.680 193.250 1334.880 193.450 ;
  LAYER VI3 ;
  RECT 1334.680 192.850 1334.880 193.050 ;
  LAYER VI3 ;
  RECT 1334.280 193.250 1334.480 193.450 ;
  LAYER VI3 ;
  RECT 1334.280 192.850 1334.480 193.050 ;
  LAYER VI3 ;
  RECT 1333.880 193.250 1334.080 193.450 ;
  LAYER VI3 ;
  RECT 1333.880 192.850 1334.080 193.050 ;
  LAYER VI3 ;
  RECT 1333.480 193.250 1333.680 193.450 ;
  LAYER VI3 ;
  RECT 1333.480 192.850 1333.680 193.050 ;
  LAYER VI3 ;
  RECT 1333.080 193.250 1333.280 193.450 ;
  LAYER VI3 ;
  RECT 1333.080 192.850 1333.280 193.050 ;
  LAYER VI3 ;
  RECT 1332.680 193.250 1332.880 193.450 ;
  LAYER VI3 ;
  RECT 1332.680 192.850 1332.880 193.050 ;
  LAYER VI3 ;
  RECT 1332.280 193.250 1332.480 193.450 ;
  LAYER VI3 ;
  RECT 1332.280 192.850 1332.480 193.050 ;
  LAYER VI3 ;
  RECT 1331.880 193.250 1332.080 193.450 ;
  LAYER VI3 ;
  RECT 1331.880 192.850 1332.080 193.050 ;
  LAYER VI2 ;
  RECT 1331.880 192.790 1334.940 193.650 ;
  LAYER VI2 ;
  RECT 1334.680 193.250 1334.880 193.450 ;
  LAYER VI2 ;
  RECT 1334.680 192.850 1334.880 193.050 ;
  LAYER VI2 ;
  RECT 1334.280 193.250 1334.480 193.450 ;
  LAYER VI2 ;
  RECT 1334.280 192.850 1334.480 193.050 ;
  LAYER VI2 ;
  RECT 1333.880 193.250 1334.080 193.450 ;
  LAYER VI2 ;
  RECT 1333.880 192.850 1334.080 193.050 ;
  LAYER VI2 ;
  RECT 1333.480 193.250 1333.680 193.450 ;
  LAYER VI2 ;
  RECT 1333.480 192.850 1333.680 193.050 ;
  LAYER VI2 ;
  RECT 1333.080 193.250 1333.280 193.450 ;
  LAYER VI2 ;
  RECT 1333.080 192.850 1333.280 193.050 ;
  LAYER VI2 ;
  RECT 1332.680 193.250 1332.880 193.450 ;
  LAYER VI2 ;
  RECT 1332.680 192.850 1332.880 193.050 ;
  LAYER VI2 ;
  RECT 1332.280 193.250 1332.480 193.450 ;
  LAYER VI2 ;
  RECT 1332.280 192.850 1332.480 193.050 ;
  LAYER VI2 ;
  RECT 1331.880 193.250 1332.080 193.450 ;
  LAYER VI2 ;
  RECT 1331.880 192.850 1332.080 193.050 ;
  LAYER VI3 ;
  RECT 1356.060 192.790 1358.910 193.650 ;
  LAYER VI3 ;
  RECT 1358.460 193.250 1358.660 193.450 ;
  LAYER VI3 ;
  RECT 1358.460 192.850 1358.660 193.050 ;
  LAYER VI3 ;
  RECT 1358.060 193.250 1358.260 193.450 ;
  LAYER VI3 ;
  RECT 1358.060 192.850 1358.260 193.050 ;
  LAYER VI3 ;
  RECT 1357.660 193.250 1357.860 193.450 ;
  LAYER VI3 ;
  RECT 1357.660 192.850 1357.860 193.050 ;
  LAYER VI3 ;
  RECT 1357.260 193.250 1357.460 193.450 ;
  LAYER VI3 ;
  RECT 1357.260 192.850 1357.460 193.050 ;
  LAYER VI3 ;
  RECT 1356.860 193.250 1357.060 193.450 ;
  LAYER VI3 ;
  RECT 1356.860 192.850 1357.060 193.050 ;
  LAYER VI3 ;
  RECT 1356.460 193.250 1356.660 193.450 ;
  LAYER VI3 ;
  RECT 1356.460 192.850 1356.660 193.050 ;
  LAYER VI3 ;
  RECT 1356.060 193.250 1356.260 193.450 ;
  LAYER VI3 ;
  RECT 1356.060 192.850 1356.260 193.050 ;
  LAYER VI2 ;
  RECT 1356.060 192.790 1358.910 193.650 ;
  LAYER VI2 ;
  RECT 1358.460 193.250 1358.660 193.450 ;
  LAYER VI2 ;
  RECT 1358.460 192.850 1358.660 193.050 ;
  LAYER VI2 ;
  RECT 1358.060 193.250 1358.260 193.450 ;
  LAYER VI2 ;
  RECT 1358.060 192.850 1358.260 193.050 ;
  LAYER VI2 ;
  RECT 1357.660 193.250 1357.860 193.450 ;
  LAYER VI2 ;
  RECT 1357.660 192.850 1357.860 193.050 ;
  LAYER VI2 ;
  RECT 1357.260 193.250 1357.460 193.450 ;
  LAYER VI2 ;
  RECT 1357.260 192.850 1357.460 193.050 ;
  LAYER VI2 ;
  RECT 1356.860 193.250 1357.060 193.450 ;
  LAYER VI2 ;
  RECT 1356.860 192.850 1357.060 193.050 ;
  LAYER VI2 ;
  RECT 1356.460 193.250 1356.660 193.450 ;
  LAYER VI2 ;
  RECT 1356.460 192.850 1356.660 193.050 ;
  LAYER VI2 ;
  RECT 1356.060 193.250 1356.260 193.450 ;
  LAYER VI2 ;
  RECT 1356.060 192.850 1356.260 193.050 ;
  LAYER VI3 ;
  RECT 1360.360 192.790 1363.610 193.650 ;
  LAYER VI3 ;
  RECT 1363.160 193.250 1363.360 193.450 ;
  LAYER VI3 ;
  RECT 1363.160 192.850 1363.360 193.050 ;
  LAYER VI3 ;
  RECT 1362.760 193.250 1362.960 193.450 ;
  LAYER VI3 ;
  RECT 1362.760 192.850 1362.960 193.050 ;
  LAYER VI3 ;
  RECT 1362.360 193.250 1362.560 193.450 ;
  LAYER VI3 ;
  RECT 1362.360 192.850 1362.560 193.050 ;
  LAYER VI3 ;
  RECT 1361.960 193.250 1362.160 193.450 ;
  LAYER VI3 ;
  RECT 1361.960 192.850 1362.160 193.050 ;
  LAYER VI3 ;
  RECT 1361.560 193.250 1361.760 193.450 ;
  LAYER VI3 ;
  RECT 1361.560 192.850 1361.760 193.050 ;
  LAYER VI3 ;
  RECT 1361.160 193.250 1361.360 193.450 ;
  LAYER VI3 ;
  RECT 1361.160 192.850 1361.360 193.050 ;
  LAYER VI3 ;
  RECT 1360.760 193.250 1360.960 193.450 ;
  LAYER VI3 ;
  RECT 1360.760 192.850 1360.960 193.050 ;
  LAYER VI3 ;
  RECT 1360.360 193.250 1360.560 193.450 ;
  LAYER VI3 ;
  RECT 1360.360 192.850 1360.560 193.050 ;
  LAYER VI2 ;
  RECT 1360.360 192.790 1363.610 193.650 ;
  LAYER VI2 ;
  RECT 1363.160 193.250 1363.360 193.450 ;
  LAYER VI2 ;
  RECT 1363.160 192.850 1363.360 193.050 ;
  LAYER VI2 ;
  RECT 1362.760 193.250 1362.960 193.450 ;
  LAYER VI2 ;
  RECT 1362.760 192.850 1362.960 193.050 ;
  LAYER VI2 ;
  RECT 1362.360 193.250 1362.560 193.450 ;
  LAYER VI2 ;
  RECT 1362.360 192.850 1362.560 193.050 ;
  LAYER VI2 ;
  RECT 1361.960 193.250 1362.160 193.450 ;
  LAYER VI2 ;
  RECT 1361.960 192.850 1362.160 193.050 ;
  LAYER VI2 ;
  RECT 1361.560 193.250 1361.760 193.450 ;
  LAYER VI2 ;
  RECT 1361.560 192.850 1361.760 193.050 ;
  LAYER VI2 ;
  RECT 1361.160 193.250 1361.360 193.450 ;
  LAYER VI2 ;
  RECT 1361.160 192.850 1361.360 193.050 ;
  LAYER VI2 ;
  RECT 1360.760 193.250 1360.960 193.450 ;
  LAYER VI2 ;
  RECT 1360.760 192.850 1360.960 193.050 ;
  LAYER VI2 ;
  RECT 1360.360 193.250 1360.560 193.450 ;
  LAYER VI2 ;
  RECT 1360.360 192.850 1360.560 193.050 ;
  LAYER VI3 ;
  RECT 1329.160 192.790 1330.920 193.650 ;
  LAYER VI3 ;
  RECT 1330.360 193.250 1330.560 193.450 ;
  LAYER VI3 ;
  RECT 1330.360 192.850 1330.560 193.050 ;
  LAYER VI3 ;
  RECT 1329.960 193.250 1330.160 193.450 ;
  LAYER VI3 ;
  RECT 1329.960 192.850 1330.160 193.050 ;
  LAYER VI3 ;
  RECT 1329.560 193.250 1329.760 193.450 ;
  LAYER VI3 ;
  RECT 1329.560 192.850 1329.760 193.050 ;
  LAYER VI3 ;
  RECT 1329.160 193.250 1329.360 193.450 ;
  LAYER VI3 ;
  RECT 1329.160 192.850 1329.360 193.050 ;
  LAYER VI2 ;
  RECT 1329.160 192.790 1330.920 193.650 ;
  LAYER VI2 ;
  RECT 1330.360 193.250 1330.560 193.450 ;
  LAYER VI2 ;
  RECT 1330.360 192.850 1330.560 193.050 ;
  LAYER VI2 ;
  RECT 1329.960 193.250 1330.160 193.450 ;
  LAYER VI2 ;
  RECT 1329.960 192.850 1330.160 193.050 ;
  LAYER VI2 ;
  RECT 1329.560 193.250 1329.760 193.450 ;
  LAYER VI2 ;
  RECT 1329.560 192.850 1329.760 193.050 ;
  LAYER VI2 ;
  RECT 1329.160 193.250 1329.360 193.450 ;
  LAYER VI2 ;
  RECT 1329.160 192.850 1329.360 193.050 ;
  LAYER VI3 ;
  RECT 1319.820 192.790 1321.580 193.650 ;
  LAYER VI3 ;
  RECT 1321.020 193.250 1321.220 193.450 ;
  LAYER VI3 ;
  RECT 1321.020 192.850 1321.220 193.050 ;
  LAYER VI3 ;
  RECT 1320.620 193.250 1320.820 193.450 ;
  LAYER VI3 ;
  RECT 1320.620 192.850 1320.820 193.050 ;
  LAYER VI3 ;
  RECT 1320.220 193.250 1320.420 193.450 ;
  LAYER VI3 ;
  RECT 1320.220 192.850 1320.420 193.050 ;
  LAYER VI3 ;
  RECT 1319.820 193.250 1320.020 193.450 ;
  LAYER VI3 ;
  RECT 1319.820 192.850 1320.020 193.050 ;
  LAYER VI2 ;
  RECT 1319.820 192.790 1321.580 193.650 ;
  LAYER VI2 ;
  RECT 1321.020 193.250 1321.220 193.450 ;
  LAYER VI2 ;
  RECT 1321.020 192.850 1321.220 193.050 ;
  LAYER VI2 ;
  RECT 1320.620 193.250 1320.820 193.450 ;
  LAYER VI2 ;
  RECT 1320.620 192.850 1320.820 193.050 ;
  LAYER VI2 ;
  RECT 1320.220 193.250 1320.420 193.450 ;
  LAYER VI2 ;
  RECT 1320.220 192.850 1320.420 193.050 ;
  LAYER VI2 ;
  RECT 1319.820 193.250 1320.020 193.450 ;
  LAYER VI2 ;
  RECT 1319.820 192.850 1320.020 193.050 ;
  LAYER VI3 ;
  RECT 1323.820 192.790 1325.580 193.650 ;
  LAYER VI3 ;
  RECT 1325.020 193.250 1325.220 193.450 ;
  LAYER VI3 ;
  RECT 1325.020 192.850 1325.220 193.050 ;
  LAYER VI3 ;
  RECT 1324.620 193.250 1324.820 193.450 ;
  LAYER VI3 ;
  RECT 1324.620 192.850 1324.820 193.050 ;
  LAYER VI3 ;
  RECT 1324.220 193.250 1324.420 193.450 ;
  LAYER VI3 ;
  RECT 1324.220 192.850 1324.420 193.050 ;
  LAYER VI3 ;
  RECT 1323.820 193.250 1324.020 193.450 ;
  LAYER VI3 ;
  RECT 1323.820 192.850 1324.020 193.050 ;
  LAYER VI2 ;
  RECT 1323.820 192.790 1325.580 193.650 ;
  LAYER VI2 ;
  RECT 1325.020 193.250 1325.220 193.450 ;
  LAYER VI2 ;
  RECT 1325.020 192.850 1325.220 193.050 ;
  LAYER VI2 ;
  RECT 1324.620 193.250 1324.820 193.450 ;
  LAYER VI2 ;
  RECT 1324.620 192.850 1324.820 193.050 ;
  LAYER VI2 ;
  RECT 1324.220 193.250 1324.420 193.450 ;
  LAYER VI2 ;
  RECT 1324.220 192.850 1324.420 193.050 ;
  LAYER VI2 ;
  RECT 1323.820 193.250 1324.020 193.450 ;
  LAYER VI2 ;
  RECT 1323.820 192.850 1324.020 193.050 ;
  LAYER VI3 ;
  RECT 4.280 65.600 5.140 65.980 ;
  LAYER VI3 ;
  RECT 4.680 65.660 4.880 65.860 ;
  LAYER VI3 ;
  RECT 4.280 65.660 4.480 65.860 ;
  LAYER VI2 ;
  RECT 4.280 65.600 5.140 65.980 ;
  LAYER VI2 ;
  RECT 4.680 65.660 4.880 65.860 ;
  LAYER VI2 ;
  RECT 4.280 65.660 4.480 65.860 ;
  LAYER VI3 ;
  RECT 4.280 69.940 5.140 70.220 ;
  LAYER VI3 ;
  RECT 4.740 69.940 4.940 70.140 ;
  LAYER VI3 ;
  RECT 4.340 69.940 4.540 70.140 ;
  LAYER VI2 ;
  RECT 4.280 69.940 5.140 70.220 ;
  LAYER VI2 ;
  RECT 4.740 69.940 4.940 70.140 ;
  LAYER VI2 ;
  RECT 4.340 69.940 4.540 70.140 ;
  LAYER VI3 ;
  RECT 4.280 73.620 5.140 73.900 ;
  LAYER VI3 ;
  RECT 4.740 73.620 4.940 73.820 ;
  LAYER VI3 ;
  RECT 4.340 73.620 4.540 73.820 ;
  LAYER VI2 ;
  RECT 4.280 73.620 5.140 73.900 ;
  LAYER VI2 ;
  RECT 4.740 73.620 4.940 73.820 ;
  LAYER VI2 ;
  RECT 4.340 73.620 4.540 73.820 ;
  LAYER VI3 ;
  RECT 4.280 77.300 5.140 77.580 ;
  LAYER VI3 ;
  RECT 4.740 77.300 4.940 77.500 ;
  LAYER VI3 ;
  RECT 4.340 77.300 4.540 77.500 ;
  LAYER VI2 ;
  RECT 4.280 77.300 5.140 77.580 ;
  LAYER VI2 ;
  RECT 4.740 77.300 4.940 77.500 ;
  LAYER VI2 ;
  RECT 4.340 77.300 4.540 77.500 ;
  LAYER VI3 ;
  RECT 4.280 80.980 5.140 81.260 ;
  LAYER VI3 ;
  RECT 4.740 80.980 4.940 81.180 ;
  LAYER VI3 ;
  RECT 4.340 80.980 4.540 81.180 ;
  LAYER VI2 ;
  RECT 4.280 80.980 5.140 81.260 ;
  LAYER VI2 ;
  RECT 4.740 80.980 4.940 81.180 ;
  LAYER VI2 ;
  RECT 4.340 80.980 4.540 81.180 ;
  LAYER VI3 ;
  RECT 4.280 84.660 5.140 84.940 ;
  LAYER VI3 ;
  RECT 4.740 84.660 4.940 84.860 ;
  LAYER VI3 ;
  RECT 4.340 84.660 4.540 84.860 ;
  LAYER VI2 ;
  RECT 4.280 84.660 5.140 84.940 ;
  LAYER VI2 ;
  RECT 4.740 84.660 4.940 84.860 ;
  LAYER VI2 ;
  RECT 4.340 84.660 4.540 84.860 ;
  LAYER VI3 ;
  RECT 4.280 88.340 5.140 88.620 ;
  LAYER VI3 ;
  RECT 4.740 88.340 4.940 88.540 ;
  LAYER VI3 ;
  RECT 4.340 88.340 4.540 88.540 ;
  LAYER VI2 ;
  RECT 4.280 88.340 5.140 88.620 ;
  LAYER VI2 ;
  RECT 4.740 88.340 4.940 88.540 ;
  LAYER VI2 ;
  RECT 4.340 88.340 4.540 88.540 ;
  LAYER VI3 ;
  RECT 4.280 92.020 5.140 92.300 ;
  LAYER VI3 ;
  RECT 4.740 92.020 4.940 92.220 ;
  LAYER VI3 ;
  RECT 4.340 92.020 4.540 92.220 ;
  LAYER VI2 ;
  RECT 4.280 92.020 5.140 92.300 ;
  LAYER VI2 ;
  RECT 4.740 92.020 4.940 92.220 ;
  LAYER VI2 ;
  RECT 4.340 92.020 4.540 92.220 ;
  LAYER VI3 ;
  RECT 4.280 95.700 5.140 95.980 ;
  LAYER VI3 ;
  RECT 4.740 95.700 4.940 95.900 ;
  LAYER VI3 ;
  RECT 4.340 95.700 4.540 95.900 ;
  LAYER VI2 ;
  RECT 4.280 95.700 5.140 95.980 ;
  LAYER VI2 ;
  RECT 4.740 95.700 4.940 95.900 ;
  LAYER VI2 ;
  RECT 4.340 95.700 4.540 95.900 ;
  LAYER VI3 ;
  RECT 4.280 99.380 5.140 99.660 ;
  LAYER VI3 ;
  RECT 4.740 99.380 4.940 99.580 ;
  LAYER VI3 ;
  RECT 4.340 99.380 4.540 99.580 ;
  LAYER VI2 ;
  RECT 4.280 99.380 5.140 99.660 ;
  LAYER VI2 ;
  RECT 4.740 99.380 4.940 99.580 ;
  LAYER VI2 ;
  RECT 4.340 99.380 4.540 99.580 ;
  LAYER VI3 ;
  RECT 4.280 103.060 5.140 103.340 ;
  LAYER VI3 ;
  RECT 4.740 103.060 4.940 103.260 ;
  LAYER VI3 ;
  RECT 4.340 103.060 4.540 103.260 ;
  LAYER VI2 ;
  RECT 4.280 103.060 5.140 103.340 ;
  LAYER VI2 ;
  RECT 4.740 103.060 4.940 103.260 ;
  LAYER VI2 ;
  RECT 4.340 103.060 4.540 103.260 ;
  LAYER VI3 ;
  RECT 4.280 106.740 5.140 107.020 ;
  LAYER VI3 ;
  RECT 4.740 106.740 4.940 106.940 ;
  LAYER VI3 ;
  RECT 4.340 106.740 4.540 106.940 ;
  LAYER VI2 ;
  RECT 4.280 106.740 5.140 107.020 ;
  LAYER VI2 ;
  RECT 4.740 106.740 4.940 106.940 ;
  LAYER VI2 ;
  RECT 4.340 106.740 4.540 106.940 ;
  LAYER VI3 ;
  RECT 4.280 110.420 5.140 110.700 ;
  LAYER VI3 ;
  RECT 4.740 110.420 4.940 110.620 ;
  LAYER VI3 ;
  RECT 4.340 110.420 4.540 110.620 ;
  LAYER VI2 ;
  RECT 4.280 110.420 5.140 110.700 ;
  LAYER VI2 ;
  RECT 4.740 110.420 4.940 110.620 ;
  LAYER VI2 ;
  RECT 4.340 110.420 4.540 110.620 ;
  LAYER VI3 ;
  RECT 4.280 114.100 5.140 114.380 ;
  LAYER VI3 ;
  RECT 4.740 114.100 4.940 114.300 ;
  LAYER VI3 ;
  RECT 4.340 114.100 4.540 114.300 ;
  LAYER VI2 ;
  RECT 4.280 114.100 5.140 114.380 ;
  LAYER VI2 ;
  RECT 4.740 114.100 4.940 114.300 ;
  LAYER VI2 ;
  RECT 4.340 114.100 4.540 114.300 ;
  LAYER VI3 ;
  RECT 4.280 117.780 5.140 118.060 ;
  LAYER VI3 ;
  RECT 4.740 117.780 4.940 117.980 ;
  LAYER VI3 ;
  RECT 4.340 117.780 4.540 117.980 ;
  LAYER VI2 ;
  RECT 4.280 117.780 5.140 118.060 ;
  LAYER VI2 ;
  RECT 4.740 117.780 4.940 117.980 ;
  LAYER VI2 ;
  RECT 4.340 117.780 4.540 117.980 ;
  LAYER VI3 ;
  RECT 4.280 121.460 5.140 121.740 ;
  LAYER VI3 ;
  RECT 4.740 121.460 4.940 121.660 ;
  LAYER VI3 ;
  RECT 4.340 121.460 4.540 121.660 ;
  LAYER VI2 ;
  RECT 4.280 121.460 5.140 121.740 ;
  LAYER VI2 ;
  RECT 4.740 121.460 4.940 121.660 ;
  LAYER VI2 ;
  RECT 4.340 121.460 4.540 121.660 ;
  LAYER VI3 ;
  RECT 4.280 125.140 5.140 125.420 ;
  LAYER VI3 ;
  RECT 4.740 125.140 4.940 125.340 ;
  LAYER VI3 ;
  RECT 4.340 125.140 4.540 125.340 ;
  LAYER VI2 ;
  RECT 4.280 125.140 5.140 125.420 ;
  LAYER VI2 ;
  RECT 4.740 125.140 4.940 125.340 ;
  LAYER VI2 ;
  RECT 4.340 125.140 4.540 125.340 ;
  LAYER VI3 ;
  RECT 4.280 128.820 5.140 129.100 ;
  LAYER VI3 ;
  RECT 4.740 128.820 4.940 129.020 ;
  LAYER VI3 ;
  RECT 4.340 128.820 4.540 129.020 ;
  LAYER VI2 ;
  RECT 4.280 128.820 5.140 129.100 ;
  LAYER VI2 ;
  RECT 4.740 128.820 4.940 129.020 ;
  LAYER VI2 ;
  RECT 4.340 128.820 4.540 129.020 ;
  LAYER VI3 ;
  RECT 4.280 132.500 5.140 132.780 ;
  LAYER VI3 ;
  RECT 4.740 132.500 4.940 132.700 ;
  LAYER VI3 ;
  RECT 4.340 132.500 4.540 132.700 ;
  LAYER VI2 ;
  RECT 4.280 132.500 5.140 132.780 ;
  LAYER VI2 ;
  RECT 4.740 132.500 4.940 132.700 ;
  LAYER VI2 ;
  RECT 4.340 132.500 4.540 132.700 ;
  LAYER VI3 ;
  RECT 4.280 136.180 5.140 136.460 ;
  LAYER VI3 ;
  RECT 4.740 136.180 4.940 136.380 ;
  LAYER VI3 ;
  RECT 4.340 136.180 4.540 136.380 ;
  LAYER VI2 ;
  RECT 4.280 136.180 5.140 136.460 ;
  LAYER VI2 ;
  RECT 4.740 136.180 4.940 136.380 ;
  LAYER VI2 ;
  RECT 4.340 136.180 4.540 136.380 ;
  LAYER VI3 ;
  RECT 4.280 139.860 5.140 140.140 ;
  LAYER VI3 ;
  RECT 4.740 139.860 4.940 140.060 ;
  LAYER VI3 ;
  RECT 4.340 139.860 4.540 140.060 ;
  LAYER VI2 ;
  RECT 4.280 139.860 5.140 140.140 ;
  LAYER VI2 ;
  RECT 4.740 139.860 4.940 140.060 ;
  LAYER VI2 ;
  RECT 4.340 139.860 4.540 140.060 ;
  LAYER VI3 ;
  RECT 4.280 143.540 5.140 143.820 ;
  LAYER VI3 ;
  RECT 4.740 143.540 4.940 143.740 ;
  LAYER VI3 ;
  RECT 4.340 143.540 4.540 143.740 ;
  LAYER VI2 ;
  RECT 4.280 143.540 5.140 143.820 ;
  LAYER VI2 ;
  RECT 4.740 143.540 4.940 143.740 ;
  LAYER VI2 ;
  RECT 4.340 143.540 4.540 143.740 ;
  LAYER VI3 ;
  RECT 4.280 147.220 5.140 147.500 ;
  LAYER VI3 ;
  RECT 4.740 147.220 4.940 147.420 ;
  LAYER VI3 ;
  RECT 4.340 147.220 4.540 147.420 ;
  LAYER VI2 ;
  RECT 4.280 147.220 5.140 147.500 ;
  LAYER VI2 ;
  RECT 4.740 147.220 4.940 147.420 ;
  LAYER VI2 ;
  RECT 4.340 147.220 4.540 147.420 ;
  LAYER VI3 ;
  RECT 4.280 150.900 5.140 151.180 ;
  LAYER VI3 ;
  RECT 4.740 150.900 4.940 151.100 ;
  LAYER VI3 ;
  RECT 4.340 150.900 4.540 151.100 ;
  LAYER VI2 ;
  RECT 4.280 150.900 5.140 151.180 ;
  LAYER VI2 ;
  RECT 4.740 150.900 4.940 151.100 ;
  LAYER VI2 ;
  RECT 4.340 150.900 4.540 151.100 ;
  LAYER VI3 ;
  RECT 4.280 154.580 5.140 154.860 ;
  LAYER VI3 ;
  RECT 4.740 154.580 4.940 154.780 ;
  LAYER VI3 ;
  RECT 4.340 154.580 4.540 154.780 ;
  LAYER VI2 ;
  RECT 4.280 154.580 5.140 154.860 ;
  LAYER VI2 ;
  RECT 4.740 154.580 4.940 154.780 ;
  LAYER VI2 ;
  RECT 4.340 154.580 4.540 154.780 ;
  LAYER VI3 ;
  RECT 4.280 158.260 5.140 158.540 ;
  LAYER VI3 ;
  RECT 4.740 158.260 4.940 158.460 ;
  LAYER VI3 ;
  RECT 4.340 158.260 4.540 158.460 ;
  LAYER VI2 ;
  RECT 4.280 158.260 5.140 158.540 ;
  LAYER VI2 ;
  RECT 4.740 158.260 4.940 158.460 ;
  LAYER VI2 ;
  RECT 4.340 158.260 4.540 158.460 ;
  LAYER VI3 ;
  RECT 4.280 161.940 5.140 162.220 ;
  LAYER VI3 ;
  RECT 4.740 161.940 4.940 162.140 ;
  LAYER VI3 ;
  RECT 4.340 161.940 4.540 162.140 ;
  LAYER VI2 ;
  RECT 4.280 161.940 5.140 162.220 ;
  LAYER VI2 ;
  RECT 4.740 161.940 4.940 162.140 ;
  LAYER VI2 ;
  RECT 4.340 161.940 4.540 162.140 ;
  LAYER VI3 ;
  RECT 4.280 165.620 5.140 165.900 ;
  LAYER VI3 ;
  RECT 4.740 165.620 4.940 165.820 ;
  LAYER VI3 ;
  RECT 4.340 165.620 4.540 165.820 ;
  LAYER VI2 ;
  RECT 4.280 165.620 5.140 165.900 ;
  LAYER VI2 ;
  RECT 4.740 165.620 4.940 165.820 ;
  LAYER VI2 ;
  RECT 4.340 165.620 4.540 165.820 ;
  LAYER VI3 ;
  RECT 4.280 169.300 5.140 169.580 ;
  LAYER VI3 ;
  RECT 4.740 169.300 4.940 169.500 ;
  LAYER VI3 ;
  RECT 4.340 169.300 4.540 169.500 ;
  LAYER VI2 ;
  RECT 4.280 169.300 5.140 169.580 ;
  LAYER VI2 ;
  RECT 4.740 169.300 4.940 169.500 ;
  LAYER VI2 ;
  RECT 4.340 169.300 4.540 169.500 ;
  LAYER VI3 ;
  RECT 4.280 172.980 5.140 173.260 ;
  LAYER VI3 ;
  RECT 4.740 172.980 4.940 173.180 ;
  LAYER VI3 ;
  RECT 4.340 172.980 4.540 173.180 ;
  LAYER VI2 ;
  RECT 4.280 172.980 5.140 173.260 ;
  LAYER VI2 ;
  RECT 4.740 172.980 4.940 173.180 ;
  LAYER VI2 ;
  RECT 4.340 172.980 4.540 173.180 ;
  LAYER VI3 ;
  RECT 4.280 176.660 5.140 176.940 ;
  LAYER VI3 ;
  RECT 4.740 176.660 4.940 176.860 ;
  LAYER VI3 ;
  RECT 4.340 176.660 4.540 176.860 ;
  LAYER VI2 ;
  RECT 4.280 176.660 5.140 176.940 ;
  LAYER VI2 ;
  RECT 4.740 176.660 4.940 176.860 ;
  LAYER VI2 ;
  RECT 4.340 176.660 4.540 176.860 ;
  LAYER VI3 ;
  RECT 4.280 180.340 5.140 180.620 ;
  LAYER VI3 ;
  RECT 4.740 180.340 4.940 180.540 ;
  LAYER VI3 ;
  RECT 4.340 180.340 4.540 180.540 ;
  LAYER VI2 ;
  RECT 4.280 180.340 5.140 180.620 ;
  LAYER VI2 ;
  RECT 4.740 180.340 4.940 180.540 ;
  LAYER VI2 ;
  RECT 4.340 180.340 4.540 180.540 ;
  LAYER VI3 ;
  RECT 4.280 184.020 5.140 184.300 ;
  LAYER VI3 ;
  RECT 4.740 184.020 4.940 184.220 ;
  LAYER VI3 ;
  RECT 4.340 184.020 4.540 184.220 ;
  LAYER VI2 ;
  RECT 4.280 184.020 5.140 184.300 ;
  LAYER VI2 ;
  RECT 4.740 184.020 4.940 184.220 ;
  LAYER VI2 ;
  RECT 4.340 184.020 4.540 184.220 ;
  LAYER VI3 ;
  RECT 4.280 191.940 5.140 192.320 ;
  LAYER VI3 ;
  RECT 4.680 192.000 4.880 192.200 ;
  LAYER VI3 ;
  RECT 4.280 192.000 4.480 192.200 ;
  LAYER VI2 ;
  RECT 4.280 191.940 5.140 192.320 ;
  LAYER VI2 ;
  RECT 4.680 192.000 4.880 192.200 ;
  LAYER VI2 ;
  RECT 4.280 192.000 4.480 192.200 ;
  LAYER VI3 ;
  RECT 47.350 192.790 47.600 193.650 ;
  LAYER VI3 ;
  RECT 47.350 193.250 47.550 193.450 ;
  LAYER VI3 ;
  RECT 47.350 192.850 47.550 193.050 ;
  LAYER VI2 ;
  RECT 47.350 192.790 47.600 193.650 ;
  LAYER VI2 ;
  RECT 47.350 193.250 47.550 193.450 ;
  LAYER VI2 ;
  RECT 47.350 192.850 47.550 193.050 ;
  LAYER VI3 ;
  RECT 88.270 192.790 88.520 193.650 ;
  LAYER VI3 ;
  RECT 88.270 193.250 88.470 193.450 ;
  LAYER VI3 ;
  RECT 88.270 192.850 88.470 193.050 ;
  LAYER VI2 ;
  RECT 88.270 192.790 88.520 193.650 ;
  LAYER VI2 ;
  RECT 88.270 193.250 88.470 193.450 ;
  LAYER VI2 ;
  RECT 88.270 192.850 88.470 193.050 ;
  LAYER VI3 ;
  RECT 129.190 192.790 129.440 193.650 ;
  LAYER VI3 ;
  RECT 129.190 193.250 129.390 193.450 ;
  LAYER VI3 ;
  RECT 129.190 192.850 129.390 193.050 ;
  LAYER VI2 ;
  RECT 129.190 192.790 129.440 193.650 ;
  LAYER VI2 ;
  RECT 129.190 193.250 129.390 193.450 ;
  LAYER VI2 ;
  RECT 129.190 192.850 129.390 193.050 ;
  LAYER VI3 ;
  RECT 170.110 192.790 170.360 193.650 ;
  LAYER VI3 ;
  RECT 170.110 193.250 170.310 193.450 ;
  LAYER VI3 ;
  RECT 170.110 192.850 170.310 193.050 ;
  LAYER VI2 ;
  RECT 170.110 192.790 170.360 193.650 ;
  LAYER VI2 ;
  RECT 170.110 193.250 170.310 193.450 ;
  LAYER VI2 ;
  RECT 170.110 192.850 170.310 193.050 ;
  LAYER VI3 ;
  RECT 211.030 192.790 211.280 193.650 ;
  LAYER VI3 ;
  RECT 211.030 193.250 211.230 193.450 ;
  LAYER VI3 ;
  RECT 211.030 192.850 211.230 193.050 ;
  LAYER VI2 ;
  RECT 211.030 192.790 211.280 193.650 ;
  LAYER VI2 ;
  RECT 211.030 193.250 211.230 193.450 ;
  LAYER VI2 ;
  RECT 211.030 192.850 211.230 193.050 ;
  LAYER VI3 ;
  RECT 251.950 192.790 252.200 193.650 ;
  LAYER VI3 ;
  RECT 251.950 193.250 252.150 193.450 ;
  LAYER VI3 ;
  RECT 251.950 192.850 252.150 193.050 ;
  LAYER VI2 ;
  RECT 251.950 192.790 252.200 193.650 ;
  LAYER VI2 ;
  RECT 251.950 193.250 252.150 193.450 ;
  LAYER VI2 ;
  RECT 251.950 192.850 252.150 193.050 ;
  LAYER VI3 ;
  RECT 292.870 192.790 293.120 193.650 ;
  LAYER VI3 ;
  RECT 292.870 193.250 293.070 193.450 ;
  LAYER VI3 ;
  RECT 292.870 192.850 293.070 193.050 ;
  LAYER VI2 ;
  RECT 292.870 192.790 293.120 193.650 ;
  LAYER VI2 ;
  RECT 292.870 193.250 293.070 193.450 ;
  LAYER VI2 ;
  RECT 292.870 192.850 293.070 193.050 ;
  LAYER VI3 ;
  RECT 333.790 192.790 334.040 193.650 ;
  LAYER VI3 ;
  RECT 333.790 193.250 333.990 193.450 ;
  LAYER VI3 ;
  RECT 333.790 192.850 333.990 193.050 ;
  LAYER VI2 ;
  RECT 333.790 192.790 334.040 193.650 ;
  LAYER VI2 ;
  RECT 333.790 193.250 333.990 193.450 ;
  LAYER VI2 ;
  RECT 333.790 192.850 333.990 193.050 ;
  LAYER VI3 ;
  RECT 374.710 192.790 374.960 193.650 ;
  LAYER VI3 ;
  RECT 374.710 193.250 374.910 193.450 ;
  LAYER VI3 ;
  RECT 374.710 192.850 374.910 193.050 ;
  LAYER VI2 ;
  RECT 374.710 192.790 374.960 193.650 ;
  LAYER VI2 ;
  RECT 374.710 193.250 374.910 193.450 ;
  LAYER VI2 ;
  RECT 374.710 192.850 374.910 193.050 ;
  LAYER VI3 ;
  RECT 415.630 192.790 415.880 193.650 ;
  LAYER VI3 ;
  RECT 415.630 193.250 415.830 193.450 ;
  LAYER VI3 ;
  RECT 415.630 192.850 415.830 193.050 ;
  LAYER VI2 ;
  RECT 415.630 192.790 415.880 193.650 ;
  LAYER VI2 ;
  RECT 415.630 193.250 415.830 193.450 ;
  LAYER VI2 ;
  RECT 415.630 192.850 415.830 193.050 ;
  LAYER VI3 ;
  RECT 456.550 192.790 456.800 193.650 ;
  LAYER VI3 ;
  RECT 456.550 193.250 456.750 193.450 ;
  LAYER VI3 ;
  RECT 456.550 192.850 456.750 193.050 ;
  LAYER VI2 ;
  RECT 456.550 192.790 456.800 193.650 ;
  LAYER VI2 ;
  RECT 456.550 193.250 456.750 193.450 ;
  LAYER VI2 ;
  RECT 456.550 192.850 456.750 193.050 ;
  LAYER VI3 ;
  RECT 497.470 192.790 497.720 193.650 ;
  LAYER VI3 ;
  RECT 497.470 193.250 497.670 193.450 ;
  LAYER VI3 ;
  RECT 497.470 192.850 497.670 193.050 ;
  LAYER VI2 ;
  RECT 497.470 192.790 497.720 193.650 ;
  LAYER VI2 ;
  RECT 497.470 193.250 497.670 193.450 ;
  LAYER VI2 ;
  RECT 497.470 192.850 497.670 193.050 ;
  LAYER VI3 ;
  RECT 538.390 192.790 538.640 193.650 ;
  LAYER VI3 ;
  RECT 538.390 193.250 538.590 193.450 ;
  LAYER VI3 ;
  RECT 538.390 192.850 538.590 193.050 ;
  LAYER VI2 ;
  RECT 538.390 192.790 538.640 193.650 ;
  LAYER VI2 ;
  RECT 538.390 193.250 538.590 193.450 ;
  LAYER VI2 ;
  RECT 538.390 192.850 538.590 193.050 ;
  LAYER VI3 ;
  RECT 579.310 192.790 579.560 193.650 ;
  LAYER VI3 ;
  RECT 579.310 193.250 579.510 193.450 ;
  LAYER VI3 ;
  RECT 579.310 192.850 579.510 193.050 ;
  LAYER VI2 ;
  RECT 579.310 192.790 579.560 193.650 ;
  LAYER VI2 ;
  RECT 579.310 193.250 579.510 193.450 ;
  LAYER VI2 ;
  RECT 579.310 192.850 579.510 193.050 ;
  LAYER VI3 ;
  RECT 620.230 192.790 620.480 193.650 ;
  LAYER VI3 ;
  RECT 620.230 193.250 620.430 193.450 ;
  LAYER VI3 ;
  RECT 620.230 192.850 620.430 193.050 ;
  LAYER VI2 ;
  RECT 620.230 192.790 620.480 193.650 ;
  LAYER VI2 ;
  RECT 620.230 193.250 620.430 193.450 ;
  LAYER VI2 ;
  RECT 620.230 192.850 620.430 193.050 ;
  LAYER VI3 ;
  RECT 661.150 192.790 661.400 193.650 ;
  LAYER VI3 ;
  RECT 661.150 193.250 661.350 193.450 ;
  LAYER VI3 ;
  RECT 661.150 192.850 661.350 193.050 ;
  LAYER VI2 ;
  RECT 661.150 192.790 661.400 193.650 ;
  LAYER VI2 ;
  RECT 661.150 193.250 661.350 193.450 ;
  LAYER VI2 ;
  RECT 661.150 192.850 661.350 193.050 ;
  LAYER VI3 ;
  RECT 702.070 192.790 702.320 193.650 ;
  LAYER VI3 ;
  RECT 702.070 193.250 702.270 193.450 ;
  LAYER VI3 ;
  RECT 702.070 192.850 702.270 193.050 ;
  LAYER VI2 ;
  RECT 702.070 192.790 702.320 193.650 ;
  LAYER VI2 ;
  RECT 702.070 193.250 702.270 193.450 ;
  LAYER VI2 ;
  RECT 702.070 192.850 702.270 193.050 ;
  LAYER VI3 ;
  RECT 742.990 192.790 743.240 193.650 ;
  LAYER VI3 ;
  RECT 742.990 193.250 743.190 193.450 ;
  LAYER VI3 ;
  RECT 742.990 192.850 743.190 193.050 ;
  LAYER VI2 ;
  RECT 742.990 192.790 743.240 193.650 ;
  LAYER VI2 ;
  RECT 742.990 193.250 743.190 193.450 ;
  LAYER VI2 ;
  RECT 742.990 192.850 743.190 193.050 ;
  LAYER VI3 ;
  RECT 783.910 192.790 784.160 193.650 ;
  LAYER VI3 ;
  RECT 783.910 193.250 784.110 193.450 ;
  LAYER VI3 ;
  RECT 783.910 192.850 784.110 193.050 ;
  LAYER VI2 ;
  RECT 783.910 192.790 784.160 193.650 ;
  LAYER VI2 ;
  RECT 783.910 193.250 784.110 193.450 ;
  LAYER VI2 ;
  RECT 783.910 192.850 784.110 193.050 ;
  LAYER VI3 ;
  RECT 824.830 192.790 825.080 193.650 ;
  LAYER VI3 ;
  RECT 824.830 193.250 825.030 193.450 ;
  LAYER VI3 ;
  RECT 824.830 192.850 825.030 193.050 ;
  LAYER VI2 ;
  RECT 824.830 192.790 825.080 193.650 ;
  LAYER VI2 ;
  RECT 824.830 193.250 825.030 193.450 ;
  LAYER VI2 ;
  RECT 824.830 192.850 825.030 193.050 ;
  LAYER VI3 ;
  RECT 865.750 192.790 866.000 193.650 ;
  LAYER VI3 ;
  RECT 865.750 193.250 865.950 193.450 ;
  LAYER VI3 ;
  RECT 865.750 192.850 865.950 193.050 ;
  LAYER VI2 ;
  RECT 865.750 192.790 866.000 193.650 ;
  LAYER VI2 ;
  RECT 865.750 193.250 865.950 193.450 ;
  LAYER VI2 ;
  RECT 865.750 192.850 865.950 193.050 ;
  LAYER VI3 ;
  RECT 906.670 192.790 906.920 193.650 ;
  LAYER VI3 ;
  RECT 906.670 193.250 906.870 193.450 ;
  LAYER VI3 ;
  RECT 906.670 192.850 906.870 193.050 ;
  LAYER VI2 ;
  RECT 906.670 192.790 906.920 193.650 ;
  LAYER VI2 ;
  RECT 906.670 193.250 906.870 193.450 ;
  LAYER VI2 ;
  RECT 906.670 192.850 906.870 193.050 ;
  LAYER VI3 ;
  RECT 947.590 192.790 947.840 193.650 ;
  LAYER VI3 ;
  RECT 947.590 193.250 947.790 193.450 ;
  LAYER VI3 ;
  RECT 947.590 192.850 947.790 193.050 ;
  LAYER VI2 ;
  RECT 947.590 192.790 947.840 193.650 ;
  LAYER VI2 ;
  RECT 947.590 193.250 947.790 193.450 ;
  LAYER VI2 ;
  RECT 947.590 192.850 947.790 193.050 ;
  LAYER VI3 ;
  RECT 988.510 192.790 988.760 193.650 ;
  LAYER VI3 ;
  RECT 988.510 193.250 988.710 193.450 ;
  LAYER VI3 ;
  RECT 988.510 192.850 988.710 193.050 ;
  LAYER VI2 ;
  RECT 988.510 192.790 988.760 193.650 ;
  LAYER VI2 ;
  RECT 988.510 193.250 988.710 193.450 ;
  LAYER VI2 ;
  RECT 988.510 192.850 988.710 193.050 ;
  LAYER VI3 ;
  RECT 1029.430 192.790 1029.680 193.650 ;
  LAYER VI3 ;
  RECT 1029.430 193.250 1029.630 193.450 ;
  LAYER VI3 ;
  RECT 1029.430 192.850 1029.630 193.050 ;
  LAYER VI2 ;
  RECT 1029.430 192.790 1029.680 193.650 ;
  LAYER VI2 ;
  RECT 1029.430 193.250 1029.630 193.450 ;
  LAYER VI2 ;
  RECT 1029.430 192.850 1029.630 193.050 ;
  LAYER VI3 ;
  RECT 1070.350 192.790 1070.600 193.650 ;
  LAYER VI3 ;
  RECT 1070.350 193.250 1070.550 193.450 ;
  LAYER VI3 ;
  RECT 1070.350 192.850 1070.550 193.050 ;
  LAYER VI2 ;
  RECT 1070.350 192.790 1070.600 193.650 ;
  LAYER VI2 ;
  RECT 1070.350 193.250 1070.550 193.450 ;
  LAYER VI2 ;
  RECT 1070.350 192.850 1070.550 193.050 ;
  LAYER VI3 ;
  RECT 1111.270 192.790 1111.520 193.650 ;
  LAYER VI3 ;
  RECT 1111.270 193.250 1111.470 193.450 ;
  LAYER VI3 ;
  RECT 1111.270 192.850 1111.470 193.050 ;
  LAYER VI2 ;
  RECT 1111.270 192.790 1111.520 193.650 ;
  LAYER VI2 ;
  RECT 1111.270 193.250 1111.470 193.450 ;
  LAYER VI2 ;
  RECT 1111.270 192.850 1111.470 193.050 ;
  LAYER VI3 ;
  RECT 1152.190 192.790 1152.440 193.650 ;
  LAYER VI3 ;
  RECT 1152.190 193.250 1152.390 193.450 ;
  LAYER VI3 ;
  RECT 1152.190 192.850 1152.390 193.050 ;
  LAYER VI2 ;
  RECT 1152.190 192.790 1152.440 193.650 ;
  LAYER VI2 ;
  RECT 1152.190 193.250 1152.390 193.450 ;
  LAYER VI2 ;
  RECT 1152.190 192.850 1152.390 193.050 ;
  LAYER VI3 ;
  RECT 1193.110 192.790 1193.360 193.650 ;
  LAYER VI3 ;
  RECT 1193.110 193.250 1193.310 193.450 ;
  LAYER VI3 ;
  RECT 1193.110 192.850 1193.310 193.050 ;
  LAYER VI2 ;
  RECT 1193.110 192.790 1193.360 193.650 ;
  LAYER VI2 ;
  RECT 1193.110 193.250 1193.310 193.450 ;
  LAYER VI2 ;
  RECT 1193.110 192.850 1193.310 193.050 ;
  LAYER VI3 ;
  RECT 1234.030 192.790 1234.280 193.650 ;
  LAYER VI3 ;
  RECT 1234.030 193.250 1234.230 193.450 ;
  LAYER VI3 ;
  RECT 1234.030 192.850 1234.230 193.050 ;
  LAYER VI2 ;
  RECT 1234.030 192.790 1234.280 193.650 ;
  LAYER VI2 ;
  RECT 1234.030 193.250 1234.230 193.450 ;
  LAYER VI2 ;
  RECT 1234.030 192.850 1234.230 193.050 ;
  LAYER VI3 ;
  RECT 1274.950 192.790 1275.200 193.650 ;
  LAYER VI3 ;
  RECT 1274.950 193.250 1275.150 193.450 ;
  LAYER VI3 ;
  RECT 1274.950 192.850 1275.150 193.050 ;
  LAYER VI2 ;
  RECT 1274.950 192.790 1275.200 193.650 ;
  LAYER VI2 ;
  RECT 1274.950 193.250 1275.150 193.450 ;
  LAYER VI2 ;
  RECT 1274.950 192.850 1275.150 193.050 ;
END
END SHKD110_1024X16X8BM1
END LIBRARY





