# ________________________________________________________________________________________________
# 
# 
#             Synchronous One-Port Register File Compiler
# 
#                 UMC 0.11um LL AE Logic Process
# 
# ________________________________________________________________________________________________
# 
#               
#         Copyright (C) 2024 Faraday Technology Corporation. All Rights Reserved.       
#                
#         This source code is an unpublished work belongs to Faraday Technology Corporation       
#         It is considered a trade secret and is not to be divulged or       
#         used by parties who have not received written authorization from       
#         Faraday Technology Corporation       
#                
#         Faraday's home page can be found at: http://www.faraday-tech.com/       
#                
# ________________________________________________________________________________________________
# 
#        IP Name            :  FSR0K_B_SY                
#        IP Version         :  1.4.0                     
#        IP Release Status  :  Active                    
#        Word               :  256                       
#        Bit                :  9                         
#        Byte               :  8                         
#        Mux                :  4                         
#        Output Loading     :  0.01                      
#        Clock Input Slew   :  0.016                     
#        Data Input Slew    :  0.016                     
#        Ring Type          :  Ringless Model            
#        Ring Width         :  0                         
#        Bus Format         :  0                         
#        Memaker Path       :  /home/mem/Desktop/memlib  
#        GUI Version        :  m20230904                 
#        Date               :  2024/09/10 14:48:14       
# ________________________________________________________________________________________________
# 

VERSION 5.5 ;
NAMESCASESENSITIVE ON ;
MACRO SYKB110_256X9X8CM4
CLASS BLOCK ;
FOREIGN SYKB110_256X9X8CM4 0.000 0.000 ;
ORIGIN 0.000 0.000 ;
SIZE 620.075 BY 98.967 ;
SYMMETRY x y r90 ;
SITE core ;
PIN VCC
  DIRECTION INOUT ;
  USE POWER ;
 PORT
  LAYER ME4 ;
  RECT 333.521 0.000 334.241 33.870 ;
 END
 PORT
  LAYER ME4 ;
  RECT 329.517 0.000 330.237 33.870 ;
 END
 PORT
  LAYER ME4 ;
  RECT 341.529 0.000 342.249 33.870 ;
 END
 PORT
  LAYER ME4 ;
  RECT 337.525 0.000 338.245 33.870 ;
 END
 PORT
  LAYER ME4 ;
  RECT 349.537 0.000 350.257 33.870 ;
 END
 PORT
  LAYER ME4 ;
  RECT 345.533 0.000 346.253 33.870 ;
 END
 PORT
  LAYER ME4 ;
  RECT 357.545 0.000 358.265 33.870 ;
 END
 PORT
  LAYER ME4 ;
  RECT 353.541 0.000 354.261 33.870 ;
 END
 PORT
  LAYER ME4 ;
  RECT 365.553 0.000 366.273 33.870 ;
 END
 PORT
  LAYER ME4 ;
  RECT 361.549 0.000 362.269 33.870 ;
 END
 PORT
  LAYER ME4 ;
  RECT 373.561 0.000 374.281 33.870 ;
 END
 PORT
  LAYER ME4 ;
  RECT 369.557 0.000 370.277 33.870 ;
 END
 PORT
  LAYER ME4 ;
  RECT 381.569 0.000 382.289 33.870 ;
 END
 PORT
  LAYER ME4 ;
  RECT 377.565 0.000 378.285 33.870 ;
 END
 PORT
  LAYER ME4 ;
  RECT 389.577 0.000 390.297 33.870 ;
 END
 PORT
  LAYER ME4 ;
  RECT 385.573 0.000 386.293 33.870 ;
 END
 PORT
  LAYER ME4 ;
  RECT 397.585 0.000 398.305 33.870 ;
 END
 PORT
  LAYER ME4 ;
  RECT 393.581 0.000 394.301 33.870 ;
 END
 PORT
  LAYER ME4 ;
  RECT 405.593 0.000 406.313 33.870 ;
 END
 PORT
  LAYER ME4 ;
  RECT 401.589 0.000 402.309 33.870 ;
 END
 PORT
  LAYER ME4 ;
  RECT 413.601 0.000 414.321 33.870 ;
 END
 PORT
  LAYER ME4 ;
  RECT 409.597 0.000 410.317 33.870 ;
 END
 PORT
  LAYER ME4 ;
  RECT 421.609 0.000 422.329 33.870 ;
 END
 PORT
  LAYER ME4 ;
  RECT 417.605 0.000 418.325 33.870 ;
 END
 PORT
  LAYER ME4 ;
  RECT 429.617 0.000 430.337 33.870 ;
 END
 PORT
  LAYER ME4 ;
  RECT 425.613 0.000 426.333 33.870 ;
 END
 PORT
  LAYER ME4 ;
  RECT 437.625 0.000 438.345 33.870 ;
 END
 PORT
  LAYER ME4 ;
  RECT 433.621 0.000 434.341 33.870 ;
 END
 PORT
  LAYER ME4 ;
  RECT 445.633 0.000 446.353 33.870 ;
 END
 PORT
  LAYER ME4 ;
  RECT 441.629 0.000 442.349 33.870 ;
 END
 PORT
  LAYER ME4 ;
  RECT 453.641 0.000 454.361 33.870 ;
 END
 PORT
  LAYER ME4 ;
  RECT 449.637 0.000 450.357 33.870 ;
 END
 PORT
  LAYER ME4 ;
  RECT 461.649 0.000 462.369 33.870 ;
 END
 PORT
  LAYER ME4 ;
  RECT 457.645 0.000 458.365 33.870 ;
 END
 PORT
  LAYER ME4 ;
  RECT 469.657 0.000 470.377 33.870 ;
 END
 PORT
  LAYER ME4 ;
  RECT 465.653 0.000 466.373 33.870 ;
 END
 PORT
  LAYER ME4 ;
  RECT 477.665 0.000 478.385 33.870 ;
 END
 PORT
  LAYER ME4 ;
  RECT 473.661 0.000 474.381 33.870 ;
 END
 PORT
  LAYER ME4 ;
  RECT 485.673 0.000 486.393 33.870 ;
 END
 PORT
  LAYER ME4 ;
  RECT 481.669 0.000 482.389 33.870 ;
 END
 PORT
  LAYER ME4 ;
  RECT 493.681 0.000 494.401 33.870 ;
 END
 PORT
  LAYER ME4 ;
  RECT 489.677 0.000 490.397 33.870 ;
 END
 PORT
  LAYER ME4 ;
  RECT 501.689 0.000 502.409 33.870 ;
 END
 PORT
  LAYER ME4 ;
  RECT 497.685 0.000 498.405 33.870 ;
 END
 PORT
  LAYER ME4 ;
  RECT 509.697 0.000 510.417 33.870 ;
 END
 PORT
  LAYER ME4 ;
  RECT 505.693 0.000 506.413 33.870 ;
 END
 PORT
  LAYER ME4 ;
  RECT 517.705 0.000 518.425 33.870 ;
 END
 PORT
  LAYER ME4 ;
  RECT 513.701 0.000 514.421 33.870 ;
 END
 PORT
  LAYER ME4 ;
  RECT 525.713 0.000 526.433 33.870 ;
 END
 PORT
  LAYER ME4 ;
  RECT 521.709 0.000 522.429 33.870 ;
 END
 PORT
  LAYER ME4 ;
  RECT 533.721 0.000 534.441 33.870 ;
 END
 PORT
  LAYER ME4 ;
  RECT 529.717 0.000 530.437 33.870 ;
 END
 PORT
  LAYER ME4 ;
  RECT 541.729 0.000 542.449 33.870 ;
 END
 PORT
  LAYER ME4 ;
  RECT 537.725 0.000 538.445 33.870 ;
 END
 PORT
  LAYER ME4 ;
  RECT 549.737 0.000 550.457 33.870 ;
 END
 PORT
  LAYER ME4 ;
  RECT 545.733 0.000 546.453 33.870 ;
 END
 PORT
  LAYER ME4 ;
  RECT 557.745 0.000 558.465 33.870 ;
 END
 PORT
  LAYER ME4 ;
  RECT 553.741 0.000 554.461 33.870 ;
 END
 PORT
  LAYER ME4 ;
  RECT 565.753 0.000 566.473 33.870 ;
 END
 PORT
  LAYER ME4 ;
  RECT 561.749 0.000 562.469 33.870 ;
 END
 PORT
  LAYER ME4 ;
  RECT 573.761 0.000 574.481 33.870 ;
 END
 PORT
  LAYER ME4 ;
  RECT 569.757 0.000 570.477 33.870 ;
 END
 PORT
  LAYER ME4 ;
  RECT 581.769 0.000 582.489 33.870 ;
 END
 PORT
  LAYER ME4 ;
  RECT 577.765 0.000 578.485 33.870 ;
 END
 PORT
  LAYER ME4 ;
  RECT 589.777 0.000 590.497 33.870 ;
 END
 PORT
  LAYER ME4 ;
  RECT 585.773 0.000 586.493 33.870 ;
 END
 PORT
  LAYER ME4 ;
  RECT 597.785 0.000 598.505 33.870 ;
 END
 PORT
  LAYER ME4 ;
  RECT 593.781 0.000 594.501 33.870 ;
 END
 PORT
  LAYER ME4 ;
  RECT 605.793 0.000 606.513 33.870 ;
 END
 PORT
  LAYER ME4 ;
  RECT 601.789 0.000 602.509 33.870 ;
 END
 PORT
  LAYER ME4 ;
  RECT 613.801 0.000 614.521 33.870 ;
 END
 PORT
  LAYER ME4 ;
  RECT 609.797 0.000 610.517 33.870 ;
 END
 PORT
  LAYER ME4 ;
  RECT 618.775 0.000 619.155 98.967 ;
 END
 PORT
  LAYER ME4 ;
  RECT 312.629 0.000 313.229 98.967 ;
 END
 PORT
  LAYER ME4 ;
  RECT 316.809 0.000 317.529 98.967 ;
 END
 PORT
  LAYER ME4 ;
  RECT 318.919 0.000 320.039 98.967 ;
 END
 PORT
  LAYER ME4 ;
  RECT 324.949 0.000 325.669 98.967 ;
 END
 PORT
  LAYER ME4 ;
  RECT 326.885 0.921 327.265 98.967 ;
 END
 PORT
  LAYER ME4 ;
  RECT 305.684 0.000 306.804 98.967 ;
 END
 PORT
  LAYER ME4 ;
  RECT 308.399 0.000 309.119 98.967 ;
 END
 PORT
  LAYER ME4 ;
  RECT 303.310 0.000 304.030 98.208 ;
 END
 PORT
  LAYER ME4 ;
  RECT 301.270 0.921 301.990 98.967 ;
 END
 PORT
  LAYER ME4 ;
  RECT 299.150 0.000 299.870 98.967 ;
 END
 PORT
  LAYER ME4 ;
  RECT 297.110 0.921 297.830 98.967 ;
 END
 PORT
  LAYER ME4 ;
  RECT 0.920 0.000 1.300 98.967 ;
 END
 PORT
  LAYER ME4 ;
  RECT 7.556 0.000 8.276 33.870 ;
 END
 PORT
  LAYER ME4 ;
  RECT 3.552 0.000 4.272 33.870 ;
 END
 PORT
  LAYER ME4 ;
  RECT 15.564 0.000 16.284 33.870 ;
 END
 PORT
  LAYER ME4 ;
  RECT 11.560 0.000 12.280 33.870 ;
 END
 PORT
  LAYER ME4 ;
  RECT 23.572 0.000 24.292 33.870 ;
 END
 PORT
  LAYER ME4 ;
  RECT 19.568 0.000 20.288 33.870 ;
 END
 PORT
  LAYER ME4 ;
  RECT 31.580 0.000 32.300 33.870 ;
 END
 PORT
  LAYER ME4 ;
  RECT 27.576 0.000 28.296 33.870 ;
 END
 PORT
  LAYER ME4 ;
  RECT 39.588 0.000 40.308 33.870 ;
 END
 PORT
  LAYER ME4 ;
  RECT 35.584 0.000 36.304 33.870 ;
 END
 PORT
  LAYER ME4 ;
  RECT 47.596 0.000 48.316 33.870 ;
 END
 PORT
  LAYER ME4 ;
  RECT 43.592 0.000 44.312 33.870 ;
 END
 PORT
  LAYER ME4 ;
  RECT 55.604 0.000 56.324 33.870 ;
 END
 PORT
  LAYER ME4 ;
  RECT 51.600 0.000 52.320 33.870 ;
 END
 PORT
  LAYER ME4 ;
  RECT 63.612 0.000 64.332 33.870 ;
 END
 PORT
  LAYER ME4 ;
  RECT 59.608 0.000 60.328 33.870 ;
 END
 PORT
  LAYER ME4 ;
  RECT 71.620 0.000 72.340 33.870 ;
 END
 PORT
  LAYER ME4 ;
  RECT 67.616 0.000 68.336 33.870 ;
 END
 PORT
  LAYER ME4 ;
  RECT 79.628 0.000 80.348 33.870 ;
 END
 PORT
  LAYER ME4 ;
  RECT 75.624 0.000 76.344 33.870 ;
 END
 PORT
  LAYER ME4 ;
  RECT 87.636 0.000 88.356 33.870 ;
 END
 PORT
  LAYER ME4 ;
  RECT 83.632 0.000 84.352 33.870 ;
 END
 PORT
  LAYER ME4 ;
  RECT 95.644 0.000 96.364 33.870 ;
 END
 PORT
  LAYER ME4 ;
  RECT 91.640 0.000 92.360 33.870 ;
 END
 PORT
  LAYER ME4 ;
  RECT 103.652 0.000 104.372 33.870 ;
 END
 PORT
  LAYER ME4 ;
  RECT 99.648 0.000 100.368 33.870 ;
 END
 PORT
  LAYER ME4 ;
  RECT 111.660 0.000 112.380 33.870 ;
 END
 PORT
  LAYER ME4 ;
  RECT 107.656 0.000 108.376 33.870 ;
 END
 PORT
  LAYER ME4 ;
  RECT 119.668 0.000 120.388 33.870 ;
 END
 PORT
  LAYER ME4 ;
  RECT 115.664 0.000 116.384 33.870 ;
 END
 PORT
  LAYER ME4 ;
  RECT 127.676 0.000 128.396 33.870 ;
 END
 PORT
  LAYER ME4 ;
  RECT 123.672 0.000 124.392 33.870 ;
 END
 PORT
  LAYER ME4 ;
  RECT 135.684 0.000 136.404 33.870 ;
 END
 PORT
  LAYER ME4 ;
  RECT 131.680 0.000 132.400 33.870 ;
 END
 PORT
  LAYER ME4 ;
  RECT 143.692 0.000 144.412 33.870 ;
 END
 PORT
  LAYER ME4 ;
  RECT 139.688 0.000 140.408 33.870 ;
 END
 PORT
  LAYER ME4 ;
  RECT 151.700 0.000 152.420 33.870 ;
 END
 PORT
  LAYER ME4 ;
  RECT 147.696 0.000 148.416 33.870 ;
 END
 PORT
  LAYER ME4 ;
  RECT 159.708 0.000 160.428 33.870 ;
 END
 PORT
  LAYER ME4 ;
  RECT 155.704 0.000 156.424 33.870 ;
 END
 PORT
  LAYER ME4 ;
  RECT 167.716 0.000 168.436 33.870 ;
 END
 PORT
  LAYER ME4 ;
  RECT 163.712 0.000 164.432 33.870 ;
 END
 PORT
  LAYER ME4 ;
  RECT 175.724 0.000 176.444 33.870 ;
 END
 PORT
  LAYER ME4 ;
  RECT 171.720 0.000 172.440 33.870 ;
 END
 PORT
  LAYER ME4 ;
  RECT 183.732 0.000 184.452 33.870 ;
 END
 PORT
  LAYER ME4 ;
  RECT 179.728 0.000 180.448 33.870 ;
 END
 PORT
  LAYER ME4 ;
  RECT 191.740 0.000 192.460 33.870 ;
 END
 PORT
  LAYER ME4 ;
  RECT 187.736 0.000 188.456 33.870 ;
 END
 PORT
  LAYER ME4 ;
  RECT 199.748 0.000 200.468 33.870 ;
 END
 PORT
  LAYER ME4 ;
  RECT 195.744 0.000 196.464 33.870 ;
 END
 PORT
  LAYER ME4 ;
  RECT 207.756 0.000 208.476 33.870 ;
 END
 PORT
  LAYER ME4 ;
  RECT 203.752 0.000 204.472 33.870 ;
 END
 PORT
  LAYER ME4 ;
  RECT 215.764 0.000 216.484 33.870 ;
 END
 PORT
  LAYER ME4 ;
  RECT 211.760 0.000 212.480 33.870 ;
 END
 PORT
  LAYER ME4 ;
  RECT 223.772 0.000 224.492 33.870 ;
 END
 PORT
  LAYER ME4 ;
  RECT 219.768 0.000 220.488 33.870 ;
 END
 PORT
  LAYER ME4 ;
  RECT 231.780 0.000 232.500 33.870 ;
 END
 PORT
  LAYER ME4 ;
  RECT 227.776 0.000 228.496 33.870 ;
 END
 PORT
  LAYER ME4 ;
  RECT 239.788 0.000 240.508 33.870 ;
 END
 PORT
  LAYER ME4 ;
  RECT 235.784 0.000 236.504 33.870 ;
 END
 PORT
  LAYER ME4 ;
  RECT 247.796 0.000 248.516 33.870 ;
 END
 PORT
  LAYER ME4 ;
  RECT 243.792 0.000 244.512 33.870 ;
 END
 PORT
  LAYER ME4 ;
  RECT 255.804 0.000 256.524 33.870 ;
 END
 PORT
  LAYER ME4 ;
  RECT 251.800 0.000 252.520 33.870 ;
 END
 PORT
  LAYER ME4 ;
  RECT 263.812 0.000 264.532 33.870 ;
 END
 PORT
  LAYER ME4 ;
  RECT 259.808 0.000 260.528 33.870 ;
 END
 PORT
  LAYER ME4 ;
  RECT 271.820 0.000 272.540 33.870 ;
 END
 PORT
  LAYER ME4 ;
  RECT 267.816 0.000 268.536 33.870 ;
 END
 PORT
  LAYER ME4 ;
  RECT 279.828 0.000 280.548 33.870 ;
 END
 PORT
  LAYER ME4 ;
  RECT 275.824 0.000 276.544 33.870 ;
 END
 PORT
  LAYER ME4 ;
  RECT 287.836 0.000 288.556 33.870 ;
 END
 PORT
  LAYER ME4 ;
  RECT 283.832 0.000 284.552 33.870 ;
 END
 PORT
  LAYER ME4 ;
  RECT 294.990 0.000 295.710 98.967 ;
 END
 PORT
  LAYER ME4 ;
  RECT 292.810 0.000 293.190 98.967 ;
 END
 PORT
  LAYER ME4 ;
  RECT 335.713 35.220 336.053 98.967 ;
 END
 PORT
  LAYER ME4 ;
  RECT 333.711 35.220 334.051 98.967 ;
 END
 PORT
  LAYER ME4 ;
  RECT 331.709 35.220 332.049 98.967 ;
 END
 PORT
  LAYER ME4 ;
  RECT 329.707 35.220 330.047 98.967 ;
 END
 PORT
  LAYER ME4 ;
  RECT 343.721 35.220 344.061 98.967 ;
 END
 PORT
  LAYER ME4 ;
  RECT 341.719 35.220 342.059 98.967 ;
 END
 PORT
  LAYER ME4 ;
  RECT 339.717 35.220 340.057 98.967 ;
 END
 PORT
  LAYER ME4 ;
  RECT 337.715 35.220 338.055 98.967 ;
 END
 PORT
  LAYER ME4 ;
  RECT 351.729 35.220 352.069 98.967 ;
 END
 PORT
  LAYER ME4 ;
  RECT 349.727 35.220 350.067 98.967 ;
 END
 PORT
  LAYER ME4 ;
  RECT 347.725 35.220 348.065 98.967 ;
 END
 PORT
  LAYER ME4 ;
  RECT 345.723 35.220 346.063 98.967 ;
 END
 PORT
  LAYER ME4 ;
  RECT 359.737 35.220 360.077 98.967 ;
 END
 PORT
  LAYER ME4 ;
  RECT 357.735 35.220 358.075 98.967 ;
 END
 PORT
  LAYER ME4 ;
  RECT 355.733 35.220 356.073 98.967 ;
 END
 PORT
  LAYER ME4 ;
  RECT 353.731 35.220 354.071 98.967 ;
 END
 PORT
  LAYER ME4 ;
  RECT 367.745 35.220 368.085 98.967 ;
 END
 PORT
  LAYER ME4 ;
  RECT 365.743 35.220 366.083 98.967 ;
 END
 PORT
  LAYER ME4 ;
  RECT 363.741 35.220 364.081 98.967 ;
 END
 PORT
  LAYER ME4 ;
  RECT 361.739 35.220 362.079 98.967 ;
 END
 PORT
  LAYER ME4 ;
  RECT 375.753 35.220 376.093 98.967 ;
 END
 PORT
  LAYER ME4 ;
  RECT 373.751 35.220 374.091 98.967 ;
 END
 PORT
  LAYER ME4 ;
  RECT 371.749 35.220 372.089 98.967 ;
 END
 PORT
  LAYER ME4 ;
  RECT 369.747 35.220 370.087 98.967 ;
 END
 PORT
  LAYER ME4 ;
  RECT 383.761 35.220 384.101 98.967 ;
 END
 PORT
  LAYER ME4 ;
  RECT 381.759 35.220 382.099 98.967 ;
 END
 PORT
  LAYER ME4 ;
  RECT 379.757 35.220 380.097 98.967 ;
 END
 PORT
  LAYER ME4 ;
  RECT 377.755 35.220 378.095 98.967 ;
 END
 PORT
  LAYER ME4 ;
  RECT 391.769 35.220 392.109 98.967 ;
 END
 PORT
  LAYER ME4 ;
  RECT 389.767 35.220 390.107 98.967 ;
 END
 PORT
  LAYER ME4 ;
  RECT 387.765 35.220 388.105 98.967 ;
 END
 PORT
  LAYER ME4 ;
  RECT 385.763 35.220 386.103 98.967 ;
 END
 PORT
  LAYER ME4 ;
  RECT 399.777 35.220 400.117 98.967 ;
 END
 PORT
  LAYER ME4 ;
  RECT 397.775 35.220 398.115 98.967 ;
 END
 PORT
  LAYER ME4 ;
  RECT 395.773 35.220 396.113 98.967 ;
 END
 PORT
  LAYER ME4 ;
  RECT 393.771 35.220 394.111 98.967 ;
 END
 PORT
  LAYER ME4 ;
  RECT 407.785 35.220 408.125 98.967 ;
 END
 PORT
  LAYER ME4 ;
  RECT 405.783 35.220 406.123 98.967 ;
 END
 PORT
  LAYER ME4 ;
  RECT 403.781 35.220 404.121 98.967 ;
 END
 PORT
  LAYER ME4 ;
  RECT 401.779 35.220 402.119 98.967 ;
 END
 PORT
  LAYER ME4 ;
  RECT 415.793 35.220 416.133 98.967 ;
 END
 PORT
  LAYER ME4 ;
  RECT 413.791 35.220 414.131 98.967 ;
 END
 PORT
  LAYER ME4 ;
  RECT 411.789 35.220 412.129 98.967 ;
 END
 PORT
  LAYER ME4 ;
  RECT 409.787 35.220 410.127 98.967 ;
 END
 PORT
  LAYER ME4 ;
  RECT 423.801 35.220 424.141 98.967 ;
 END
 PORT
  LAYER ME4 ;
  RECT 421.799 35.220 422.139 98.967 ;
 END
 PORT
  LAYER ME4 ;
  RECT 419.797 35.220 420.137 98.967 ;
 END
 PORT
  LAYER ME4 ;
  RECT 417.795 35.220 418.135 98.967 ;
 END
 PORT
  LAYER ME4 ;
  RECT 431.809 35.220 432.149 98.967 ;
 END
 PORT
  LAYER ME4 ;
  RECT 429.807 35.220 430.147 98.967 ;
 END
 PORT
  LAYER ME4 ;
  RECT 427.805 35.220 428.145 98.967 ;
 END
 PORT
  LAYER ME4 ;
  RECT 425.803 35.220 426.143 98.967 ;
 END
 PORT
  LAYER ME4 ;
  RECT 439.817 35.220 440.157 98.967 ;
 END
 PORT
  LAYER ME4 ;
  RECT 437.815 35.220 438.155 98.967 ;
 END
 PORT
  LAYER ME4 ;
  RECT 435.813 35.220 436.153 98.967 ;
 END
 PORT
  LAYER ME4 ;
  RECT 433.811 35.220 434.151 98.967 ;
 END
 PORT
  LAYER ME4 ;
  RECT 447.825 35.220 448.165 98.967 ;
 END
 PORT
  LAYER ME4 ;
  RECT 445.823 35.220 446.163 98.967 ;
 END
 PORT
  LAYER ME4 ;
  RECT 443.821 35.220 444.161 98.967 ;
 END
 PORT
  LAYER ME4 ;
  RECT 441.819 35.220 442.159 98.967 ;
 END
 PORT
  LAYER ME4 ;
  RECT 455.833 35.220 456.173 98.967 ;
 END
 PORT
  LAYER ME4 ;
  RECT 453.831 35.220 454.171 98.967 ;
 END
 PORT
  LAYER ME4 ;
  RECT 451.829 35.220 452.169 98.967 ;
 END
 PORT
  LAYER ME4 ;
  RECT 449.827 35.220 450.167 98.967 ;
 END
 PORT
  LAYER ME4 ;
  RECT 463.841 35.220 464.181 98.967 ;
 END
 PORT
  LAYER ME4 ;
  RECT 461.839 35.220 462.179 98.967 ;
 END
 PORT
  LAYER ME4 ;
  RECT 459.837 35.220 460.177 98.967 ;
 END
 PORT
  LAYER ME4 ;
  RECT 457.835 35.220 458.175 98.967 ;
 END
 PORT
  LAYER ME4 ;
  RECT 471.849 35.220 472.189 98.967 ;
 END
 PORT
  LAYER ME4 ;
  RECT 469.847 35.220 470.187 98.967 ;
 END
 PORT
  LAYER ME4 ;
  RECT 467.845 35.220 468.185 98.967 ;
 END
 PORT
  LAYER ME4 ;
  RECT 465.843 35.220 466.183 98.967 ;
 END
 PORT
  LAYER ME4 ;
  RECT 479.857 35.220 480.197 98.967 ;
 END
 PORT
  LAYER ME4 ;
  RECT 477.855 35.220 478.195 98.967 ;
 END
 PORT
  LAYER ME4 ;
  RECT 475.853 35.220 476.193 98.967 ;
 END
 PORT
  LAYER ME4 ;
  RECT 473.851 35.220 474.191 98.967 ;
 END
 PORT
  LAYER ME4 ;
  RECT 487.865 35.220 488.205 98.967 ;
 END
 PORT
  LAYER ME4 ;
  RECT 485.863 35.220 486.203 98.967 ;
 END
 PORT
  LAYER ME4 ;
  RECT 483.861 35.220 484.201 98.967 ;
 END
 PORT
  LAYER ME4 ;
  RECT 481.859 35.220 482.199 98.967 ;
 END
 PORT
  LAYER ME4 ;
  RECT 495.873 35.220 496.213 98.967 ;
 END
 PORT
  LAYER ME4 ;
  RECT 493.871 35.220 494.211 98.967 ;
 END
 PORT
  LAYER ME4 ;
  RECT 491.869 35.220 492.209 98.967 ;
 END
 PORT
  LAYER ME4 ;
  RECT 489.867 35.220 490.207 98.967 ;
 END
 PORT
  LAYER ME4 ;
  RECT 503.881 35.220 504.221 98.967 ;
 END
 PORT
  LAYER ME4 ;
  RECT 501.879 35.220 502.219 98.967 ;
 END
 PORT
  LAYER ME4 ;
  RECT 499.877 35.220 500.217 98.967 ;
 END
 PORT
  LAYER ME4 ;
  RECT 497.875 35.220 498.215 98.967 ;
 END
 PORT
  LAYER ME4 ;
  RECT 511.889 35.220 512.229 98.967 ;
 END
 PORT
  LAYER ME4 ;
  RECT 509.887 35.220 510.227 98.967 ;
 END
 PORT
  LAYER ME4 ;
  RECT 507.885 35.220 508.225 98.967 ;
 END
 PORT
  LAYER ME4 ;
  RECT 505.883 35.220 506.223 98.967 ;
 END
 PORT
  LAYER ME4 ;
  RECT 519.897 35.220 520.237 98.967 ;
 END
 PORT
  LAYER ME4 ;
  RECT 517.895 35.220 518.235 98.967 ;
 END
 PORT
  LAYER ME4 ;
  RECT 515.893 35.220 516.233 98.967 ;
 END
 PORT
  LAYER ME4 ;
  RECT 513.891 35.220 514.231 98.967 ;
 END
 PORT
  LAYER ME4 ;
  RECT 527.905 35.220 528.245 98.967 ;
 END
 PORT
  LAYER ME4 ;
  RECT 525.903 35.220 526.243 98.967 ;
 END
 PORT
  LAYER ME4 ;
  RECT 523.901 35.220 524.241 98.967 ;
 END
 PORT
  LAYER ME4 ;
  RECT 521.899 35.220 522.239 98.967 ;
 END
 PORT
  LAYER ME4 ;
  RECT 535.913 35.220 536.253 98.967 ;
 END
 PORT
  LAYER ME4 ;
  RECT 533.911 35.220 534.251 98.967 ;
 END
 PORT
  LAYER ME4 ;
  RECT 531.909 35.220 532.249 98.967 ;
 END
 PORT
  LAYER ME4 ;
  RECT 529.907 35.220 530.247 98.967 ;
 END
 PORT
  LAYER ME4 ;
  RECT 543.921 35.220 544.261 98.967 ;
 END
 PORT
  LAYER ME4 ;
  RECT 541.919 35.220 542.259 98.967 ;
 END
 PORT
  LAYER ME4 ;
  RECT 539.917 35.220 540.257 98.967 ;
 END
 PORT
  LAYER ME4 ;
  RECT 537.915 35.220 538.255 98.967 ;
 END
 PORT
  LAYER ME4 ;
  RECT 551.929 35.220 552.269 98.967 ;
 END
 PORT
  LAYER ME4 ;
  RECT 549.927 35.220 550.267 98.967 ;
 END
 PORT
  LAYER ME4 ;
  RECT 547.925 35.220 548.265 98.967 ;
 END
 PORT
  LAYER ME4 ;
  RECT 545.923 35.220 546.263 98.967 ;
 END
 PORT
  LAYER ME4 ;
  RECT 559.937 35.220 560.277 98.967 ;
 END
 PORT
  LAYER ME4 ;
  RECT 557.935 35.220 558.275 98.967 ;
 END
 PORT
  LAYER ME4 ;
  RECT 555.933 35.220 556.273 98.967 ;
 END
 PORT
  LAYER ME4 ;
  RECT 553.931 35.220 554.271 98.967 ;
 END
 PORT
  LAYER ME4 ;
  RECT 567.945 35.220 568.285 98.967 ;
 END
 PORT
  LAYER ME4 ;
  RECT 565.943 35.220 566.283 98.967 ;
 END
 PORT
  LAYER ME4 ;
  RECT 563.941 35.220 564.281 98.967 ;
 END
 PORT
  LAYER ME4 ;
  RECT 561.939 35.220 562.279 98.967 ;
 END
 PORT
  LAYER ME4 ;
  RECT 575.953 35.220 576.293 98.967 ;
 END
 PORT
  LAYER ME4 ;
  RECT 573.951 35.220 574.291 98.967 ;
 END
 PORT
  LAYER ME4 ;
  RECT 571.949 35.220 572.289 98.967 ;
 END
 PORT
  LAYER ME4 ;
  RECT 569.947 35.220 570.287 98.967 ;
 END
 PORT
  LAYER ME4 ;
  RECT 583.961 35.220 584.301 98.967 ;
 END
 PORT
  LAYER ME4 ;
  RECT 581.959 35.220 582.299 98.967 ;
 END
 PORT
  LAYER ME4 ;
  RECT 579.957 35.220 580.297 98.967 ;
 END
 PORT
  LAYER ME4 ;
  RECT 577.955 35.220 578.295 98.967 ;
 END
 PORT
  LAYER ME4 ;
  RECT 591.969 35.220 592.309 98.967 ;
 END
 PORT
  LAYER ME4 ;
  RECT 589.967 35.220 590.307 98.967 ;
 END
 PORT
  LAYER ME4 ;
  RECT 587.965 35.220 588.305 98.967 ;
 END
 PORT
  LAYER ME4 ;
  RECT 585.963 35.220 586.303 98.967 ;
 END
 PORT
  LAYER ME4 ;
  RECT 599.977 35.220 600.317 98.967 ;
 END
 PORT
  LAYER ME4 ;
  RECT 597.975 35.220 598.315 98.967 ;
 END
 PORT
  LAYER ME4 ;
  RECT 595.973 35.220 596.313 98.967 ;
 END
 PORT
  LAYER ME4 ;
  RECT 593.971 35.220 594.311 98.967 ;
 END
 PORT
  LAYER ME4 ;
  RECT 607.985 35.220 608.325 98.967 ;
 END
 PORT
  LAYER ME4 ;
  RECT 605.983 35.220 606.323 98.967 ;
 END
 PORT
  LAYER ME4 ;
  RECT 603.981 35.220 604.321 98.967 ;
 END
 PORT
  LAYER ME4 ;
  RECT 601.979 35.220 602.319 98.967 ;
 END
 PORT
  LAYER ME4 ;
  RECT 615.993 35.220 616.333 98.967 ;
 END
 PORT
  LAYER ME4 ;
  RECT 613.991 35.220 614.331 98.967 ;
 END
 PORT
  LAYER ME4 ;
  RECT 611.989 35.220 612.329 98.967 ;
 END
 PORT
  LAYER ME4 ;
  RECT 609.987 35.220 610.327 98.967 ;
 END
 PORT
  LAYER ME4 ;
  RECT 9.748 35.220 10.088 98.967 ;
 END
 PORT
  LAYER ME4 ;
  RECT 7.746 35.220 8.086 98.967 ;
 END
 PORT
  LAYER ME4 ;
  RECT 5.744 35.220 6.084 98.967 ;
 END
 PORT
  LAYER ME4 ;
  RECT 3.742 35.220 4.082 98.967 ;
 END
 PORT
  LAYER ME4 ;
  RECT 17.756 35.220 18.096 98.967 ;
 END
 PORT
  LAYER ME4 ;
  RECT 15.754 35.220 16.094 98.967 ;
 END
 PORT
  LAYER ME4 ;
  RECT 13.752 35.220 14.092 98.967 ;
 END
 PORT
  LAYER ME4 ;
  RECT 11.750 35.220 12.090 98.967 ;
 END
 PORT
  LAYER ME4 ;
  RECT 25.764 35.220 26.104 98.967 ;
 END
 PORT
  LAYER ME4 ;
  RECT 23.762 35.220 24.102 98.967 ;
 END
 PORT
  LAYER ME4 ;
  RECT 21.760 35.220 22.100 98.967 ;
 END
 PORT
  LAYER ME4 ;
  RECT 19.758 35.220 20.098 98.967 ;
 END
 PORT
  LAYER ME4 ;
  RECT 33.772 35.220 34.112 98.967 ;
 END
 PORT
  LAYER ME4 ;
  RECT 31.770 35.220 32.110 98.967 ;
 END
 PORT
  LAYER ME4 ;
  RECT 29.768 35.220 30.108 98.967 ;
 END
 PORT
  LAYER ME4 ;
  RECT 27.766 35.220 28.106 98.967 ;
 END
 PORT
  LAYER ME4 ;
  RECT 41.780 35.220 42.120 98.967 ;
 END
 PORT
  LAYER ME4 ;
  RECT 39.778 35.220 40.118 98.967 ;
 END
 PORT
  LAYER ME4 ;
  RECT 37.776 35.220 38.116 98.967 ;
 END
 PORT
  LAYER ME4 ;
  RECT 35.774 35.220 36.114 98.967 ;
 END
 PORT
  LAYER ME4 ;
  RECT 49.788 35.220 50.128 98.967 ;
 END
 PORT
  LAYER ME4 ;
  RECT 47.786 35.220 48.126 98.967 ;
 END
 PORT
  LAYER ME4 ;
  RECT 45.784 35.220 46.124 98.967 ;
 END
 PORT
  LAYER ME4 ;
  RECT 43.782 35.220 44.122 98.967 ;
 END
 PORT
  LAYER ME4 ;
  RECT 57.796 35.220 58.136 98.967 ;
 END
 PORT
  LAYER ME4 ;
  RECT 55.794 35.220 56.134 98.967 ;
 END
 PORT
  LAYER ME4 ;
  RECT 53.792 35.220 54.132 98.967 ;
 END
 PORT
  LAYER ME4 ;
  RECT 51.790 35.220 52.130 98.967 ;
 END
 PORT
  LAYER ME4 ;
  RECT 65.804 35.220 66.144 98.967 ;
 END
 PORT
  LAYER ME4 ;
  RECT 63.802 35.220 64.142 98.967 ;
 END
 PORT
  LAYER ME4 ;
  RECT 61.800 35.220 62.140 98.967 ;
 END
 PORT
  LAYER ME4 ;
  RECT 59.798 35.220 60.138 98.967 ;
 END
 PORT
  LAYER ME4 ;
  RECT 73.812 35.220 74.152 98.967 ;
 END
 PORT
  LAYER ME4 ;
  RECT 71.810 35.220 72.150 98.967 ;
 END
 PORT
  LAYER ME4 ;
  RECT 69.808 35.220 70.148 98.967 ;
 END
 PORT
  LAYER ME4 ;
  RECT 67.806 35.220 68.146 98.967 ;
 END
 PORT
  LAYER ME4 ;
  RECT 81.820 35.220 82.160 98.967 ;
 END
 PORT
  LAYER ME4 ;
  RECT 79.818 35.220 80.158 98.967 ;
 END
 PORT
  LAYER ME4 ;
  RECT 77.816 35.220 78.156 98.967 ;
 END
 PORT
  LAYER ME4 ;
  RECT 75.814 35.220 76.154 98.967 ;
 END
 PORT
  LAYER ME4 ;
  RECT 89.828 35.220 90.168 98.967 ;
 END
 PORT
  LAYER ME4 ;
  RECT 87.826 35.220 88.166 98.967 ;
 END
 PORT
  LAYER ME4 ;
  RECT 85.824 35.220 86.164 98.967 ;
 END
 PORT
  LAYER ME4 ;
  RECT 83.822 35.220 84.162 98.967 ;
 END
 PORT
  LAYER ME4 ;
  RECT 97.836 35.220 98.176 98.967 ;
 END
 PORT
  LAYER ME4 ;
  RECT 95.834 35.220 96.174 98.967 ;
 END
 PORT
  LAYER ME4 ;
  RECT 93.832 35.220 94.172 98.967 ;
 END
 PORT
  LAYER ME4 ;
  RECT 91.830 35.220 92.170 98.967 ;
 END
 PORT
  LAYER ME4 ;
  RECT 105.844 35.220 106.184 98.967 ;
 END
 PORT
  LAYER ME4 ;
  RECT 103.842 35.220 104.182 98.967 ;
 END
 PORT
  LAYER ME4 ;
  RECT 101.840 35.220 102.180 98.967 ;
 END
 PORT
  LAYER ME4 ;
  RECT 99.838 35.220 100.178 98.967 ;
 END
 PORT
  LAYER ME4 ;
  RECT 113.852 35.220 114.192 98.967 ;
 END
 PORT
  LAYER ME4 ;
  RECT 111.850 35.220 112.190 98.967 ;
 END
 PORT
  LAYER ME4 ;
  RECT 109.848 35.220 110.188 98.967 ;
 END
 PORT
  LAYER ME4 ;
  RECT 107.846 35.220 108.186 98.967 ;
 END
 PORT
  LAYER ME4 ;
  RECT 121.860 35.220 122.200 98.967 ;
 END
 PORT
  LAYER ME4 ;
  RECT 119.858 35.220 120.198 98.967 ;
 END
 PORT
  LAYER ME4 ;
  RECT 117.856 35.220 118.196 98.967 ;
 END
 PORT
  LAYER ME4 ;
  RECT 115.854 35.220 116.194 98.967 ;
 END
 PORT
  LAYER ME4 ;
  RECT 129.868 35.220 130.208 98.967 ;
 END
 PORT
  LAYER ME4 ;
  RECT 127.866 35.220 128.206 98.967 ;
 END
 PORT
  LAYER ME4 ;
  RECT 125.864 35.220 126.204 98.967 ;
 END
 PORT
  LAYER ME4 ;
  RECT 123.862 35.220 124.202 98.967 ;
 END
 PORT
  LAYER ME4 ;
  RECT 137.876 35.220 138.216 98.967 ;
 END
 PORT
  LAYER ME4 ;
  RECT 135.874 35.220 136.214 98.967 ;
 END
 PORT
  LAYER ME4 ;
  RECT 133.872 35.220 134.212 98.967 ;
 END
 PORT
  LAYER ME4 ;
  RECT 131.870 35.220 132.210 98.967 ;
 END
 PORT
  LAYER ME4 ;
  RECT 145.884 35.220 146.224 98.967 ;
 END
 PORT
  LAYER ME4 ;
  RECT 143.882 35.220 144.222 98.967 ;
 END
 PORT
  LAYER ME4 ;
  RECT 141.880 35.220 142.220 98.967 ;
 END
 PORT
  LAYER ME4 ;
  RECT 139.878 35.220 140.218 98.967 ;
 END
 PORT
  LAYER ME4 ;
  RECT 153.892 35.220 154.232 98.967 ;
 END
 PORT
  LAYER ME4 ;
  RECT 151.890 35.220 152.230 98.967 ;
 END
 PORT
  LAYER ME4 ;
  RECT 149.888 35.220 150.228 98.967 ;
 END
 PORT
  LAYER ME4 ;
  RECT 147.886 35.220 148.226 98.967 ;
 END
 PORT
  LAYER ME4 ;
  RECT 161.900 35.220 162.240 98.967 ;
 END
 PORT
  LAYER ME4 ;
  RECT 159.898 35.220 160.238 98.967 ;
 END
 PORT
  LAYER ME4 ;
  RECT 157.896 35.220 158.236 98.967 ;
 END
 PORT
  LAYER ME4 ;
  RECT 155.894 35.220 156.234 98.967 ;
 END
 PORT
  LAYER ME4 ;
  RECT 169.908 35.220 170.248 98.967 ;
 END
 PORT
  LAYER ME4 ;
  RECT 167.906 35.220 168.246 98.967 ;
 END
 PORT
  LAYER ME4 ;
  RECT 165.904 35.220 166.244 98.967 ;
 END
 PORT
  LAYER ME4 ;
  RECT 163.902 35.220 164.242 98.967 ;
 END
 PORT
  LAYER ME4 ;
  RECT 177.916 35.220 178.256 98.967 ;
 END
 PORT
  LAYER ME4 ;
  RECT 175.914 35.220 176.254 98.967 ;
 END
 PORT
  LAYER ME4 ;
  RECT 173.912 35.220 174.252 98.967 ;
 END
 PORT
  LAYER ME4 ;
  RECT 171.910 35.220 172.250 98.967 ;
 END
 PORT
  LAYER ME4 ;
  RECT 185.924 35.220 186.264 98.967 ;
 END
 PORT
  LAYER ME4 ;
  RECT 183.922 35.220 184.262 98.967 ;
 END
 PORT
  LAYER ME4 ;
  RECT 181.920 35.220 182.260 98.967 ;
 END
 PORT
  LAYER ME4 ;
  RECT 179.918 35.220 180.258 98.967 ;
 END
 PORT
  LAYER ME4 ;
  RECT 193.932 35.220 194.272 98.967 ;
 END
 PORT
  LAYER ME4 ;
  RECT 191.930 35.220 192.270 98.967 ;
 END
 PORT
  LAYER ME4 ;
  RECT 189.928 35.220 190.268 98.967 ;
 END
 PORT
  LAYER ME4 ;
  RECT 187.926 35.220 188.266 98.967 ;
 END
 PORT
  LAYER ME4 ;
  RECT 201.940 35.220 202.280 98.967 ;
 END
 PORT
  LAYER ME4 ;
  RECT 199.938 35.220 200.278 98.967 ;
 END
 PORT
  LAYER ME4 ;
  RECT 197.936 35.220 198.276 98.967 ;
 END
 PORT
  LAYER ME4 ;
  RECT 195.934 35.220 196.274 98.967 ;
 END
 PORT
  LAYER ME4 ;
  RECT 209.948 35.220 210.288 98.967 ;
 END
 PORT
  LAYER ME4 ;
  RECT 207.946 35.220 208.286 98.967 ;
 END
 PORT
  LAYER ME4 ;
  RECT 205.944 35.220 206.284 98.967 ;
 END
 PORT
  LAYER ME4 ;
  RECT 203.942 35.220 204.282 98.967 ;
 END
 PORT
  LAYER ME4 ;
  RECT 217.956 35.220 218.296 98.967 ;
 END
 PORT
  LAYER ME4 ;
  RECT 215.954 35.220 216.294 98.967 ;
 END
 PORT
  LAYER ME4 ;
  RECT 213.952 35.220 214.292 98.967 ;
 END
 PORT
  LAYER ME4 ;
  RECT 211.950 35.220 212.290 98.967 ;
 END
 PORT
  LAYER ME4 ;
  RECT 225.964 35.220 226.304 98.967 ;
 END
 PORT
  LAYER ME4 ;
  RECT 223.962 35.220 224.302 98.967 ;
 END
 PORT
  LAYER ME4 ;
  RECT 221.960 35.220 222.300 98.967 ;
 END
 PORT
  LAYER ME4 ;
  RECT 219.958 35.220 220.298 98.967 ;
 END
 PORT
  LAYER ME4 ;
  RECT 233.972 35.220 234.312 98.967 ;
 END
 PORT
  LAYER ME4 ;
  RECT 231.970 35.220 232.310 98.967 ;
 END
 PORT
  LAYER ME4 ;
  RECT 229.968 35.220 230.308 98.967 ;
 END
 PORT
  LAYER ME4 ;
  RECT 227.966 35.220 228.306 98.967 ;
 END
 PORT
  LAYER ME4 ;
  RECT 241.980 35.220 242.320 98.967 ;
 END
 PORT
  LAYER ME4 ;
  RECT 239.978 35.220 240.318 98.967 ;
 END
 PORT
  LAYER ME4 ;
  RECT 237.976 35.220 238.316 98.967 ;
 END
 PORT
  LAYER ME4 ;
  RECT 235.974 35.220 236.314 98.967 ;
 END
 PORT
  LAYER ME4 ;
  RECT 249.988 35.220 250.328 98.967 ;
 END
 PORT
  LAYER ME4 ;
  RECT 247.986 35.220 248.326 98.967 ;
 END
 PORT
  LAYER ME4 ;
  RECT 245.984 35.220 246.324 98.967 ;
 END
 PORT
  LAYER ME4 ;
  RECT 243.982 35.220 244.322 98.967 ;
 END
 PORT
  LAYER ME4 ;
  RECT 257.996 35.220 258.336 98.967 ;
 END
 PORT
  LAYER ME4 ;
  RECT 255.994 35.220 256.334 98.967 ;
 END
 PORT
  LAYER ME4 ;
  RECT 253.992 35.220 254.332 98.967 ;
 END
 PORT
  LAYER ME4 ;
  RECT 251.990 35.220 252.330 98.967 ;
 END
 PORT
  LAYER ME4 ;
  RECT 266.004 35.220 266.344 98.967 ;
 END
 PORT
  LAYER ME4 ;
  RECT 264.002 35.220 264.342 98.967 ;
 END
 PORT
  LAYER ME4 ;
  RECT 262.000 35.220 262.340 98.967 ;
 END
 PORT
  LAYER ME4 ;
  RECT 259.998 35.220 260.338 98.967 ;
 END
 PORT
  LAYER ME4 ;
  RECT 274.012 35.220 274.352 98.967 ;
 END
 PORT
  LAYER ME4 ;
  RECT 272.010 35.220 272.350 98.967 ;
 END
 PORT
  LAYER ME4 ;
  RECT 270.008 35.220 270.348 98.967 ;
 END
 PORT
  LAYER ME4 ;
  RECT 268.006 35.220 268.346 98.967 ;
 END
 PORT
  LAYER ME4 ;
  RECT 282.020 35.220 282.360 98.967 ;
 END
 PORT
  LAYER ME4 ;
  RECT 280.018 35.220 280.358 98.967 ;
 END
 PORT
  LAYER ME4 ;
  RECT 278.016 35.220 278.356 98.967 ;
 END
 PORT
  LAYER ME4 ;
  RECT 276.014 35.220 276.354 98.967 ;
 END
 PORT
  LAYER ME4 ;
  RECT 290.028 35.220 290.368 98.967 ;
 END
 PORT
  LAYER ME4 ;
  RECT 288.026 35.220 288.366 98.967 ;
 END
 PORT
  LAYER ME4 ;
  RECT 286.024 35.220 286.364 98.967 ;
 END
 PORT
  LAYER ME4 ;
  RECT 284.022 35.220 284.362 98.967 ;
 END
END VCC
PIN GND
  DIRECTION INOUT ;
  USE GROUND ;
 PORT
  LAYER ME4 ;
  RECT 328.706 0.921 329.046 98.967 ;
 END
 PORT
  LAYER ME4 ;
  RECT 335.523 0.000 336.243 31.570 ;
 END
 PORT
  LAYER ME4 ;
  RECT 336.714 0.000 337.054 98.967 ;
 END
 PORT
  LAYER ME4 ;
  RECT 330.708 0.000 331.048 98.967 ;
 END
 PORT
  LAYER ME4 ;
  RECT 331.519 0.000 332.239 31.570 ;
 END
 PORT
  LAYER ME4 ;
  RECT 332.710 0.921 333.050 98.967 ;
 END
 PORT
  LAYER ME4 ;
  RECT 334.712 0.921 335.052 98.967 ;
 END
 PORT
  LAYER ME4 ;
  RECT 343.531 0.000 344.251 31.570 ;
 END
 PORT
  LAYER ME4 ;
  RECT 344.722 0.000 345.062 98.967 ;
 END
 PORT
  LAYER ME4 ;
  RECT 338.716 0.000 339.056 98.967 ;
 END
 PORT
  LAYER ME4 ;
  RECT 339.527 0.000 340.247 31.570 ;
 END
 PORT
  LAYER ME4 ;
  RECT 340.718 0.921 341.058 98.967 ;
 END
 PORT
  LAYER ME4 ;
  RECT 342.720 0.921 343.060 98.967 ;
 END
 PORT
  LAYER ME4 ;
  RECT 351.539 0.000 352.259 31.570 ;
 END
 PORT
  LAYER ME4 ;
  RECT 352.730 0.000 353.070 98.967 ;
 END
 PORT
  LAYER ME4 ;
  RECT 346.724 0.000 347.064 98.967 ;
 END
 PORT
  LAYER ME4 ;
  RECT 347.535 0.000 348.255 31.570 ;
 END
 PORT
  LAYER ME4 ;
  RECT 348.726 0.921 349.066 98.967 ;
 END
 PORT
  LAYER ME4 ;
  RECT 350.728 0.921 351.068 98.967 ;
 END
 PORT
  LAYER ME4 ;
  RECT 359.547 0.000 360.267 31.570 ;
 END
 PORT
  LAYER ME4 ;
  RECT 360.738 0.000 361.078 98.967 ;
 END
 PORT
  LAYER ME4 ;
  RECT 354.732 0.000 355.072 98.967 ;
 END
 PORT
  LAYER ME4 ;
  RECT 355.543 0.000 356.263 31.570 ;
 END
 PORT
  LAYER ME4 ;
  RECT 356.734 0.921 357.074 98.967 ;
 END
 PORT
  LAYER ME4 ;
  RECT 358.736 0.921 359.076 98.967 ;
 END
 PORT
  LAYER ME4 ;
  RECT 367.555 0.000 368.275 31.570 ;
 END
 PORT
  LAYER ME4 ;
  RECT 368.746 0.000 369.086 98.967 ;
 END
 PORT
  LAYER ME4 ;
  RECT 362.740 0.000 363.080 98.967 ;
 END
 PORT
  LAYER ME4 ;
  RECT 363.551 0.000 364.271 31.570 ;
 END
 PORT
  LAYER ME4 ;
  RECT 364.742 0.921 365.082 98.967 ;
 END
 PORT
  LAYER ME4 ;
  RECT 366.744 0.921 367.084 98.967 ;
 END
 PORT
  LAYER ME4 ;
  RECT 375.563 0.000 376.283 31.570 ;
 END
 PORT
  LAYER ME4 ;
  RECT 376.754 0.000 377.094 98.967 ;
 END
 PORT
  LAYER ME4 ;
  RECT 370.748 0.000 371.088 98.967 ;
 END
 PORT
  LAYER ME4 ;
  RECT 371.559 0.000 372.279 31.570 ;
 END
 PORT
  LAYER ME4 ;
  RECT 372.750 0.921 373.090 98.967 ;
 END
 PORT
  LAYER ME4 ;
  RECT 374.752 0.921 375.092 98.967 ;
 END
 PORT
  LAYER ME4 ;
  RECT 383.571 0.000 384.291 31.570 ;
 END
 PORT
  LAYER ME4 ;
  RECT 384.762 0.000 385.102 98.967 ;
 END
 PORT
  LAYER ME4 ;
  RECT 378.756 0.000 379.096 98.967 ;
 END
 PORT
  LAYER ME4 ;
  RECT 379.567 0.000 380.287 31.570 ;
 END
 PORT
  LAYER ME4 ;
  RECT 380.758 0.921 381.098 98.967 ;
 END
 PORT
  LAYER ME4 ;
  RECT 382.760 0.921 383.100 98.967 ;
 END
 PORT
  LAYER ME4 ;
  RECT 391.579 0.000 392.299 31.570 ;
 END
 PORT
  LAYER ME4 ;
  RECT 392.770 0.000 393.110 98.967 ;
 END
 PORT
  LAYER ME4 ;
  RECT 386.764 0.000 387.104 98.967 ;
 END
 PORT
  LAYER ME4 ;
  RECT 387.575 0.000 388.295 31.570 ;
 END
 PORT
  LAYER ME4 ;
  RECT 388.766 0.921 389.106 98.967 ;
 END
 PORT
  LAYER ME4 ;
  RECT 390.768 0.921 391.108 98.967 ;
 END
 PORT
  LAYER ME4 ;
  RECT 399.587 0.000 400.307 31.570 ;
 END
 PORT
  LAYER ME4 ;
  RECT 400.778 0.000 401.118 98.967 ;
 END
 PORT
  LAYER ME4 ;
  RECT 394.772 0.000 395.112 98.967 ;
 END
 PORT
  LAYER ME4 ;
  RECT 395.583 0.000 396.303 31.570 ;
 END
 PORT
  LAYER ME4 ;
  RECT 396.774 0.921 397.114 98.967 ;
 END
 PORT
  LAYER ME4 ;
  RECT 398.776 0.921 399.116 98.967 ;
 END
 PORT
  LAYER ME4 ;
  RECT 407.595 0.000 408.315 31.570 ;
 END
 PORT
  LAYER ME4 ;
  RECT 408.786 0.000 409.126 98.967 ;
 END
 PORT
  LAYER ME4 ;
  RECT 402.780 0.000 403.120 98.967 ;
 END
 PORT
  LAYER ME4 ;
  RECT 403.591 0.000 404.311 31.570 ;
 END
 PORT
  LAYER ME4 ;
  RECT 404.782 0.921 405.122 98.967 ;
 END
 PORT
  LAYER ME4 ;
  RECT 406.784 0.921 407.124 98.967 ;
 END
 PORT
  LAYER ME4 ;
  RECT 415.603 0.000 416.323 31.570 ;
 END
 PORT
  LAYER ME4 ;
  RECT 416.794 0.000 417.134 98.967 ;
 END
 PORT
  LAYER ME4 ;
  RECT 410.788 0.000 411.128 98.967 ;
 END
 PORT
  LAYER ME4 ;
  RECT 411.599 0.000 412.319 31.570 ;
 END
 PORT
  LAYER ME4 ;
  RECT 412.790 0.921 413.130 98.967 ;
 END
 PORT
  LAYER ME4 ;
  RECT 414.792 0.921 415.132 98.967 ;
 END
 PORT
  LAYER ME4 ;
  RECT 423.611 0.000 424.331 31.570 ;
 END
 PORT
  LAYER ME4 ;
  RECT 424.802 0.000 425.142 98.967 ;
 END
 PORT
  LAYER ME4 ;
  RECT 418.796 0.000 419.136 98.967 ;
 END
 PORT
  LAYER ME4 ;
  RECT 419.607 0.000 420.327 31.570 ;
 END
 PORT
  LAYER ME4 ;
  RECT 420.798 0.921 421.138 98.967 ;
 END
 PORT
  LAYER ME4 ;
  RECT 422.800 0.921 423.140 98.967 ;
 END
 PORT
  LAYER ME4 ;
  RECT 431.619 0.000 432.339 31.570 ;
 END
 PORT
  LAYER ME4 ;
  RECT 432.810 0.000 433.150 98.967 ;
 END
 PORT
  LAYER ME4 ;
  RECT 426.804 0.000 427.144 98.967 ;
 END
 PORT
  LAYER ME4 ;
  RECT 427.615 0.000 428.335 31.570 ;
 END
 PORT
  LAYER ME4 ;
  RECT 428.806 0.921 429.146 98.967 ;
 END
 PORT
  LAYER ME4 ;
  RECT 430.808 0.921 431.148 98.967 ;
 END
 PORT
  LAYER ME4 ;
  RECT 439.627 0.000 440.347 31.570 ;
 END
 PORT
  LAYER ME4 ;
  RECT 440.818 0.000 441.158 98.967 ;
 END
 PORT
  LAYER ME4 ;
  RECT 434.812 0.000 435.152 98.967 ;
 END
 PORT
  LAYER ME4 ;
  RECT 435.623 0.000 436.343 31.570 ;
 END
 PORT
  LAYER ME4 ;
  RECT 436.814 0.921 437.154 98.967 ;
 END
 PORT
  LAYER ME4 ;
  RECT 438.816 0.921 439.156 98.967 ;
 END
 PORT
  LAYER ME4 ;
  RECT 447.635 0.000 448.355 31.570 ;
 END
 PORT
  LAYER ME4 ;
  RECT 448.826 0.000 449.166 98.967 ;
 END
 PORT
  LAYER ME4 ;
  RECT 442.820 0.000 443.160 98.967 ;
 END
 PORT
  LAYER ME4 ;
  RECT 443.631 0.000 444.351 31.570 ;
 END
 PORT
  LAYER ME4 ;
  RECT 444.822 0.921 445.162 98.967 ;
 END
 PORT
  LAYER ME4 ;
  RECT 446.824 0.921 447.164 98.967 ;
 END
 PORT
  LAYER ME4 ;
  RECT 455.643 0.000 456.363 31.570 ;
 END
 PORT
  LAYER ME4 ;
  RECT 456.834 0.000 457.174 98.967 ;
 END
 PORT
  LAYER ME4 ;
  RECT 450.828 0.000 451.168 98.967 ;
 END
 PORT
  LAYER ME4 ;
  RECT 451.639 0.000 452.359 31.570 ;
 END
 PORT
  LAYER ME4 ;
  RECT 452.830 0.921 453.170 98.967 ;
 END
 PORT
  LAYER ME4 ;
  RECT 454.832 0.921 455.172 98.967 ;
 END
 PORT
  LAYER ME4 ;
  RECT 463.651 0.000 464.371 31.570 ;
 END
 PORT
  LAYER ME4 ;
  RECT 464.842 0.000 465.182 98.967 ;
 END
 PORT
  LAYER ME4 ;
  RECT 458.836 0.000 459.176 98.967 ;
 END
 PORT
  LAYER ME4 ;
  RECT 459.647 0.000 460.367 31.570 ;
 END
 PORT
  LAYER ME4 ;
  RECT 460.838 0.921 461.178 98.967 ;
 END
 PORT
  LAYER ME4 ;
  RECT 462.840 0.921 463.180 98.967 ;
 END
 PORT
  LAYER ME4 ;
  RECT 471.659 0.000 472.379 31.570 ;
 END
 PORT
  LAYER ME4 ;
  RECT 472.850 0.000 473.190 98.967 ;
 END
 PORT
  LAYER ME4 ;
  RECT 466.844 0.000 467.184 98.967 ;
 END
 PORT
  LAYER ME4 ;
  RECT 467.655 0.000 468.375 31.570 ;
 END
 PORT
  LAYER ME4 ;
  RECT 468.846 0.921 469.186 98.967 ;
 END
 PORT
  LAYER ME4 ;
  RECT 470.848 0.921 471.188 98.967 ;
 END
 PORT
  LAYER ME4 ;
  RECT 479.667 0.000 480.387 31.570 ;
 END
 PORT
  LAYER ME4 ;
  RECT 480.858 0.000 481.198 98.967 ;
 END
 PORT
  LAYER ME4 ;
  RECT 474.852 0.000 475.192 98.967 ;
 END
 PORT
  LAYER ME4 ;
  RECT 475.663 0.000 476.383 31.570 ;
 END
 PORT
  LAYER ME4 ;
  RECT 476.854 0.921 477.194 98.967 ;
 END
 PORT
  LAYER ME4 ;
  RECT 478.856 0.921 479.196 98.967 ;
 END
 PORT
  LAYER ME4 ;
  RECT 487.675 0.000 488.395 31.570 ;
 END
 PORT
  LAYER ME4 ;
  RECT 488.866 0.000 489.206 98.967 ;
 END
 PORT
  LAYER ME4 ;
  RECT 482.860 0.000 483.200 98.967 ;
 END
 PORT
  LAYER ME4 ;
  RECT 483.671 0.000 484.391 31.570 ;
 END
 PORT
  LAYER ME4 ;
  RECT 484.862 0.921 485.202 98.967 ;
 END
 PORT
  LAYER ME4 ;
  RECT 486.864 0.921 487.204 98.967 ;
 END
 PORT
  LAYER ME4 ;
  RECT 495.683 0.000 496.403 31.570 ;
 END
 PORT
  LAYER ME4 ;
  RECT 496.874 0.000 497.214 98.967 ;
 END
 PORT
  LAYER ME4 ;
  RECT 490.868 0.000 491.208 98.967 ;
 END
 PORT
  LAYER ME4 ;
  RECT 491.679 0.000 492.399 31.570 ;
 END
 PORT
  LAYER ME4 ;
  RECT 492.870 0.921 493.210 98.967 ;
 END
 PORT
  LAYER ME4 ;
  RECT 494.872 0.921 495.212 98.967 ;
 END
 PORT
  LAYER ME4 ;
  RECT 503.691 0.000 504.411 31.570 ;
 END
 PORT
  LAYER ME4 ;
  RECT 504.882 0.000 505.222 98.967 ;
 END
 PORT
  LAYER ME4 ;
  RECT 498.876 0.000 499.216 98.967 ;
 END
 PORT
  LAYER ME4 ;
  RECT 499.687 0.000 500.407 31.570 ;
 END
 PORT
  LAYER ME4 ;
  RECT 500.878 0.921 501.218 98.967 ;
 END
 PORT
  LAYER ME4 ;
  RECT 502.880 0.921 503.220 98.967 ;
 END
 PORT
  LAYER ME4 ;
  RECT 511.699 0.000 512.419 31.570 ;
 END
 PORT
  LAYER ME4 ;
  RECT 512.890 0.000 513.230 98.967 ;
 END
 PORT
  LAYER ME4 ;
  RECT 506.884 0.000 507.224 98.967 ;
 END
 PORT
  LAYER ME4 ;
  RECT 507.695 0.000 508.415 31.570 ;
 END
 PORT
  LAYER ME4 ;
  RECT 508.886 0.921 509.226 98.967 ;
 END
 PORT
  LAYER ME4 ;
  RECT 510.888 0.921 511.228 98.967 ;
 END
 PORT
  LAYER ME4 ;
  RECT 519.707 0.000 520.427 31.570 ;
 END
 PORT
  LAYER ME4 ;
  RECT 520.898 0.000 521.238 98.967 ;
 END
 PORT
  LAYER ME4 ;
  RECT 514.892 0.000 515.232 98.967 ;
 END
 PORT
  LAYER ME4 ;
  RECT 515.703 0.000 516.423 31.570 ;
 END
 PORT
  LAYER ME4 ;
  RECT 516.894 0.921 517.234 98.967 ;
 END
 PORT
  LAYER ME4 ;
  RECT 518.896 0.921 519.236 98.967 ;
 END
 PORT
  LAYER ME4 ;
  RECT 527.715 0.000 528.435 31.570 ;
 END
 PORT
  LAYER ME4 ;
  RECT 528.906 0.000 529.246 98.967 ;
 END
 PORT
  LAYER ME4 ;
  RECT 522.900 0.000 523.240 98.967 ;
 END
 PORT
  LAYER ME4 ;
  RECT 523.711 0.000 524.431 31.570 ;
 END
 PORT
  LAYER ME4 ;
  RECT 524.902 0.921 525.242 98.967 ;
 END
 PORT
  LAYER ME4 ;
  RECT 526.904 0.921 527.244 98.967 ;
 END
 PORT
  LAYER ME4 ;
  RECT 535.723 0.000 536.443 31.570 ;
 END
 PORT
  LAYER ME4 ;
  RECT 536.914 0.000 537.254 98.967 ;
 END
 PORT
  LAYER ME4 ;
  RECT 530.908 0.000 531.248 98.967 ;
 END
 PORT
  LAYER ME4 ;
  RECT 531.719 0.000 532.439 31.570 ;
 END
 PORT
  LAYER ME4 ;
  RECT 532.910 0.921 533.250 98.967 ;
 END
 PORT
  LAYER ME4 ;
  RECT 534.912 0.921 535.252 98.967 ;
 END
 PORT
  LAYER ME4 ;
  RECT 543.731 0.000 544.451 31.570 ;
 END
 PORT
  LAYER ME4 ;
  RECT 544.922 0.000 545.262 98.967 ;
 END
 PORT
  LAYER ME4 ;
  RECT 538.916 0.000 539.256 98.967 ;
 END
 PORT
  LAYER ME4 ;
  RECT 539.727 0.000 540.447 31.570 ;
 END
 PORT
  LAYER ME4 ;
  RECT 540.918 0.921 541.258 98.967 ;
 END
 PORT
  LAYER ME4 ;
  RECT 542.920 0.921 543.260 98.967 ;
 END
 PORT
  LAYER ME4 ;
  RECT 551.739 0.000 552.459 31.570 ;
 END
 PORT
  LAYER ME4 ;
  RECT 552.930 0.000 553.270 98.967 ;
 END
 PORT
  LAYER ME4 ;
  RECT 546.924 0.000 547.264 98.967 ;
 END
 PORT
  LAYER ME4 ;
  RECT 547.735 0.000 548.455 31.570 ;
 END
 PORT
  LAYER ME4 ;
  RECT 548.926 0.921 549.266 98.967 ;
 END
 PORT
  LAYER ME4 ;
  RECT 550.928 0.921 551.268 98.967 ;
 END
 PORT
  LAYER ME4 ;
  RECT 559.747 0.000 560.467 31.570 ;
 END
 PORT
  LAYER ME4 ;
  RECT 560.938 0.000 561.278 98.967 ;
 END
 PORT
  LAYER ME4 ;
  RECT 554.932 0.000 555.272 98.967 ;
 END
 PORT
  LAYER ME4 ;
  RECT 555.743 0.000 556.463 31.570 ;
 END
 PORT
  LAYER ME4 ;
  RECT 556.934 0.921 557.274 98.967 ;
 END
 PORT
  LAYER ME4 ;
  RECT 558.936 0.921 559.276 98.967 ;
 END
 PORT
  LAYER ME4 ;
  RECT 567.755 0.000 568.475 31.570 ;
 END
 PORT
  LAYER ME4 ;
  RECT 568.946 0.000 569.286 98.967 ;
 END
 PORT
  LAYER ME4 ;
  RECT 562.940 0.000 563.280 98.967 ;
 END
 PORT
  LAYER ME4 ;
  RECT 563.751 0.000 564.471 31.570 ;
 END
 PORT
  LAYER ME4 ;
  RECT 564.942 0.921 565.282 98.967 ;
 END
 PORT
  LAYER ME4 ;
  RECT 566.944 0.921 567.284 98.967 ;
 END
 PORT
  LAYER ME4 ;
  RECT 575.763 0.000 576.483 31.570 ;
 END
 PORT
  LAYER ME4 ;
  RECT 576.954 0.000 577.294 98.967 ;
 END
 PORT
  LAYER ME4 ;
  RECT 570.948 0.000 571.288 98.967 ;
 END
 PORT
  LAYER ME4 ;
  RECT 571.759 0.000 572.479 31.570 ;
 END
 PORT
  LAYER ME4 ;
  RECT 572.950 0.921 573.290 98.967 ;
 END
 PORT
  LAYER ME4 ;
  RECT 574.952 0.921 575.292 98.967 ;
 END
 PORT
  LAYER ME4 ;
  RECT 583.771 0.000 584.491 31.570 ;
 END
 PORT
  LAYER ME4 ;
  RECT 584.962 0.000 585.302 98.967 ;
 END
 PORT
  LAYER ME4 ;
  RECT 578.956 0.000 579.296 98.967 ;
 END
 PORT
  LAYER ME4 ;
  RECT 579.767 0.000 580.487 31.570 ;
 END
 PORT
  LAYER ME4 ;
  RECT 580.958 0.921 581.298 98.967 ;
 END
 PORT
  LAYER ME4 ;
  RECT 582.960 0.921 583.300 98.967 ;
 END
 PORT
  LAYER ME4 ;
  RECT 591.779 0.000 592.499 31.570 ;
 END
 PORT
  LAYER ME4 ;
  RECT 592.970 0.000 593.310 98.967 ;
 END
 PORT
  LAYER ME4 ;
  RECT 586.964 0.000 587.304 98.967 ;
 END
 PORT
  LAYER ME4 ;
  RECT 587.775 0.000 588.495 31.570 ;
 END
 PORT
  LAYER ME4 ;
  RECT 588.966 0.921 589.306 98.967 ;
 END
 PORT
  LAYER ME4 ;
  RECT 590.968 0.921 591.308 98.967 ;
 END
 PORT
  LAYER ME4 ;
  RECT 599.787 0.000 600.507 31.570 ;
 END
 PORT
  LAYER ME4 ;
  RECT 600.978 0.000 601.318 98.967 ;
 END
 PORT
  LAYER ME4 ;
  RECT 594.972 0.000 595.312 98.967 ;
 END
 PORT
  LAYER ME4 ;
  RECT 595.783 0.000 596.503 31.570 ;
 END
 PORT
  LAYER ME4 ;
  RECT 596.974 0.921 597.314 98.967 ;
 END
 PORT
  LAYER ME4 ;
  RECT 598.976 0.921 599.316 98.967 ;
 END
 PORT
  LAYER ME4 ;
  RECT 607.795 0.000 608.515 31.570 ;
 END
 PORT
  LAYER ME4 ;
  RECT 608.986 0.000 609.326 98.967 ;
 END
 PORT
  LAYER ME4 ;
  RECT 602.980 0.000 603.320 98.967 ;
 END
 PORT
  LAYER ME4 ;
  RECT 603.791 0.000 604.511 31.570 ;
 END
 PORT
  LAYER ME4 ;
  RECT 604.982 0.921 605.322 98.967 ;
 END
 PORT
  LAYER ME4 ;
  RECT 606.984 0.921 607.324 98.967 ;
 END
 PORT
  LAYER ME4 ;
  RECT 615.803 0.000 616.523 31.570 ;
 END
 PORT
  LAYER ME4 ;
  RECT 616.994 0.000 617.334 98.967 ;
 END
 PORT
  LAYER ME4 ;
  RECT 610.988 0.000 611.328 98.967 ;
 END
 PORT
  LAYER ME4 ;
  RECT 611.799 0.000 612.519 31.570 ;
 END
 PORT
  LAYER ME4 ;
  RECT 612.990 0.921 613.330 98.967 ;
 END
 PORT
  LAYER ME4 ;
  RECT 614.992 0.921 615.332 98.967 ;
 END
 PORT
  LAYER ME4 ;
  RECT 617.995 0.000 618.335 98.967 ;
 END
 PORT
  LAYER ME4 ;
  RECT 309.849 0.000 310.569 98.967 ;
 END
 PORT
  LAYER ME4 ;
  RECT 315.843 0.000 316.563 98.967 ;
 END
 PORT
  LAYER ME4 ;
  RECT 321.314 0.000 322.034 98.967 ;
 END
 PORT
  LAYER ME4 ;
  RECT 323.029 0.000 323.749 98.967 ;
 END
 PORT
  LAYER ME4 ;
  RECT 326.025 0.000 326.625 98.967 ;
 END
 PORT
  LAYER ME4 ;
  RECT 327.705 0.921 328.045 98.967 ;
 END
 PORT
  LAYER ME4 ;
  RECT 302.290 0.000 303.010 98.967 ;
 END
 PORT
  LAYER ME4 ;
  RECT 300.250 0.921 300.970 98.208 ;
 END
 PORT
  LAYER ME4 ;
  RECT 298.130 0.000 298.850 98.967 ;
 END
 PORT
  LAYER ME4 ;
  RECT 296.090 0.921 296.810 98.967 ;
 END
 PORT
  LAYER ME4 ;
  RECT 1.740 0.000 2.080 98.967 ;
 END
 PORT
  LAYER ME4 ;
  RECT 2.741 0.921 3.081 98.967 ;
 END
 PORT
  LAYER ME4 ;
  RECT 9.558 0.000 10.278 31.570 ;
 END
 PORT
  LAYER ME4 ;
  RECT 10.749 0.000 11.089 98.967 ;
 END
 PORT
  LAYER ME4 ;
  RECT 4.743 0.000 5.083 98.967 ;
 END
 PORT
  LAYER ME4 ;
  RECT 5.554 0.000 6.274 31.570 ;
 END
 PORT
  LAYER ME4 ;
  RECT 6.745 0.921 7.085 98.967 ;
 END
 PORT
  LAYER ME4 ;
  RECT 8.747 0.921 9.087 98.967 ;
 END
 PORT
  LAYER ME4 ;
  RECT 17.566 0.000 18.286 31.570 ;
 END
 PORT
  LAYER ME4 ;
  RECT 18.757 0.000 19.097 98.967 ;
 END
 PORT
  LAYER ME4 ;
  RECT 12.751 0.000 13.091 98.967 ;
 END
 PORT
  LAYER ME4 ;
  RECT 13.562 0.000 14.282 31.570 ;
 END
 PORT
  LAYER ME4 ;
  RECT 14.753 0.921 15.093 98.967 ;
 END
 PORT
  LAYER ME4 ;
  RECT 16.755 0.921 17.095 98.967 ;
 END
 PORT
  LAYER ME4 ;
  RECT 25.574 0.000 26.294 31.570 ;
 END
 PORT
  LAYER ME4 ;
  RECT 26.765 0.000 27.105 98.967 ;
 END
 PORT
  LAYER ME4 ;
  RECT 20.759 0.000 21.099 98.967 ;
 END
 PORT
  LAYER ME4 ;
  RECT 21.570 0.000 22.290 31.570 ;
 END
 PORT
  LAYER ME4 ;
  RECT 22.761 0.921 23.101 98.967 ;
 END
 PORT
  LAYER ME4 ;
  RECT 24.763 0.921 25.103 98.967 ;
 END
 PORT
  LAYER ME4 ;
  RECT 33.582 0.000 34.302 31.570 ;
 END
 PORT
  LAYER ME4 ;
  RECT 34.773 0.000 35.113 98.967 ;
 END
 PORT
  LAYER ME4 ;
  RECT 28.767 0.000 29.107 98.967 ;
 END
 PORT
  LAYER ME4 ;
  RECT 29.578 0.000 30.298 31.570 ;
 END
 PORT
  LAYER ME4 ;
  RECT 30.769 0.921 31.109 98.967 ;
 END
 PORT
  LAYER ME4 ;
  RECT 32.771 0.921 33.111 98.967 ;
 END
 PORT
  LAYER ME4 ;
  RECT 41.590 0.000 42.310 31.570 ;
 END
 PORT
  LAYER ME4 ;
  RECT 42.781 0.000 43.121 98.967 ;
 END
 PORT
  LAYER ME4 ;
  RECT 36.775 0.000 37.115 98.967 ;
 END
 PORT
  LAYER ME4 ;
  RECT 37.586 0.000 38.306 31.570 ;
 END
 PORT
  LAYER ME4 ;
  RECT 38.777 0.921 39.117 98.967 ;
 END
 PORT
  LAYER ME4 ;
  RECT 40.779 0.921 41.119 98.967 ;
 END
 PORT
  LAYER ME4 ;
  RECT 49.598 0.000 50.318 31.570 ;
 END
 PORT
  LAYER ME4 ;
  RECT 50.789 0.000 51.129 98.967 ;
 END
 PORT
  LAYER ME4 ;
  RECT 44.783 0.000 45.123 98.967 ;
 END
 PORT
  LAYER ME4 ;
  RECT 45.594 0.000 46.314 31.570 ;
 END
 PORT
  LAYER ME4 ;
  RECT 46.785 0.921 47.125 98.967 ;
 END
 PORT
  LAYER ME4 ;
  RECT 48.787 0.921 49.127 98.967 ;
 END
 PORT
  LAYER ME4 ;
  RECT 57.606 0.000 58.326 31.570 ;
 END
 PORT
  LAYER ME4 ;
  RECT 58.797 0.000 59.137 98.967 ;
 END
 PORT
  LAYER ME4 ;
  RECT 52.791 0.000 53.131 98.967 ;
 END
 PORT
  LAYER ME4 ;
  RECT 53.602 0.000 54.322 31.570 ;
 END
 PORT
  LAYER ME4 ;
  RECT 54.793 0.921 55.133 98.967 ;
 END
 PORT
  LAYER ME4 ;
  RECT 56.795 0.921 57.135 98.967 ;
 END
 PORT
  LAYER ME4 ;
  RECT 65.614 0.000 66.334 31.570 ;
 END
 PORT
  LAYER ME4 ;
  RECT 66.805 0.000 67.145 98.967 ;
 END
 PORT
  LAYER ME4 ;
  RECT 60.799 0.000 61.139 98.967 ;
 END
 PORT
  LAYER ME4 ;
  RECT 61.610 0.000 62.330 31.570 ;
 END
 PORT
  LAYER ME4 ;
  RECT 62.801 0.921 63.141 98.967 ;
 END
 PORT
  LAYER ME4 ;
  RECT 64.803 0.921 65.143 98.967 ;
 END
 PORT
  LAYER ME4 ;
  RECT 73.622 0.000 74.342 31.570 ;
 END
 PORT
  LAYER ME4 ;
  RECT 74.813 0.000 75.153 98.967 ;
 END
 PORT
  LAYER ME4 ;
  RECT 68.807 0.000 69.147 98.967 ;
 END
 PORT
  LAYER ME4 ;
  RECT 69.618 0.000 70.338 31.570 ;
 END
 PORT
  LAYER ME4 ;
  RECT 70.809 0.921 71.149 98.967 ;
 END
 PORT
  LAYER ME4 ;
  RECT 72.811 0.921 73.151 98.967 ;
 END
 PORT
  LAYER ME4 ;
  RECT 81.630 0.000 82.350 31.570 ;
 END
 PORT
  LAYER ME4 ;
  RECT 82.821 0.000 83.161 98.967 ;
 END
 PORT
  LAYER ME4 ;
  RECT 76.815 0.000 77.155 98.967 ;
 END
 PORT
  LAYER ME4 ;
  RECT 77.626 0.000 78.346 31.570 ;
 END
 PORT
  LAYER ME4 ;
  RECT 78.817 0.921 79.157 98.967 ;
 END
 PORT
  LAYER ME4 ;
  RECT 80.819 0.921 81.159 98.967 ;
 END
 PORT
  LAYER ME4 ;
  RECT 89.638 0.000 90.358 31.570 ;
 END
 PORT
  LAYER ME4 ;
  RECT 90.829 0.000 91.169 98.967 ;
 END
 PORT
  LAYER ME4 ;
  RECT 84.823 0.000 85.163 98.967 ;
 END
 PORT
  LAYER ME4 ;
  RECT 85.634 0.000 86.354 31.570 ;
 END
 PORT
  LAYER ME4 ;
  RECT 86.825 0.921 87.165 98.967 ;
 END
 PORT
  LAYER ME4 ;
  RECT 88.827 0.921 89.167 98.967 ;
 END
 PORT
  LAYER ME4 ;
  RECT 97.646 0.000 98.366 31.570 ;
 END
 PORT
  LAYER ME4 ;
  RECT 98.837 0.000 99.177 98.967 ;
 END
 PORT
  LAYER ME4 ;
  RECT 92.831 0.000 93.171 98.967 ;
 END
 PORT
  LAYER ME4 ;
  RECT 93.642 0.000 94.362 31.570 ;
 END
 PORT
  LAYER ME4 ;
  RECT 94.833 0.921 95.173 98.967 ;
 END
 PORT
  LAYER ME4 ;
  RECT 96.835 0.921 97.175 98.967 ;
 END
 PORT
  LAYER ME4 ;
  RECT 105.654 0.000 106.374 31.570 ;
 END
 PORT
  LAYER ME4 ;
  RECT 106.845 0.000 107.185 98.967 ;
 END
 PORT
  LAYER ME4 ;
  RECT 100.839 0.000 101.179 98.967 ;
 END
 PORT
  LAYER ME4 ;
  RECT 101.650 0.000 102.370 31.570 ;
 END
 PORT
  LAYER ME4 ;
  RECT 102.841 0.921 103.181 98.967 ;
 END
 PORT
  LAYER ME4 ;
  RECT 104.843 0.921 105.183 98.967 ;
 END
 PORT
  LAYER ME4 ;
  RECT 113.662 0.000 114.382 31.570 ;
 END
 PORT
  LAYER ME4 ;
  RECT 114.853 0.000 115.193 98.967 ;
 END
 PORT
  LAYER ME4 ;
  RECT 108.847 0.000 109.187 98.967 ;
 END
 PORT
  LAYER ME4 ;
  RECT 109.658 0.000 110.378 31.570 ;
 END
 PORT
  LAYER ME4 ;
  RECT 110.849 0.921 111.189 98.967 ;
 END
 PORT
  LAYER ME4 ;
  RECT 112.851 0.921 113.191 98.967 ;
 END
 PORT
  LAYER ME4 ;
  RECT 121.670 0.000 122.390 31.570 ;
 END
 PORT
  LAYER ME4 ;
  RECT 122.861 0.000 123.201 98.967 ;
 END
 PORT
  LAYER ME4 ;
  RECT 116.855 0.000 117.195 98.967 ;
 END
 PORT
  LAYER ME4 ;
  RECT 117.666 0.000 118.386 31.570 ;
 END
 PORT
  LAYER ME4 ;
  RECT 118.857 0.921 119.197 98.967 ;
 END
 PORT
  LAYER ME4 ;
  RECT 120.859 0.921 121.199 98.967 ;
 END
 PORT
  LAYER ME4 ;
  RECT 129.678 0.000 130.398 31.570 ;
 END
 PORT
  LAYER ME4 ;
  RECT 130.869 0.000 131.209 98.967 ;
 END
 PORT
  LAYER ME4 ;
  RECT 124.863 0.000 125.203 98.967 ;
 END
 PORT
  LAYER ME4 ;
  RECT 125.674 0.000 126.394 31.570 ;
 END
 PORT
  LAYER ME4 ;
  RECT 126.865 0.921 127.205 98.967 ;
 END
 PORT
  LAYER ME4 ;
  RECT 128.867 0.921 129.207 98.967 ;
 END
 PORT
  LAYER ME4 ;
  RECT 137.686 0.000 138.406 31.570 ;
 END
 PORT
  LAYER ME4 ;
  RECT 138.877 0.000 139.217 98.967 ;
 END
 PORT
  LAYER ME4 ;
  RECT 132.871 0.000 133.211 98.967 ;
 END
 PORT
  LAYER ME4 ;
  RECT 133.682 0.000 134.402 31.570 ;
 END
 PORT
  LAYER ME4 ;
  RECT 134.873 0.921 135.213 98.967 ;
 END
 PORT
  LAYER ME4 ;
  RECT 136.875 0.921 137.215 98.967 ;
 END
 PORT
  LAYER ME4 ;
  RECT 145.694 0.000 146.414 31.570 ;
 END
 PORT
  LAYER ME4 ;
  RECT 146.885 0.000 147.225 98.967 ;
 END
 PORT
  LAYER ME4 ;
  RECT 140.879 0.000 141.219 98.967 ;
 END
 PORT
  LAYER ME4 ;
  RECT 141.690 0.000 142.410 31.570 ;
 END
 PORT
  LAYER ME4 ;
  RECT 142.881 0.921 143.221 98.967 ;
 END
 PORT
  LAYER ME4 ;
  RECT 144.883 0.921 145.223 98.967 ;
 END
 PORT
  LAYER ME4 ;
  RECT 153.702 0.000 154.422 31.570 ;
 END
 PORT
  LAYER ME4 ;
  RECT 154.893 0.000 155.233 98.967 ;
 END
 PORT
  LAYER ME4 ;
  RECT 148.887 0.000 149.227 98.967 ;
 END
 PORT
  LAYER ME4 ;
  RECT 149.698 0.000 150.418 31.570 ;
 END
 PORT
  LAYER ME4 ;
  RECT 150.889 0.921 151.229 98.967 ;
 END
 PORT
  LAYER ME4 ;
  RECT 152.891 0.921 153.231 98.967 ;
 END
 PORT
  LAYER ME4 ;
  RECT 161.710 0.000 162.430 31.570 ;
 END
 PORT
  LAYER ME4 ;
  RECT 162.901 0.000 163.241 98.967 ;
 END
 PORT
  LAYER ME4 ;
  RECT 156.895 0.000 157.235 98.967 ;
 END
 PORT
  LAYER ME4 ;
  RECT 157.706 0.000 158.426 31.570 ;
 END
 PORT
  LAYER ME4 ;
  RECT 158.897 0.921 159.237 98.967 ;
 END
 PORT
  LAYER ME4 ;
  RECT 160.899 0.921 161.239 98.967 ;
 END
 PORT
  LAYER ME4 ;
  RECT 169.718 0.000 170.438 31.570 ;
 END
 PORT
  LAYER ME4 ;
  RECT 170.909 0.000 171.249 98.967 ;
 END
 PORT
  LAYER ME4 ;
  RECT 164.903 0.000 165.243 98.967 ;
 END
 PORT
  LAYER ME4 ;
  RECT 165.714 0.000 166.434 31.570 ;
 END
 PORT
  LAYER ME4 ;
  RECT 166.905 0.921 167.245 98.967 ;
 END
 PORT
  LAYER ME4 ;
  RECT 168.907 0.921 169.247 98.967 ;
 END
 PORT
  LAYER ME4 ;
  RECT 177.726 0.000 178.446 31.570 ;
 END
 PORT
  LAYER ME4 ;
  RECT 178.917 0.000 179.257 98.967 ;
 END
 PORT
  LAYER ME4 ;
  RECT 172.911 0.000 173.251 98.967 ;
 END
 PORT
  LAYER ME4 ;
  RECT 173.722 0.000 174.442 31.570 ;
 END
 PORT
  LAYER ME4 ;
  RECT 174.913 0.921 175.253 98.967 ;
 END
 PORT
  LAYER ME4 ;
  RECT 176.915 0.921 177.255 98.967 ;
 END
 PORT
  LAYER ME4 ;
  RECT 185.734 0.000 186.454 31.570 ;
 END
 PORT
  LAYER ME4 ;
  RECT 186.925 0.000 187.265 98.967 ;
 END
 PORT
  LAYER ME4 ;
  RECT 180.919 0.000 181.259 98.967 ;
 END
 PORT
  LAYER ME4 ;
  RECT 181.730 0.000 182.450 31.570 ;
 END
 PORT
  LAYER ME4 ;
  RECT 182.921 0.921 183.261 98.967 ;
 END
 PORT
  LAYER ME4 ;
  RECT 184.923 0.921 185.263 98.967 ;
 END
 PORT
  LAYER ME4 ;
  RECT 193.742 0.000 194.462 31.570 ;
 END
 PORT
  LAYER ME4 ;
  RECT 194.933 0.000 195.273 98.967 ;
 END
 PORT
  LAYER ME4 ;
  RECT 188.927 0.000 189.267 98.967 ;
 END
 PORT
  LAYER ME4 ;
  RECT 189.738 0.000 190.458 31.570 ;
 END
 PORT
  LAYER ME4 ;
  RECT 190.929 0.921 191.269 98.967 ;
 END
 PORT
  LAYER ME4 ;
  RECT 192.931 0.921 193.271 98.967 ;
 END
 PORT
  LAYER ME4 ;
  RECT 201.750 0.000 202.470 31.570 ;
 END
 PORT
  LAYER ME4 ;
  RECT 202.941 0.000 203.281 98.967 ;
 END
 PORT
  LAYER ME4 ;
  RECT 196.935 0.000 197.275 98.967 ;
 END
 PORT
  LAYER ME4 ;
  RECT 197.746 0.000 198.466 31.570 ;
 END
 PORT
  LAYER ME4 ;
  RECT 198.937 0.921 199.277 98.967 ;
 END
 PORT
  LAYER ME4 ;
  RECT 200.939 0.921 201.279 98.967 ;
 END
 PORT
  LAYER ME4 ;
  RECT 209.758 0.000 210.478 31.570 ;
 END
 PORT
  LAYER ME4 ;
  RECT 210.949 0.000 211.289 98.967 ;
 END
 PORT
  LAYER ME4 ;
  RECT 204.943 0.000 205.283 98.967 ;
 END
 PORT
  LAYER ME4 ;
  RECT 205.754 0.000 206.474 31.570 ;
 END
 PORT
  LAYER ME4 ;
  RECT 206.945 0.921 207.285 98.967 ;
 END
 PORT
  LAYER ME4 ;
  RECT 208.947 0.921 209.287 98.967 ;
 END
 PORT
  LAYER ME4 ;
  RECT 217.766 0.000 218.486 31.570 ;
 END
 PORT
  LAYER ME4 ;
  RECT 218.957 0.000 219.297 98.967 ;
 END
 PORT
  LAYER ME4 ;
  RECT 212.951 0.000 213.291 98.967 ;
 END
 PORT
  LAYER ME4 ;
  RECT 213.762 0.000 214.482 31.570 ;
 END
 PORT
  LAYER ME4 ;
  RECT 214.953 0.921 215.293 98.967 ;
 END
 PORT
  LAYER ME4 ;
  RECT 216.955 0.921 217.295 98.967 ;
 END
 PORT
  LAYER ME4 ;
  RECT 225.774 0.000 226.494 31.570 ;
 END
 PORT
  LAYER ME4 ;
  RECT 226.965 0.000 227.305 98.967 ;
 END
 PORT
  LAYER ME4 ;
  RECT 220.959 0.000 221.299 98.967 ;
 END
 PORT
  LAYER ME4 ;
  RECT 221.770 0.000 222.490 31.570 ;
 END
 PORT
  LAYER ME4 ;
  RECT 222.961 0.921 223.301 98.967 ;
 END
 PORT
  LAYER ME4 ;
  RECT 224.963 0.921 225.303 98.967 ;
 END
 PORT
  LAYER ME4 ;
  RECT 233.782 0.000 234.502 31.570 ;
 END
 PORT
  LAYER ME4 ;
  RECT 234.973 0.000 235.313 98.967 ;
 END
 PORT
  LAYER ME4 ;
  RECT 228.967 0.000 229.307 98.967 ;
 END
 PORT
  LAYER ME4 ;
  RECT 229.778 0.000 230.498 31.570 ;
 END
 PORT
  LAYER ME4 ;
  RECT 230.969 0.921 231.309 98.967 ;
 END
 PORT
  LAYER ME4 ;
  RECT 232.971 0.921 233.311 98.967 ;
 END
 PORT
  LAYER ME4 ;
  RECT 241.790 0.000 242.510 31.570 ;
 END
 PORT
  LAYER ME4 ;
  RECT 242.981 0.000 243.321 98.967 ;
 END
 PORT
  LAYER ME4 ;
  RECT 236.975 0.000 237.315 98.967 ;
 END
 PORT
  LAYER ME4 ;
  RECT 237.786 0.000 238.506 31.570 ;
 END
 PORT
  LAYER ME4 ;
  RECT 238.977 0.921 239.317 98.967 ;
 END
 PORT
  LAYER ME4 ;
  RECT 240.979 0.921 241.319 98.967 ;
 END
 PORT
  LAYER ME4 ;
  RECT 249.798 0.000 250.518 31.570 ;
 END
 PORT
  LAYER ME4 ;
  RECT 250.989 0.000 251.329 98.967 ;
 END
 PORT
  LAYER ME4 ;
  RECT 244.983 0.000 245.323 98.967 ;
 END
 PORT
  LAYER ME4 ;
  RECT 245.794 0.000 246.514 31.570 ;
 END
 PORT
  LAYER ME4 ;
  RECT 246.985 0.921 247.325 98.967 ;
 END
 PORT
  LAYER ME4 ;
  RECT 248.987 0.921 249.327 98.967 ;
 END
 PORT
  LAYER ME4 ;
  RECT 257.806 0.000 258.526 31.570 ;
 END
 PORT
  LAYER ME4 ;
  RECT 258.997 0.000 259.337 98.967 ;
 END
 PORT
  LAYER ME4 ;
  RECT 252.991 0.000 253.331 98.967 ;
 END
 PORT
  LAYER ME4 ;
  RECT 253.802 0.000 254.522 31.570 ;
 END
 PORT
  LAYER ME4 ;
  RECT 254.993 0.921 255.333 98.967 ;
 END
 PORT
  LAYER ME4 ;
  RECT 256.995 0.921 257.335 98.967 ;
 END
 PORT
  LAYER ME4 ;
  RECT 265.814 0.000 266.534 31.570 ;
 END
 PORT
  LAYER ME4 ;
  RECT 267.005 0.000 267.345 98.967 ;
 END
 PORT
  LAYER ME4 ;
  RECT 260.999 0.000 261.339 98.967 ;
 END
 PORT
  LAYER ME4 ;
  RECT 261.810 0.000 262.530 31.570 ;
 END
 PORT
  LAYER ME4 ;
  RECT 263.001 0.921 263.341 98.967 ;
 END
 PORT
  LAYER ME4 ;
  RECT 265.003 0.921 265.343 98.967 ;
 END
 PORT
  LAYER ME4 ;
  RECT 273.822 0.000 274.542 31.570 ;
 END
 PORT
  LAYER ME4 ;
  RECT 275.013 0.000 275.353 98.967 ;
 END
 PORT
  LAYER ME4 ;
  RECT 269.007 0.000 269.347 98.967 ;
 END
 PORT
  LAYER ME4 ;
  RECT 269.818 0.000 270.538 31.570 ;
 END
 PORT
  LAYER ME4 ;
  RECT 271.009 0.921 271.349 98.967 ;
 END
 PORT
  LAYER ME4 ;
  RECT 273.011 0.921 273.351 98.967 ;
 END
 PORT
  LAYER ME4 ;
  RECT 281.830 0.000 282.550 31.570 ;
 END
 PORT
  LAYER ME4 ;
  RECT 283.021 0.000 283.361 98.967 ;
 END
 PORT
  LAYER ME4 ;
  RECT 277.015 0.000 277.355 98.967 ;
 END
 PORT
  LAYER ME4 ;
  RECT 277.826 0.000 278.546 31.570 ;
 END
 PORT
  LAYER ME4 ;
  RECT 279.017 0.921 279.357 98.967 ;
 END
 PORT
  LAYER ME4 ;
  RECT 281.019 0.921 281.359 98.967 ;
 END
 PORT
  LAYER ME4 ;
  RECT 289.838 0.000 290.558 31.570 ;
 END
 PORT
  LAYER ME4 ;
  RECT 291.029 0.000 291.369 98.967 ;
 END
 PORT
  LAYER ME4 ;
  RECT 285.023 0.000 285.363 98.967 ;
 END
 PORT
  LAYER ME4 ;
  RECT 285.834 0.000 286.554 31.570 ;
 END
 PORT
  LAYER ME4 ;
  RECT 287.025 0.921 287.365 98.967 ;
 END
 PORT
  LAYER ME4 ;
  RECT 289.027 0.921 289.367 98.967 ;
 END
 PORT
  LAYER ME4 ;
  RECT 293.970 0.000 294.690 98.967 ;
 END
 PORT
  LAYER ME4 ;
  RECT 292.030 0.000 292.370 98.967 ;
 END
END GND
PIN DI35
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 288.886 0.000 289.166 0.720 ;
  LAYER ME3 ;
  RECT 288.886 0.000 289.166 0.720 ;
  LAYER ME2 ;
  RECT 288.886 0.000 289.166 0.720 ;
  LAYER ME1 ;
  RECT 288.886 0.000 289.166 0.720 ;
 END
 ANTENNAPARTIALMETALAREA                  0.805 LAYER ME1 ;
 ANTENNAGATEAREA                          0.072 LAYER ME1 ;
 ANTENNAGATEAREA                          0.072 LAYER ME2 ;
 ANTENNAGATEAREA                          0.072 LAYER ME3 ;
 ANTENNAGATEAREA                          0.072 LAYER ME4 ;
 ANTENNADIFFAREA                          0.218 LAYER ME1 ;
 ANTENNADIFFAREA                          0.218 LAYER ME2 ;
 ANTENNADIFFAREA                          0.218 LAYER ME3 ;
 ANTENNADIFFAREA                          0.218 LAYER ME4 ;
 ANTENNAMAXAREACAR                       13.984 LAYER ME1 ;
 ANTENNAMAXAREACAR                       16.784 LAYER ME2 ;
 ANTENNAMAXAREACAR                       19.584 LAYER ME3 ;
 ANTENNAMAXAREACAR                       22.384 LAYER ME4 ;
END DI35
PIN DO35
  DIRECTION OUTPUT ;
 PORT
  LAYER ME4 ;
  RECT 286.908 0.000 287.188 0.720 ;
  LAYER ME3 ;
  RECT 286.908 0.000 287.188 0.720 ;
  LAYER ME2 ;
  RECT 286.908 0.000 287.188 0.720 ;
  LAYER ME1 ;
  RECT 286.908 0.000 287.188 0.720 ;
 END
 ANTENNAPARTIALMETALAREA                  2.030 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME3 ;
 ANTENNADIFFAREA                          1.293 LAYER ME4 ;
END DO35
PIN DI34
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 280.878 0.000 281.158 0.720 ;
  LAYER ME3 ;
  RECT 280.878 0.000 281.158 0.720 ;
  LAYER ME2 ;
  RECT 280.878 0.000 281.158 0.720 ;
  LAYER ME1 ;
  RECT 280.878 0.000 281.158 0.720 ;
 END
 ANTENNAPARTIALMETALAREA                  0.805 LAYER ME1 ;
 ANTENNAGATEAREA                          0.072 LAYER ME1 ;
 ANTENNAGATEAREA                          0.072 LAYER ME2 ;
 ANTENNAGATEAREA                          0.072 LAYER ME3 ;
 ANTENNAGATEAREA                          0.072 LAYER ME4 ;
 ANTENNADIFFAREA                          0.218 LAYER ME1 ;
 ANTENNADIFFAREA                          0.218 LAYER ME2 ;
 ANTENNADIFFAREA                          0.218 LAYER ME3 ;
 ANTENNADIFFAREA                          0.218 LAYER ME4 ;
 ANTENNAMAXAREACAR                       13.984 LAYER ME1 ;
 ANTENNAMAXAREACAR                       16.784 LAYER ME2 ;
 ANTENNAMAXAREACAR                       19.584 LAYER ME3 ;
 ANTENNAMAXAREACAR                       22.384 LAYER ME4 ;
END DI34
PIN DO34
  DIRECTION OUTPUT ;
 PORT
  LAYER ME4 ;
  RECT 278.900 0.000 279.180 0.720 ;
  LAYER ME3 ;
  RECT 278.900 0.000 279.180 0.720 ;
  LAYER ME2 ;
  RECT 278.900 0.000 279.180 0.720 ;
  LAYER ME1 ;
  RECT 278.900 0.000 279.180 0.720 ;
 END
 ANTENNAPARTIALMETALAREA                  2.030 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME3 ;
 ANTENNADIFFAREA                          1.293 LAYER ME4 ;
END DO34
PIN DI33
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 272.870 0.000 273.150 0.720 ;
  LAYER ME3 ;
  RECT 272.870 0.000 273.150 0.720 ;
  LAYER ME2 ;
  RECT 272.870 0.000 273.150 0.720 ;
  LAYER ME1 ;
  RECT 272.870 0.000 273.150 0.720 ;
 END
 ANTENNAPARTIALMETALAREA                  0.805 LAYER ME1 ;
 ANTENNAGATEAREA                          0.072 LAYER ME1 ;
 ANTENNAGATEAREA                          0.072 LAYER ME2 ;
 ANTENNAGATEAREA                          0.072 LAYER ME3 ;
 ANTENNAGATEAREA                          0.072 LAYER ME4 ;
 ANTENNADIFFAREA                          0.218 LAYER ME1 ;
 ANTENNADIFFAREA                          0.218 LAYER ME2 ;
 ANTENNADIFFAREA                          0.218 LAYER ME3 ;
 ANTENNADIFFAREA                          0.218 LAYER ME4 ;
 ANTENNAMAXAREACAR                       13.984 LAYER ME1 ;
 ANTENNAMAXAREACAR                       16.784 LAYER ME2 ;
 ANTENNAMAXAREACAR                       19.584 LAYER ME3 ;
 ANTENNAMAXAREACAR                       22.384 LAYER ME4 ;
END DI33
PIN DO33
  DIRECTION OUTPUT ;
 PORT
  LAYER ME4 ;
  RECT 270.892 0.000 271.172 0.720 ;
  LAYER ME3 ;
  RECT 270.892 0.000 271.172 0.720 ;
  LAYER ME2 ;
  RECT 270.892 0.000 271.172 0.720 ;
  LAYER ME1 ;
  RECT 270.892 0.000 271.172 0.720 ;
 END
 ANTENNAPARTIALMETALAREA                  2.030 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME3 ;
 ANTENNADIFFAREA                          1.293 LAYER ME4 ;
END DO33
PIN DI32
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 264.862 0.000 265.142 0.720 ;
  LAYER ME3 ;
  RECT 264.862 0.000 265.142 0.720 ;
  LAYER ME2 ;
  RECT 264.862 0.000 265.142 0.720 ;
  LAYER ME1 ;
  RECT 264.862 0.000 265.142 0.720 ;
 END
 ANTENNAPARTIALMETALAREA                  0.805 LAYER ME1 ;
 ANTENNAGATEAREA                          0.072 LAYER ME1 ;
 ANTENNAGATEAREA                          0.072 LAYER ME2 ;
 ANTENNAGATEAREA                          0.072 LAYER ME3 ;
 ANTENNAGATEAREA                          0.072 LAYER ME4 ;
 ANTENNADIFFAREA                          0.218 LAYER ME1 ;
 ANTENNADIFFAREA                          0.218 LAYER ME2 ;
 ANTENNADIFFAREA                          0.218 LAYER ME3 ;
 ANTENNADIFFAREA                          0.218 LAYER ME4 ;
 ANTENNAMAXAREACAR                       13.984 LAYER ME1 ;
 ANTENNAMAXAREACAR                       16.784 LAYER ME2 ;
 ANTENNAMAXAREACAR                       19.584 LAYER ME3 ;
 ANTENNAMAXAREACAR                       22.384 LAYER ME4 ;
END DI32
PIN DO32
  DIRECTION OUTPUT ;
 PORT
  LAYER ME4 ;
  RECT 262.884 0.000 263.164 0.720 ;
  LAYER ME3 ;
  RECT 262.884 0.000 263.164 0.720 ;
  LAYER ME2 ;
  RECT 262.884 0.000 263.164 0.720 ;
  LAYER ME1 ;
  RECT 262.884 0.000 263.164 0.720 ;
 END
 ANTENNAPARTIALMETALAREA                  2.030 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME3 ;
 ANTENNADIFFAREA                          1.293 LAYER ME4 ;
END DO32
PIN DI31
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 256.854 0.000 257.134 0.720 ;
  LAYER ME3 ;
  RECT 256.854 0.000 257.134 0.720 ;
  LAYER ME2 ;
  RECT 256.854 0.000 257.134 0.720 ;
  LAYER ME1 ;
  RECT 256.854 0.000 257.134 0.720 ;
 END
 ANTENNAPARTIALMETALAREA                  0.805 LAYER ME1 ;
 ANTENNAGATEAREA                          0.072 LAYER ME1 ;
 ANTENNAGATEAREA                          0.072 LAYER ME2 ;
 ANTENNAGATEAREA                          0.072 LAYER ME3 ;
 ANTENNAGATEAREA                          0.072 LAYER ME4 ;
 ANTENNADIFFAREA                          0.218 LAYER ME1 ;
 ANTENNADIFFAREA                          0.218 LAYER ME2 ;
 ANTENNADIFFAREA                          0.218 LAYER ME3 ;
 ANTENNADIFFAREA                          0.218 LAYER ME4 ;
 ANTENNAMAXAREACAR                       13.984 LAYER ME1 ;
 ANTENNAMAXAREACAR                       16.784 LAYER ME2 ;
 ANTENNAMAXAREACAR                       19.584 LAYER ME3 ;
 ANTENNAMAXAREACAR                       22.384 LAYER ME4 ;
END DI31
PIN DO31
  DIRECTION OUTPUT ;
 PORT
  LAYER ME4 ;
  RECT 254.876 0.000 255.156 0.720 ;
  LAYER ME3 ;
  RECT 254.876 0.000 255.156 0.720 ;
  LAYER ME2 ;
  RECT 254.876 0.000 255.156 0.720 ;
  LAYER ME1 ;
  RECT 254.876 0.000 255.156 0.720 ;
 END
 ANTENNAPARTIALMETALAREA                  2.030 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME3 ;
 ANTENNADIFFAREA                          1.293 LAYER ME4 ;
END DO31
PIN DI30
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 248.846 0.000 249.126 0.720 ;
  LAYER ME3 ;
  RECT 248.846 0.000 249.126 0.720 ;
  LAYER ME2 ;
  RECT 248.846 0.000 249.126 0.720 ;
  LAYER ME1 ;
  RECT 248.846 0.000 249.126 0.720 ;
 END
 ANTENNAPARTIALMETALAREA                  0.805 LAYER ME1 ;
 ANTENNAGATEAREA                          0.072 LAYER ME1 ;
 ANTENNAGATEAREA                          0.072 LAYER ME2 ;
 ANTENNAGATEAREA                          0.072 LAYER ME3 ;
 ANTENNAGATEAREA                          0.072 LAYER ME4 ;
 ANTENNADIFFAREA                          0.218 LAYER ME1 ;
 ANTENNADIFFAREA                          0.218 LAYER ME2 ;
 ANTENNADIFFAREA                          0.218 LAYER ME3 ;
 ANTENNADIFFAREA                          0.218 LAYER ME4 ;
 ANTENNAMAXAREACAR                       13.984 LAYER ME1 ;
 ANTENNAMAXAREACAR                       16.784 LAYER ME2 ;
 ANTENNAMAXAREACAR                       19.584 LAYER ME3 ;
 ANTENNAMAXAREACAR                       22.384 LAYER ME4 ;
END DI30
PIN DO30
  DIRECTION OUTPUT ;
 PORT
  LAYER ME4 ;
  RECT 246.868 0.000 247.148 0.720 ;
  LAYER ME3 ;
  RECT 246.868 0.000 247.148 0.720 ;
  LAYER ME2 ;
  RECT 246.868 0.000 247.148 0.720 ;
  LAYER ME1 ;
  RECT 246.868 0.000 247.148 0.720 ;
 END
 ANTENNAPARTIALMETALAREA                  2.030 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME3 ;
 ANTENNADIFFAREA                          1.293 LAYER ME4 ;
END DO30
PIN DI29
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 240.838 0.000 241.118 0.720 ;
  LAYER ME3 ;
  RECT 240.838 0.000 241.118 0.720 ;
  LAYER ME2 ;
  RECT 240.838 0.000 241.118 0.720 ;
  LAYER ME1 ;
  RECT 240.838 0.000 241.118 0.720 ;
 END
 ANTENNAPARTIALMETALAREA                  0.805 LAYER ME1 ;
 ANTENNAGATEAREA                          0.072 LAYER ME1 ;
 ANTENNAGATEAREA                          0.072 LAYER ME2 ;
 ANTENNAGATEAREA                          0.072 LAYER ME3 ;
 ANTENNAGATEAREA                          0.072 LAYER ME4 ;
 ANTENNADIFFAREA                          0.218 LAYER ME1 ;
 ANTENNADIFFAREA                          0.218 LAYER ME2 ;
 ANTENNADIFFAREA                          0.218 LAYER ME3 ;
 ANTENNADIFFAREA                          0.218 LAYER ME4 ;
 ANTENNAMAXAREACAR                       13.984 LAYER ME1 ;
 ANTENNAMAXAREACAR                       16.784 LAYER ME2 ;
 ANTENNAMAXAREACAR                       19.584 LAYER ME3 ;
 ANTENNAMAXAREACAR                       22.384 LAYER ME4 ;
END DI29
PIN DO29
  DIRECTION OUTPUT ;
 PORT
  LAYER ME4 ;
  RECT 238.860 0.000 239.140 0.720 ;
  LAYER ME3 ;
  RECT 238.860 0.000 239.140 0.720 ;
  LAYER ME2 ;
  RECT 238.860 0.000 239.140 0.720 ;
  LAYER ME1 ;
  RECT 238.860 0.000 239.140 0.720 ;
 END
 ANTENNAPARTIALMETALAREA                  2.030 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME3 ;
 ANTENNADIFFAREA                          1.293 LAYER ME4 ;
END DO29
PIN DI28
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 232.830 0.000 233.110 0.720 ;
  LAYER ME3 ;
  RECT 232.830 0.000 233.110 0.720 ;
  LAYER ME2 ;
  RECT 232.830 0.000 233.110 0.720 ;
  LAYER ME1 ;
  RECT 232.830 0.000 233.110 0.720 ;
 END
 ANTENNAPARTIALMETALAREA                  0.805 LAYER ME1 ;
 ANTENNAGATEAREA                          0.072 LAYER ME1 ;
 ANTENNAGATEAREA                          0.072 LAYER ME2 ;
 ANTENNAGATEAREA                          0.072 LAYER ME3 ;
 ANTENNAGATEAREA                          0.072 LAYER ME4 ;
 ANTENNADIFFAREA                          0.218 LAYER ME1 ;
 ANTENNADIFFAREA                          0.218 LAYER ME2 ;
 ANTENNADIFFAREA                          0.218 LAYER ME3 ;
 ANTENNADIFFAREA                          0.218 LAYER ME4 ;
 ANTENNAMAXAREACAR                       13.984 LAYER ME1 ;
 ANTENNAMAXAREACAR                       16.784 LAYER ME2 ;
 ANTENNAMAXAREACAR                       19.584 LAYER ME3 ;
 ANTENNAMAXAREACAR                       22.384 LAYER ME4 ;
END DI28
PIN DO28
  DIRECTION OUTPUT ;
 PORT
  LAYER ME4 ;
  RECT 230.852 0.000 231.132 0.720 ;
  LAYER ME3 ;
  RECT 230.852 0.000 231.132 0.720 ;
  LAYER ME2 ;
  RECT 230.852 0.000 231.132 0.720 ;
  LAYER ME1 ;
  RECT 230.852 0.000 231.132 0.720 ;
 END
 ANTENNAPARTIALMETALAREA                  2.030 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME3 ;
 ANTENNADIFFAREA                          1.293 LAYER ME4 ;
END DO28
PIN DI27
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 224.822 0.000 225.102 0.720 ;
  LAYER ME3 ;
  RECT 224.822 0.000 225.102 0.720 ;
  LAYER ME2 ;
  RECT 224.822 0.000 225.102 0.720 ;
  LAYER ME1 ;
  RECT 224.822 0.000 225.102 0.720 ;
 END
 ANTENNAPARTIALMETALAREA                  0.522 LAYER ME1 ;
 ANTENNAGATEAREA                          0.072 LAYER ME1 ;
 ANTENNAGATEAREA                          0.072 LAYER ME2 ;
 ANTENNAGATEAREA                          0.072 LAYER ME3 ;
 ANTENNAGATEAREA                          0.072 LAYER ME4 ;
 ANTENNADIFFAREA                          0.218 LAYER ME1 ;
 ANTENNADIFFAREA                          0.218 LAYER ME2 ;
 ANTENNADIFFAREA                          0.218 LAYER ME3 ;
 ANTENNADIFFAREA                          0.218 LAYER ME4 ;
 ANTENNAMAXAREACAR                       10.048 LAYER ME1 ;
 ANTENNAMAXAREACAR                       12.848 LAYER ME2 ;
 ANTENNAMAXAREACAR                       15.648 LAYER ME3 ;
 ANTENNAMAXAREACAR                       18.448 LAYER ME4 ;
END DI27
PIN DO27
  DIRECTION OUTPUT ;
 PORT
  LAYER ME4 ;
  RECT 222.764 0.000 223.044 0.720 ;
  LAYER ME3 ;
  RECT 222.764 0.000 223.044 0.720 ;
  LAYER ME2 ;
  RECT 222.764 0.000 223.044 0.720 ;
  LAYER ME1 ;
  RECT 222.764 0.000 223.044 0.720 ;
 END
 ANTENNAPARTIALMETALAREA                  2.030 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME3 ;
 ANTENNADIFFAREA                          1.293 LAYER ME4 ;
END DO27
PIN WEB3
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 223.244 0.000 223.524 0.720 ;
  LAYER ME3 ;
  RECT 223.244 0.000 223.524 0.720 ;
  LAYER ME2 ;
  RECT 223.244 0.000 223.524 0.720 ;
  LAYER ME1 ;
  RECT 223.244 0.000 223.524 0.720 ;
 END
 ANTENNAPARTIALMETALAREA                  0.436 LAYER ME2 ;
 ANTENNAGATEAREA                          0.288 LAYER ME2 ;
 ANTENNAGATEAREA                          0.288 LAYER ME3 ;
 ANTENNAGATEAREA                          0.288 LAYER ME4 ;
 ANTENNADIFFAREA                          0.218 LAYER ME2 ;
 ANTENNADIFFAREA                          0.218 LAYER ME3 ;
 ANTENNADIFFAREA                          0.218 LAYER ME4 ;
 ANTENNAMAXAREACAR                        4.602 LAYER ME2 ;
 ANTENNAMAXAREACAR                        5.302 LAYER ME3 ;
 ANTENNAMAXAREACAR                        6.002 LAYER ME4 ;
END WEB3
PIN DI26
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 216.814 0.000 217.094 0.720 ;
  LAYER ME3 ;
  RECT 216.814 0.000 217.094 0.720 ;
  LAYER ME2 ;
  RECT 216.814 0.000 217.094 0.720 ;
  LAYER ME1 ;
  RECT 216.814 0.000 217.094 0.720 ;
 END
 ANTENNAPARTIALMETALAREA                  0.805 LAYER ME1 ;
 ANTENNAGATEAREA                          0.072 LAYER ME1 ;
 ANTENNAGATEAREA                          0.072 LAYER ME2 ;
 ANTENNAGATEAREA                          0.072 LAYER ME3 ;
 ANTENNAGATEAREA                          0.072 LAYER ME4 ;
 ANTENNADIFFAREA                          0.218 LAYER ME1 ;
 ANTENNADIFFAREA                          0.218 LAYER ME2 ;
 ANTENNADIFFAREA                          0.218 LAYER ME3 ;
 ANTENNADIFFAREA                          0.218 LAYER ME4 ;
 ANTENNAMAXAREACAR                       13.984 LAYER ME1 ;
 ANTENNAMAXAREACAR                       16.784 LAYER ME2 ;
 ANTENNAMAXAREACAR                       19.584 LAYER ME3 ;
 ANTENNAMAXAREACAR                       22.384 LAYER ME4 ;
END DI26
PIN DO26
  DIRECTION OUTPUT ;
 PORT
  LAYER ME4 ;
  RECT 214.836 0.000 215.116 0.720 ;
  LAYER ME3 ;
  RECT 214.836 0.000 215.116 0.720 ;
  LAYER ME2 ;
  RECT 214.836 0.000 215.116 0.720 ;
  LAYER ME1 ;
  RECT 214.836 0.000 215.116 0.720 ;
 END
 ANTENNAPARTIALMETALAREA                  2.030 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME3 ;
 ANTENNADIFFAREA                          1.293 LAYER ME4 ;
END DO26
PIN DI25
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 208.806 0.000 209.086 0.720 ;
  LAYER ME3 ;
  RECT 208.806 0.000 209.086 0.720 ;
  LAYER ME2 ;
  RECT 208.806 0.000 209.086 0.720 ;
  LAYER ME1 ;
  RECT 208.806 0.000 209.086 0.720 ;
 END
 ANTENNAPARTIALMETALAREA                  0.805 LAYER ME1 ;
 ANTENNAGATEAREA                          0.072 LAYER ME1 ;
 ANTENNAGATEAREA                          0.072 LAYER ME2 ;
 ANTENNAGATEAREA                          0.072 LAYER ME3 ;
 ANTENNAGATEAREA                          0.072 LAYER ME4 ;
 ANTENNADIFFAREA                          0.218 LAYER ME1 ;
 ANTENNADIFFAREA                          0.218 LAYER ME2 ;
 ANTENNADIFFAREA                          0.218 LAYER ME3 ;
 ANTENNADIFFAREA                          0.218 LAYER ME4 ;
 ANTENNAMAXAREACAR                       13.984 LAYER ME1 ;
 ANTENNAMAXAREACAR                       16.784 LAYER ME2 ;
 ANTENNAMAXAREACAR                       19.584 LAYER ME3 ;
 ANTENNAMAXAREACAR                       22.384 LAYER ME4 ;
END DI25
PIN DO25
  DIRECTION OUTPUT ;
 PORT
  LAYER ME4 ;
  RECT 206.828 0.000 207.108 0.720 ;
  LAYER ME3 ;
  RECT 206.828 0.000 207.108 0.720 ;
  LAYER ME2 ;
  RECT 206.828 0.000 207.108 0.720 ;
  LAYER ME1 ;
  RECT 206.828 0.000 207.108 0.720 ;
 END
 ANTENNAPARTIALMETALAREA                  2.030 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME3 ;
 ANTENNADIFFAREA                          1.293 LAYER ME4 ;
END DO25
PIN DI24
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 200.798 0.000 201.078 0.720 ;
  LAYER ME3 ;
  RECT 200.798 0.000 201.078 0.720 ;
  LAYER ME2 ;
  RECT 200.798 0.000 201.078 0.720 ;
  LAYER ME1 ;
  RECT 200.798 0.000 201.078 0.720 ;
 END
 ANTENNAPARTIALMETALAREA                  0.805 LAYER ME1 ;
 ANTENNAGATEAREA                          0.072 LAYER ME1 ;
 ANTENNAGATEAREA                          0.072 LAYER ME2 ;
 ANTENNAGATEAREA                          0.072 LAYER ME3 ;
 ANTENNAGATEAREA                          0.072 LAYER ME4 ;
 ANTENNADIFFAREA                          0.218 LAYER ME1 ;
 ANTENNADIFFAREA                          0.218 LAYER ME2 ;
 ANTENNADIFFAREA                          0.218 LAYER ME3 ;
 ANTENNADIFFAREA                          0.218 LAYER ME4 ;
 ANTENNAMAXAREACAR                       13.984 LAYER ME1 ;
 ANTENNAMAXAREACAR                       16.784 LAYER ME2 ;
 ANTENNAMAXAREACAR                       19.584 LAYER ME3 ;
 ANTENNAMAXAREACAR                       22.384 LAYER ME4 ;
END DI24
PIN DO24
  DIRECTION OUTPUT ;
 PORT
  LAYER ME4 ;
  RECT 198.820 0.000 199.100 0.720 ;
  LAYER ME3 ;
  RECT 198.820 0.000 199.100 0.720 ;
  LAYER ME2 ;
  RECT 198.820 0.000 199.100 0.720 ;
  LAYER ME1 ;
  RECT 198.820 0.000 199.100 0.720 ;
 END
 ANTENNAPARTIALMETALAREA                  2.030 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME3 ;
 ANTENNADIFFAREA                          1.293 LAYER ME4 ;
END DO24
PIN DI23
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 192.790 0.000 193.070 0.720 ;
  LAYER ME3 ;
  RECT 192.790 0.000 193.070 0.720 ;
  LAYER ME2 ;
  RECT 192.790 0.000 193.070 0.720 ;
  LAYER ME1 ;
  RECT 192.790 0.000 193.070 0.720 ;
 END
 ANTENNAPARTIALMETALAREA                  0.805 LAYER ME1 ;
 ANTENNAGATEAREA                          0.072 LAYER ME1 ;
 ANTENNAGATEAREA                          0.072 LAYER ME2 ;
 ANTENNAGATEAREA                          0.072 LAYER ME3 ;
 ANTENNAGATEAREA                          0.072 LAYER ME4 ;
 ANTENNADIFFAREA                          0.218 LAYER ME1 ;
 ANTENNADIFFAREA                          0.218 LAYER ME2 ;
 ANTENNADIFFAREA                          0.218 LAYER ME3 ;
 ANTENNADIFFAREA                          0.218 LAYER ME4 ;
 ANTENNAMAXAREACAR                       13.984 LAYER ME1 ;
 ANTENNAMAXAREACAR                       16.784 LAYER ME2 ;
 ANTENNAMAXAREACAR                       19.584 LAYER ME3 ;
 ANTENNAMAXAREACAR                       22.384 LAYER ME4 ;
END DI23
PIN DO23
  DIRECTION OUTPUT ;
 PORT
  LAYER ME4 ;
  RECT 190.812 0.000 191.092 0.720 ;
  LAYER ME3 ;
  RECT 190.812 0.000 191.092 0.720 ;
  LAYER ME2 ;
  RECT 190.812 0.000 191.092 0.720 ;
  LAYER ME1 ;
  RECT 190.812 0.000 191.092 0.720 ;
 END
 ANTENNAPARTIALMETALAREA                  2.030 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME3 ;
 ANTENNADIFFAREA                          1.293 LAYER ME4 ;
END DO23
PIN DI22
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 184.782 0.000 185.062 0.720 ;
  LAYER ME3 ;
  RECT 184.782 0.000 185.062 0.720 ;
  LAYER ME2 ;
  RECT 184.782 0.000 185.062 0.720 ;
  LAYER ME1 ;
  RECT 184.782 0.000 185.062 0.720 ;
 END
 ANTENNAPARTIALMETALAREA                  0.805 LAYER ME1 ;
 ANTENNAGATEAREA                          0.072 LAYER ME1 ;
 ANTENNAGATEAREA                          0.072 LAYER ME2 ;
 ANTENNAGATEAREA                          0.072 LAYER ME3 ;
 ANTENNAGATEAREA                          0.072 LAYER ME4 ;
 ANTENNADIFFAREA                          0.218 LAYER ME1 ;
 ANTENNADIFFAREA                          0.218 LAYER ME2 ;
 ANTENNADIFFAREA                          0.218 LAYER ME3 ;
 ANTENNADIFFAREA                          0.218 LAYER ME4 ;
 ANTENNAMAXAREACAR                       13.984 LAYER ME1 ;
 ANTENNAMAXAREACAR                       16.784 LAYER ME2 ;
 ANTENNAMAXAREACAR                       19.584 LAYER ME3 ;
 ANTENNAMAXAREACAR                       22.384 LAYER ME4 ;
END DI22
PIN DO22
  DIRECTION OUTPUT ;
 PORT
  LAYER ME4 ;
  RECT 182.804 0.000 183.084 0.720 ;
  LAYER ME3 ;
  RECT 182.804 0.000 183.084 0.720 ;
  LAYER ME2 ;
  RECT 182.804 0.000 183.084 0.720 ;
  LAYER ME1 ;
  RECT 182.804 0.000 183.084 0.720 ;
 END
 ANTENNAPARTIALMETALAREA                  2.030 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME3 ;
 ANTENNADIFFAREA                          1.293 LAYER ME4 ;
END DO22
PIN DI21
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 176.774 0.000 177.054 0.720 ;
  LAYER ME3 ;
  RECT 176.774 0.000 177.054 0.720 ;
  LAYER ME2 ;
  RECT 176.774 0.000 177.054 0.720 ;
  LAYER ME1 ;
  RECT 176.774 0.000 177.054 0.720 ;
 END
 ANTENNAPARTIALMETALAREA                  0.805 LAYER ME1 ;
 ANTENNAGATEAREA                          0.072 LAYER ME1 ;
 ANTENNAGATEAREA                          0.072 LAYER ME2 ;
 ANTENNAGATEAREA                          0.072 LAYER ME3 ;
 ANTENNAGATEAREA                          0.072 LAYER ME4 ;
 ANTENNADIFFAREA                          0.218 LAYER ME1 ;
 ANTENNADIFFAREA                          0.218 LAYER ME2 ;
 ANTENNADIFFAREA                          0.218 LAYER ME3 ;
 ANTENNADIFFAREA                          0.218 LAYER ME4 ;
 ANTENNAMAXAREACAR                       13.984 LAYER ME1 ;
 ANTENNAMAXAREACAR                       16.784 LAYER ME2 ;
 ANTENNAMAXAREACAR                       19.584 LAYER ME3 ;
 ANTENNAMAXAREACAR                       22.384 LAYER ME4 ;
END DI21
PIN DO21
  DIRECTION OUTPUT ;
 PORT
  LAYER ME4 ;
  RECT 174.796 0.000 175.076 0.720 ;
  LAYER ME3 ;
  RECT 174.796 0.000 175.076 0.720 ;
  LAYER ME2 ;
  RECT 174.796 0.000 175.076 0.720 ;
  LAYER ME1 ;
  RECT 174.796 0.000 175.076 0.720 ;
 END
 ANTENNAPARTIALMETALAREA                  2.030 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME3 ;
 ANTENNADIFFAREA                          1.293 LAYER ME4 ;
END DO21
PIN DI20
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 168.766 0.000 169.046 0.720 ;
  LAYER ME3 ;
  RECT 168.766 0.000 169.046 0.720 ;
  LAYER ME2 ;
  RECT 168.766 0.000 169.046 0.720 ;
  LAYER ME1 ;
  RECT 168.766 0.000 169.046 0.720 ;
 END
 ANTENNAPARTIALMETALAREA                  0.805 LAYER ME1 ;
 ANTENNAGATEAREA                          0.072 LAYER ME1 ;
 ANTENNAGATEAREA                          0.072 LAYER ME2 ;
 ANTENNAGATEAREA                          0.072 LAYER ME3 ;
 ANTENNAGATEAREA                          0.072 LAYER ME4 ;
 ANTENNADIFFAREA                          0.218 LAYER ME1 ;
 ANTENNADIFFAREA                          0.218 LAYER ME2 ;
 ANTENNADIFFAREA                          0.218 LAYER ME3 ;
 ANTENNADIFFAREA                          0.218 LAYER ME4 ;
 ANTENNAMAXAREACAR                       13.984 LAYER ME1 ;
 ANTENNAMAXAREACAR                       16.784 LAYER ME2 ;
 ANTENNAMAXAREACAR                       19.584 LAYER ME3 ;
 ANTENNAMAXAREACAR                       22.384 LAYER ME4 ;
END DI20
PIN DO20
  DIRECTION OUTPUT ;
 PORT
  LAYER ME4 ;
  RECT 166.788 0.000 167.068 0.720 ;
  LAYER ME3 ;
  RECT 166.788 0.000 167.068 0.720 ;
  LAYER ME2 ;
  RECT 166.788 0.000 167.068 0.720 ;
  LAYER ME1 ;
  RECT 166.788 0.000 167.068 0.720 ;
 END
 ANTENNAPARTIALMETALAREA                  2.030 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME3 ;
 ANTENNADIFFAREA                          1.293 LAYER ME4 ;
END DO20
PIN DI19
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 160.758 0.000 161.038 0.720 ;
  LAYER ME3 ;
  RECT 160.758 0.000 161.038 0.720 ;
  LAYER ME2 ;
  RECT 160.758 0.000 161.038 0.720 ;
  LAYER ME1 ;
  RECT 160.758 0.000 161.038 0.720 ;
 END
 ANTENNAPARTIALMETALAREA                  0.805 LAYER ME1 ;
 ANTENNAGATEAREA                          0.072 LAYER ME1 ;
 ANTENNAGATEAREA                          0.072 LAYER ME2 ;
 ANTENNAGATEAREA                          0.072 LAYER ME3 ;
 ANTENNAGATEAREA                          0.072 LAYER ME4 ;
 ANTENNADIFFAREA                          0.218 LAYER ME1 ;
 ANTENNADIFFAREA                          0.218 LAYER ME2 ;
 ANTENNADIFFAREA                          0.218 LAYER ME3 ;
 ANTENNADIFFAREA                          0.218 LAYER ME4 ;
 ANTENNAMAXAREACAR                       13.984 LAYER ME1 ;
 ANTENNAMAXAREACAR                       16.784 LAYER ME2 ;
 ANTENNAMAXAREACAR                       19.584 LAYER ME3 ;
 ANTENNAMAXAREACAR                       22.384 LAYER ME4 ;
END DI19
PIN DO19
  DIRECTION OUTPUT ;
 PORT
  LAYER ME4 ;
  RECT 158.780 0.000 159.060 0.720 ;
  LAYER ME3 ;
  RECT 158.780 0.000 159.060 0.720 ;
  LAYER ME2 ;
  RECT 158.780 0.000 159.060 0.720 ;
  LAYER ME1 ;
  RECT 158.780 0.000 159.060 0.720 ;
 END
 ANTENNAPARTIALMETALAREA                  2.030 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME3 ;
 ANTENNADIFFAREA                          1.293 LAYER ME4 ;
END DO19
PIN DI18
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 152.750 0.000 153.030 0.720 ;
  LAYER ME3 ;
  RECT 152.750 0.000 153.030 0.720 ;
  LAYER ME2 ;
  RECT 152.750 0.000 153.030 0.720 ;
  LAYER ME1 ;
  RECT 152.750 0.000 153.030 0.720 ;
 END
 ANTENNAPARTIALMETALAREA                  0.522 LAYER ME1 ;
 ANTENNAGATEAREA                          0.072 LAYER ME1 ;
 ANTENNAGATEAREA                          0.072 LAYER ME2 ;
 ANTENNAGATEAREA                          0.072 LAYER ME3 ;
 ANTENNAGATEAREA                          0.072 LAYER ME4 ;
 ANTENNADIFFAREA                          0.218 LAYER ME1 ;
 ANTENNADIFFAREA                          0.218 LAYER ME2 ;
 ANTENNADIFFAREA                          0.218 LAYER ME3 ;
 ANTENNADIFFAREA                          0.218 LAYER ME4 ;
 ANTENNAMAXAREACAR                       10.048 LAYER ME1 ;
 ANTENNAMAXAREACAR                       12.848 LAYER ME2 ;
 ANTENNAMAXAREACAR                       15.648 LAYER ME3 ;
 ANTENNAMAXAREACAR                       18.448 LAYER ME4 ;
END DI18
PIN DO18
  DIRECTION OUTPUT ;
 PORT
  LAYER ME4 ;
  RECT 150.692 0.000 150.972 0.720 ;
  LAYER ME3 ;
  RECT 150.692 0.000 150.972 0.720 ;
  LAYER ME2 ;
  RECT 150.692 0.000 150.972 0.720 ;
  LAYER ME1 ;
  RECT 150.692 0.000 150.972 0.720 ;
 END
 ANTENNAPARTIALMETALAREA                  2.030 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME3 ;
 ANTENNADIFFAREA                          1.293 LAYER ME4 ;
END DO18
PIN WEB2
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 151.172 0.000 151.452 0.720 ;
  LAYER ME3 ;
  RECT 151.172 0.000 151.452 0.720 ;
  LAYER ME2 ;
  RECT 151.172 0.000 151.452 0.720 ;
  LAYER ME1 ;
  RECT 151.172 0.000 151.452 0.720 ;
 END
 ANTENNAPARTIALMETALAREA                  0.436 LAYER ME2 ;
 ANTENNAGATEAREA                          0.288 LAYER ME2 ;
 ANTENNAGATEAREA                          0.288 LAYER ME3 ;
 ANTENNAGATEAREA                          0.288 LAYER ME4 ;
 ANTENNADIFFAREA                          0.218 LAYER ME2 ;
 ANTENNADIFFAREA                          0.218 LAYER ME3 ;
 ANTENNADIFFAREA                          0.218 LAYER ME4 ;
 ANTENNAMAXAREACAR                        4.602 LAYER ME2 ;
 ANTENNAMAXAREACAR                        5.302 LAYER ME3 ;
 ANTENNAMAXAREACAR                        6.002 LAYER ME4 ;
END WEB2
PIN DI17
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 144.742 0.000 145.022 0.720 ;
  LAYER ME3 ;
  RECT 144.742 0.000 145.022 0.720 ;
  LAYER ME2 ;
  RECT 144.742 0.000 145.022 0.720 ;
  LAYER ME1 ;
  RECT 144.742 0.000 145.022 0.720 ;
 END
 ANTENNAPARTIALMETALAREA                  0.805 LAYER ME1 ;
 ANTENNAGATEAREA                          0.072 LAYER ME1 ;
 ANTENNAGATEAREA                          0.072 LAYER ME2 ;
 ANTENNAGATEAREA                          0.072 LAYER ME3 ;
 ANTENNAGATEAREA                          0.072 LAYER ME4 ;
 ANTENNADIFFAREA                          0.218 LAYER ME1 ;
 ANTENNADIFFAREA                          0.218 LAYER ME2 ;
 ANTENNADIFFAREA                          0.218 LAYER ME3 ;
 ANTENNADIFFAREA                          0.218 LAYER ME4 ;
 ANTENNAMAXAREACAR                       13.984 LAYER ME1 ;
 ANTENNAMAXAREACAR                       16.784 LAYER ME2 ;
 ANTENNAMAXAREACAR                       19.584 LAYER ME3 ;
 ANTENNAMAXAREACAR                       22.384 LAYER ME4 ;
END DI17
PIN DO17
  DIRECTION OUTPUT ;
 PORT
  LAYER ME4 ;
  RECT 142.764 0.000 143.044 0.720 ;
  LAYER ME3 ;
  RECT 142.764 0.000 143.044 0.720 ;
  LAYER ME2 ;
  RECT 142.764 0.000 143.044 0.720 ;
  LAYER ME1 ;
  RECT 142.764 0.000 143.044 0.720 ;
 END
 ANTENNAPARTIALMETALAREA                  2.030 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME3 ;
 ANTENNADIFFAREA                          1.293 LAYER ME4 ;
END DO17
PIN DI16
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 136.734 0.000 137.014 0.720 ;
  LAYER ME3 ;
  RECT 136.734 0.000 137.014 0.720 ;
  LAYER ME2 ;
  RECT 136.734 0.000 137.014 0.720 ;
  LAYER ME1 ;
  RECT 136.734 0.000 137.014 0.720 ;
 END
 ANTENNAPARTIALMETALAREA                  0.805 LAYER ME1 ;
 ANTENNAGATEAREA                          0.072 LAYER ME1 ;
 ANTENNAGATEAREA                          0.072 LAYER ME2 ;
 ANTENNAGATEAREA                          0.072 LAYER ME3 ;
 ANTENNAGATEAREA                          0.072 LAYER ME4 ;
 ANTENNADIFFAREA                          0.218 LAYER ME1 ;
 ANTENNADIFFAREA                          0.218 LAYER ME2 ;
 ANTENNADIFFAREA                          0.218 LAYER ME3 ;
 ANTENNADIFFAREA                          0.218 LAYER ME4 ;
 ANTENNAMAXAREACAR                       13.984 LAYER ME1 ;
 ANTENNAMAXAREACAR                       16.784 LAYER ME2 ;
 ANTENNAMAXAREACAR                       19.584 LAYER ME3 ;
 ANTENNAMAXAREACAR                       22.384 LAYER ME4 ;
END DI16
PIN DO16
  DIRECTION OUTPUT ;
 PORT
  LAYER ME4 ;
  RECT 134.756 0.000 135.036 0.720 ;
  LAYER ME3 ;
  RECT 134.756 0.000 135.036 0.720 ;
  LAYER ME2 ;
  RECT 134.756 0.000 135.036 0.720 ;
  LAYER ME1 ;
  RECT 134.756 0.000 135.036 0.720 ;
 END
 ANTENNAPARTIALMETALAREA                  2.030 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME3 ;
 ANTENNADIFFAREA                          1.293 LAYER ME4 ;
END DO16
PIN DI15
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 128.726 0.000 129.006 0.720 ;
  LAYER ME3 ;
  RECT 128.726 0.000 129.006 0.720 ;
  LAYER ME2 ;
  RECT 128.726 0.000 129.006 0.720 ;
  LAYER ME1 ;
  RECT 128.726 0.000 129.006 0.720 ;
 END
 ANTENNAPARTIALMETALAREA                  0.805 LAYER ME1 ;
 ANTENNAGATEAREA                          0.072 LAYER ME1 ;
 ANTENNAGATEAREA                          0.072 LAYER ME2 ;
 ANTENNAGATEAREA                          0.072 LAYER ME3 ;
 ANTENNAGATEAREA                          0.072 LAYER ME4 ;
 ANTENNADIFFAREA                          0.218 LAYER ME1 ;
 ANTENNADIFFAREA                          0.218 LAYER ME2 ;
 ANTENNADIFFAREA                          0.218 LAYER ME3 ;
 ANTENNADIFFAREA                          0.218 LAYER ME4 ;
 ANTENNAMAXAREACAR                       13.984 LAYER ME1 ;
 ANTENNAMAXAREACAR                       16.784 LAYER ME2 ;
 ANTENNAMAXAREACAR                       19.584 LAYER ME3 ;
 ANTENNAMAXAREACAR                       22.384 LAYER ME4 ;
END DI15
PIN DO15
  DIRECTION OUTPUT ;
 PORT
  LAYER ME4 ;
  RECT 126.748 0.000 127.028 0.720 ;
  LAYER ME3 ;
  RECT 126.748 0.000 127.028 0.720 ;
  LAYER ME2 ;
  RECT 126.748 0.000 127.028 0.720 ;
  LAYER ME1 ;
  RECT 126.748 0.000 127.028 0.720 ;
 END
 ANTENNAPARTIALMETALAREA                  2.030 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME3 ;
 ANTENNADIFFAREA                          1.293 LAYER ME4 ;
END DO15
PIN DI14
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 120.718 0.000 120.998 0.720 ;
  LAYER ME3 ;
  RECT 120.718 0.000 120.998 0.720 ;
  LAYER ME2 ;
  RECT 120.718 0.000 120.998 0.720 ;
  LAYER ME1 ;
  RECT 120.718 0.000 120.998 0.720 ;
 END
 ANTENNAPARTIALMETALAREA                  0.805 LAYER ME1 ;
 ANTENNAGATEAREA                          0.072 LAYER ME1 ;
 ANTENNAGATEAREA                          0.072 LAYER ME2 ;
 ANTENNAGATEAREA                          0.072 LAYER ME3 ;
 ANTENNAGATEAREA                          0.072 LAYER ME4 ;
 ANTENNADIFFAREA                          0.218 LAYER ME1 ;
 ANTENNADIFFAREA                          0.218 LAYER ME2 ;
 ANTENNADIFFAREA                          0.218 LAYER ME3 ;
 ANTENNADIFFAREA                          0.218 LAYER ME4 ;
 ANTENNAMAXAREACAR                       13.984 LAYER ME1 ;
 ANTENNAMAXAREACAR                       16.784 LAYER ME2 ;
 ANTENNAMAXAREACAR                       19.584 LAYER ME3 ;
 ANTENNAMAXAREACAR                       22.384 LAYER ME4 ;
END DI14
PIN DO14
  DIRECTION OUTPUT ;
 PORT
  LAYER ME4 ;
  RECT 118.740 0.000 119.020 0.720 ;
  LAYER ME3 ;
  RECT 118.740 0.000 119.020 0.720 ;
  LAYER ME2 ;
  RECT 118.740 0.000 119.020 0.720 ;
  LAYER ME1 ;
  RECT 118.740 0.000 119.020 0.720 ;
 END
 ANTENNAPARTIALMETALAREA                  2.030 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME3 ;
 ANTENNADIFFAREA                          1.293 LAYER ME4 ;
END DO14
PIN DI13
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 112.710 0.000 112.990 0.720 ;
  LAYER ME3 ;
  RECT 112.710 0.000 112.990 0.720 ;
  LAYER ME2 ;
  RECT 112.710 0.000 112.990 0.720 ;
  LAYER ME1 ;
  RECT 112.710 0.000 112.990 0.720 ;
 END
 ANTENNAPARTIALMETALAREA                  0.805 LAYER ME1 ;
 ANTENNAGATEAREA                          0.072 LAYER ME1 ;
 ANTENNAGATEAREA                          0.072 LAYER ME2 ;
 ANTENNAGATEAREA                          0.072 LAYER ME3 ;
 ANTENNAGATEAREA                          0.072 LAYER ME4 ;
 ANTENNADIFFAREA                          0.218 LAYER ME1 ;
 ANTENNADIFFAREA                          0.218 LAYER ME2 ;
 ANTENNADIFFAREA                          0.218 LAYER ME3 ;
 ANTENNADIFFAREA                          0.218 LAYER ME4 ;
 ANTENNAMAXAREACAR                       13.984 LAYER ME1 ;
 ANTENNAMAXAREACAR                       16.784 LAYER ME2 ;
 ANTENNAMAXAREACAR                       19.584 LAYER ME3 ;
 ANTENNAMAXAREACAR                       22.384 LAYER ME4 ;
END DI13
PIN DO13
  DIRECTION OUTPUT ;
 PORT
  LAYER ME4 ;
  RECT 110.732 0.000 111.012 0.720 ;
  LAYER ME3 ;
  RECT 110.732 0.000 111.012 0.720 ;
  LAYER ME2 ;
  RECT 110.732 0.000 111.012 0.720 ;
  LAYER ME1 ;
  RECT 110.732 0.000 111.012 0.720 ;
 END
 ANTENNAPARTIALMETALAREA                  2.030 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME3 ;
 ANTENNADIFFAREA                          1.293 LAYER ME4 ;
END DO13
PIN DI12
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 104.702 0.000 104.982 0.720 ;
  LAYER ME3 ;
  RECT 104.702 0.000 104.982 0.720 ;
  LAYER ME2 ;
  RECT 104.702 0.000 104.982 0.720 ;
  LAYER ME1 ;
  RECT 104.702 0.000 104.982 0.720 ;
 END
 ANTENNAPARTIALMETALAREA                  0.805 LAYER ME1 ;
 ANTENNAGATEAREA                          0.072 LAYER ME1 ;
 ANTENNAGATEAREA                          0.072 LAYER ME2 ;
 ANTENNAGATEAREA                          0.072 LAYER ME3 ;
 ANTENNAGATEAREA                          0.072 LAYER ME4 ;
 ANTENNADIFFAREA                          0.218 LAYER ME1 ;
 ANTENNADIFFAREA                          0.218 LAYER ME2 ;
 ANTENNADIFFAREA                          0.218 LAYER ME3 ;
 ANTENNADIFFAREA                          0.218 LAYER ME4 ;
 ANTENNAMAXAREACAR                       13.984 LAYER ME1 ;
 ANTENNAMAXAREACAR                       16.784 LAYER ME2 ;
 ANTENNAMAXAREACAR                       19.584 LAYER ME3 ;
 ANTENNAMAXAREACAR                       22.384 LAYER ME4 ;
END DI12
PIN DO12
  DIRECTION OUTPUT ;
 PORT
  LAYER ME4 ;
  RECT 102.724 0.000 103.004 0.720 ;
  LAYER ME3 ;
  RECT 102.724 0.000 103.004 0.720 ;
  LAYER ME2 ;
  RECT 102.724 0.000 103.004 0.720 ;
  LAYER ME1 ;
  RECT 102.724 0.000 103.004 0.720 ;
 END
 ANTENNAPARTIALMETALAREA                  2.030 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME3 ;
 ANTENNADIFFAREA                          1.293 LAYER ME4 ;
END DO12
PIN DI11
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 96.694 0.000 96.974 0.720 ;
  LAYER ME3 ;
  RECT 96.694 0.000 96.974 0.720 ;
  LAYER ME2 ;
  RECT 96.694 0.000 96.974 0.720 ;
  LAYER ME1 ;
  RECT 96.694 0.000 96.974 0.720 ;
 END
 ANTENNAPARTIALMETALAREA                  0.805 LAYER ME1 ;
 ANTENNAGATEAREA                          0.072 LAYER ME1 ;
 ANTENNAGATEAREA                          0.072 LAYER ME2 ;
 ANTENNAGATEAREA                          0.072 LAYER ME3 ;
 ANTENNAGATEAREA                          0.072 LAYER ME4 ;
 ANTENNADIFFAREA                          0.218 LAYER ME1 ;
 ANTENNADIFFAREA                          0.218 LAYER ME2 ;
 ANTENNADIFFAREA                          0.218 LAYER ME3 ;
 ANTENNADIFFAREA                          0.218 LAYER ME4 ;
 ANTENNAMAXAREACAR                       13.984 LAYER ME1 ;
 ANTENNAMAXAREACAR                       16.784 LAYER ME2 ;
 ANTENNAMAXAREACAR                       19.584 LAYER ME3 ;
 ANTENNAMAXAREACAR                       22.384 LAYER ME4 ;
END DI11
PIN DO11
  DIRECTION OUTPUT ;
 PORT
  LAYER ME4 ;
  RECT 94.716 0.000 94.996 0.720 ;
  LAYER ME3 ;
  RECT 94.716 0.000 94.996 0.720 ;
  LAYER ME2 ;
  RECT 94.716 0.000 94.996 0.720 ;
  LAYER ME1 ;
  RECT 94.716 0.000 94.996 0.720 ;
 END
 ANTENNAPARTIALMETALAREA                  2.030 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME3 ;
 ANTENNADIFFAREA                          1.293 LAYER ME4 ;
END DO11
PIN DI10
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 88.686 0.000 88.966 0.720 ;
  LAYER ME3 ;
  RECT 88.686 0.000 88.966 0.720 ;
  LAYER ME2 ;
  RECT 88.686 0.000 88.966 0.720 ;
  LAYER ME1 ;
  RECT 88.686 0.000 88.966 0.720 ;
 END
 ANTENNAPARTIALMETALAREA                  0.805 LAYER ME1 ;
 ANTENNAGATEAREA                          0.072 LAYER ME1 ;
 ANTENNAGATEAREA                          0.072 LAYER ME2 ;
 ANTENNAGATEAREA                          0.072 LAYER ME3 ;
 ANTENNAGATEAREA                          0.072 LAYER ME4 ;
 ANTENNADIFFAREA                          0.218 LAYER ME1 ;
 ANTENNADIFFAREA                          0.218 LAYER ME2 ;
 ANTENNADIFFAREA                          0.218 LAYER ME3 ;
 ANTENNADIFFAREA                          0.218 LAYER ME4 ;
 ANTENNAMAXAREACAR                       13.984 LAYER ME1 ;
 ANTENNAMAXAREACAR                       16.784 LAYER ME2 ;
 ANTENNAMAXAREACAR                       19.584 LAYER ME3 ;
 ANTENNAMAXAREACAR                       22.384 LAYER ME4 ;
END DI10
PIN DO10
  DIRECTION OUTPUT ;
 PORT
  LAYER ME4 ;
  RECT 86.708 0.000 86.988 0.720 ;
  LAYER ME3 ;
  RECT 86.708 0.000 86.988 0.720 ;
  LAYER ME2 ;
  RECT 86.708 0.000 86.988 0.720 ;
  LAYER ME1 ;
  RECT 86.708 0.000 86.988 0.720 ;
 END
 ANTENNAPARTIALMETALAREA                  2.030 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME3 ;
 ANTENNADIFFAREA                          1.293 LAYER ME4 ;
END DO10
PIN DI9
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 80.678 0.000 80.958 0.720 ;
  LAYER ME3 ;
  RECT 80.678 0.000 80.958 0.720 ;
  LAYER ME2 ;
  RECT 80.678 0.000 80.958 0.720 ;
  LAYER ME1 ;
  RECT 80.678 0.000 80.958 0.720 ;
 END
 ANTENNAPARTIALMETALAREA                  0.522 LAYER ME1 ;
 ANTENNAGATEAREA                          0.072 LAYER ME1 ;
 ANTENNAGATEAREA                          0.072 LAYER ME2 ;
 ANTENNAGATEAREA                          0.072 LAYER ME3 ;
 ANTENNAGATEAREA                          0.072 LAYER ME4 ;
 ANTENNADIFFAREA                          0.218 LAYER ME1 ;
 ANTENNADIFFAREA                          0.218 LAYER ME2 ;
 ANTENNADIFFAREA                          0.218 LAYER ME3 ;
 ANTENNADIFFAREA                          0.218 LAYER ME4 ;
 ANTENNAMAXAREACAR                       10.048 LAYER ME1 ;
 ANTENNAMAXAREACAR                       12.848 LAYER ME2 ;
 ANTENNAMAXAREACAR                       15.648 LAYER ME3 ;
 ANTENNAMAXAREACAR                       18.448 LAYER ME4 ;
END DI9
PIN DO9
  DIRECTION OUTPUT ;
 PORT
  LAYER ME4 ;
  RECT 78.620 0.000 78.900 0.720 ;
  LAYER ME3 ;
  RECT 78.620 0.000 78.900 0.720 ;
  LAYER ME2 ;
  RECT 78.620 0.000 78.900 0.720 ;
  LAYER ME1 ;
  RECT 78.620 0.000 78.900 0.720 ;
 END
 ANTENNAPARTIALMETALAREA                  2.030 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME3 ;
 ANTENNADIFFAREA                          1.293 LAYER ME4 ;
END DO9
PIN WEB1
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 79.100 0.000 79.380 0.720 ;
  LAYER ME3 ;
  RECT 79.100 0.000 79.380 0.720 ;
  LAYER ME2 ;
  RECT 79.100 0.000 79.380 0.720 ;
  LAYER ME1 ;
  RECT 79.100 0.000 79.380 0.720 ;
 END
 ANTENNAPARTIALMETALAREA                  0.436 LAYER ME2 ;
 ANTENNAGATEAREA                          0.288 LAYER ME2 ;
 ANTENNAGATEAREA                          0.288 LAYER ME3 ;
 ANTENNAGATEAREA                          0.288 LAYER ME4 ;
 ANTENNADIFFAREA                          0.218 LAYER ME2 ;
 ANTENNADIFFAREA                          0.218 LAYER ME3 ;
 ANTENNADIFFAREA                          0.218 LAYER ME4 ;
 ANTENNAMAXAREACAR                        4.602 LAYER ME2 ;
 ANTENNAMAXAREACAR                        5.302 LAYER ME3 ;
 ANTENNAMAXAREACAR                        6.002 LAYER ME4 ;
END WEB1
PIN DI8
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 72.670 0.000 72.950 0.720 ;
  LAYER ME3 ;
  RECT 72.670 0.000 72.950 0.720 ;
  LAYER ME2 ;
  RECT 72.670 0.000 72.950 0.720 ;
  LAYER ME1 ;
  RECT 72.670 0.000 72.950 0.720 ;
 END
 ANTENNAPARTIALMETALAREA                  0.805 LAYER ME1 ;
 ANTENNAGATEAREA                          0.072 LAYER ME1 ;
 ANTENNAGATEAREA                          0.072 LAYER ME2 ;
 ANTENNAGATEAREA                          0.072 LAYER ME3 ;
 ANTENNAGATEAREA                          0.072 LAYER ME4 ;
 ANTENNADIFFAREA                          0.218 LAYER ME1 ;
 ANTENNADIFFAREA                          0.218 LAYER ME2 ;
 ANTENNADIFFAREA                          0.218 LAYER ME3 ;
 ANTENNADIFFAREA                          0.218 LAYER ME4 ;
 ANTENNAMAXAREACAR                       13.984 LAYER ME1 ;
 ANTENNAMAXAREACAR                       16.784 LAYER ME2 ;
 ANTENNAMAXAREACAR                       19.584 LAYER ME3 ;
 ANTENNAMAXAREACAR                       22.384 LAYER ME4 ;
END DI8
PIN DO8
  DIRECTION OUTPUT ;
 PORT
  LAYER ME4 ;
  RECT 70.692 0.000 70.972 0.720 ;
  LAYER ME3 ;
  RECT 70.692 0.000 70.972 0.720 ;
  LAYER ME2 ;
  RECT 70.692 0.000 70.972 0.720 ;
  LAYER ME1 ;
  RECT 70.692 0.000 70.972 0.720 ;
 END
 ANTENNAPARTIALMETALAREA                  2.030 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME3 ;
 ANTENNADIFFAREA                          1.293 LAYER ME4 ;
END DO8
PIN DI7
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 64.662 0.000 64.942 0.720 ;
  LAYER ME3 ;
  RECT 64.662 0.000 64.942 0.720 ;
  LAYER ME2 ;
  RECT 64.662 0.000 64.942 0.720 ;
  LAYER ME1 ;
  RECT 64.662 0.000 64.942 0.720 ;
 END
 ANTENNAPARTIALMETALAREA                  0.805 LAYER ME1 ;
 ANTENNAGATEAREA                          0.072 LAYER ME1 ;
 ANTENNAGATEAREA                          0.072 LAYER ME2 ;
 ANTENNAGATEAREA                          0.072 LAYER ME3 ;
 ANTENNAGATEAREA                          0.072 LAYER ME4 ;
 ANTENNADIFFAREA                          0.218 LAYER ME1 ;
 ANTENNADIFFAREA                          0.218 LAYER ME2 ;
 ANTENNADIFFAREA                          0.218 LAYER ME3 ;
 ANTENNADIFFAREA                          0.218 LAYER ME4 ;
 ANTENNAMAXAREACAR                       13.984 LAYER ME1 ;
 ANTENNAMAXAREACAR                       16.784 LAYER ME2 ;
 ANTENNAMAXAREACAR                       19.584 LAYER ME3 ;
 ANTENNAMAXAREACAR                       22.384 LAYER ME4 ;
END DI7
PIN DO7
  DIRECTION OUTPUT ;
 PORT
  LAYER ME4 ;
  RECT 62.684 0.000 62.964 0.720 ;
  LAYER ME3 ;
  RECT 62.684 0.000 62.964 0.720 ;
  LAYER ME2 ;
  RECT 62.684 0.000 62.964 0.720 ;
  LAYER ME1 ;
  RECT 62.684 0.000 62.964 0.720 ;
 END
 ANTENNAPARTIALMETALAREA                  2.030 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME3 ;
 ANTENNADIFFAREA                          1.293 LAYER ME4 ;
END DO7
PIN DI6
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 56.654 0.000 56.934 0.720 ;
  LAYER ME3 ;
  RECT 56.654 0.000 56.934 0.720 ;
  LAYER ME2 ;
  RECT 56.654 0.000 56.934 0.720 ;
  LAYER ME1 ;
  RECT 56.654 0.000 56.934 0.720 ;
 END
 ANTENNAPARTIALMETALAREA                  0.805 LAYER ME1 ;
 ANTENNAGATEAREA                          0.072 LAYER ME1 ;
 ANTENNAGATEAREA                          0.072 LAYER ME2 ;
 ANTENNAGATEAREA                          0.072 LAYER ME3 ;
 ANTENNAGATEAREA                          0.072 LAYER ME4 ;
 ANTENNADIFFAREA                          0.218 LAYER ME1 ;
 ANTENNADIFFAREA                          0.218 LAYER ME2 ;
 ANTENNADIFFAREA                          0.218 LAYER ME3 ;
 ANTENNADIFFAREA                          0.218 LAYER ME4 ;
 ANTENNAMAXAREACAR                       13.984 LAYER ME1 ;
 ANTENNAMAXAREACAR                       16.784 LAYER ME2 ;
 ANTENNAMAXAREACAR                       19.584 LAYER ME3 ;
 ANTENNAMAXAREACAR                       22.384 LAYER ME4 ;
END DI6
PIN DO6
  DIRECTION OUTPUT ;
 PORT
  LAYER ME4 ;
  RECT 54.676 0.000 54.956 0.720 ;
  LAYER ME3 ;
  RECT 54.676 0.000 54.956 0.720 ;
  LAYER ME2 ;
  RECT 54.676 0.000 54.956 0.720 ;
  LAYER ME1 ;
  RECT 54.676 0.000 54.956 0.720 ;
 END
 ANTENNAPARTIALMETALAREA                  2.030 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME3 ;
 ANTENNADIFFAREA                          1.293 LAYER ME4 ;
END DO6
PIN DI5
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 48.646 0.000 48.926 0.720 ;
  LAYER ME3 ;
  RECT 48.646 0.000 48.926 0.720 ;
  LAYER ME2 ;
  RECT 48.646 0.000 48.926 0.720 ;
  LAYER ME1 ;
  RECT 48.646 0.000 48.926 0.720 ;
 END
 ANTENNAPARTIALMETALAREA                  0.805 LAYER ME1 ;
 ANTENNAGATEAREA                          0.072 LAYER ME1 ;
 ANTENNAGATEAREA                          0.072 LAYER ME2 ;
 ANTENNAGATEAREA                          0.072 LAYER ME3 ;
 ANTENNAGATEAREA                          0.072 LAYER ME4 ;
 ANTENNADIFFAREA                          0.218 LAYER ME1 ;
 ANTENNADIFFAREA                          0.218 LAYER ME2 ;
 ANTENNADIFFAREA                          0.218 LAYER ME3 ;
 ANTENNADIFFAREA                          0.218 LAYER ME4 ;
 ANTENNAMAXAREACAR                       13.984 LAYER ME1 ;
 ANTENNAMAXAREACAR                       16.784 LAYER ME2 ;
 ANTENNAMAXAREACAR                       19.584 LAYER ME3 ;
 ANTENNAMAXAREACAR                       22.384 LAYER ME4 ;
END DI5
PIN DO5
  DIRECTION OUTPUT ;
 PORT
  LAYER ME4 ;
  RECT 46.668 0.000 46.948 0.720 ;
  LAYER ME3 ;
  RECT 46.668 0.000 46.948 0.720 ;
  LAYER ME2 ;
  RECT 46.668 0.000 46.948 0.720 ;
  LAYER ME1 ;
  RECT 46.668 0.000 46.948 0.720 ;
 END
 ANTENNAPARTIALMETALAREA                  2.030 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME3 ;
 ANTENNADIFFAREA                          1.293 LAYER ME4 ;
END DO5
PIN DI4
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 40.638 0.000 40.918 0.720 ;
  LAYER ME3 ;
  RECT 40.638 0.000 40.918 0.720 ;
  LAYER ME2 ;
  RECT 40.638 0.000 40.918 0.720 ;
  LAYER ME1 ;
  RECT 40.638 0.000 40.918 0.720 ;
 END
 ANTENNAPARTIALMETALAREA                  0.805 LAYER ME1 ;
 ANTENNAGATEAREA                          0.072 LAYER ME1 ;
 ANTENNAGATEAREA                          0.072 LAYER ME2 ;
 ANTENNAGATEAREA                          0.072 LAYER ME3 ;
 ANTENNAGATEAREA                          0.072 LAYER ME4 ;
 ANTENNADIFFAREA                          0.218 LAYER ME1 ;
 ANTENNADIFFAREA                          0.218 LAYER ME2 ;
 ANTENNADIFFAREA                          0.218 LAYER ME3 ;
 ANTENNADIFFAREA                          0.218 LAYER ME4 ;
 ANTENNAMAXAREACAR                       13.984 LAYER ME1 ;
 ANTENNAMAXAREACAR                       16.784 LAYER ME2 ;
 ANTENNAMAXAREACAR                       19.584 LAYER ME3 ;
 ANTENNAMAXAREACAR                       22.384 LAYER ME4 ;
END DI4
PIN DO4
  DIRECTION OUTPUT ;
 PORT
  LAYER ME4 ;
  RECT 38.660 0.000 38.940 0.720 ;
  LAYER ME3 ;
  RECT 38.660 0.000 38.940 0.720 ;
  LAYER ME2 ;
  RECT 38.660 0.000 38.940 0.720 ;
  LAYER ME1 ;
  RECT 38.660 0.000 38.940 0.720 ;
 END
 ANTENNAPARTIALMETALAREA                  2.030 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME3 ;
 ANTENNADIFFAREA                          1.293 LAYER ME4 ;
END DO4
PIN DI3
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 32.630 0.000 32.910 0.720 ;
  LAYER ME3 ;
  RECT 32.630 0.000 32.910 0.720 ;
  LAYER ME2 ;
  RECT 32.630 0.000 32.910 0.720 ;
  LAYER ME1 ;
  RECT 32.630 0.000 32.910 0.720 ;
 END
 ANTENNAPARTIALMETALAREA                  0.805 LAYER ME1 ;
 ANTENNAGATEAREA                          0.072 LAYER ME1 ;
 ANTENNAGATEAREA                          0.072 LAYER ME2 ;
 ANTENNAGATEAREA                          0.072 LAYER ME3 ;
 ANTENNAGATEAREA                          0.072 LAYER ME4 ;
 ANTENNADIFFAREA                          0.218 LAYER ME1 ;
 ANTENNADIFFAREA                          0.218 LAYER ME2 ;
 ANTENNADIFFAREA                          0.218 LAYER ME3 ;
 ANTENNADIFFAREA                          0.218 LAYER ME4 ;
 ANTENNAMAXAREACAR                       13.984 LAYER ME1 ;
 ANTENNAMAXAREACAR                       16.784 LAYER ME2 ;
 ANTENNAMAXAREACAR                       19.584 LAYER ME3 ;
 ANTENNAMAXAREACAR                       22.384 LAYER ME4 ;
END DI3
PIN DO3
  DIRECTION OUTPUT ;
 PORT
  LAYER ME4 ;
  RECT 30.652 0.000 30.932 0.720 ;
  LAYER ME3 ;
  RECT 30.652 0.000 30.932 0.720 ;
  LAYER ME2 ;
  RECT 30.652 0.000 30.932 0.720 ;
  LAYER ME1 ;
  RECT 30.652 0.000 30.932 0.720 ;
 END
 ANTENNAPARTIALMETALAREA                  2.030 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME3 ;
 ANTENNADIFFAREA                          1.293 LAYER ME4 ;
END DO3
PIN DI2
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 24.622 0.000 24.902 0.720 ;
  LAYER ME3 ;
  RECT 24.622 0.000 24.902 0.720 ;
  LAYER ME2 ;
  RECT 24.622 0.000 24.902 0.720 ;
  LAYER ME1 ;
  RECT 24.622 0.000 24.902 0.720 ;
 END
 ANTENNAPARTIALMETALAREA                  0.805 LAYER ME1 ;
 ANTENNAGATEAREA                          0.072 LAYER ME1 ;
 ANTENNAGATEAREA                          0.072 LAYER ME2 ;
 ANTENNAGATEAREA                          0.072 LAYER ME3 ;
 ANTENNAGATEAREA                          0.072 LAYER ME4 ;
 ANTENNADIFFAREA                          0.218 LAYER ME1 ;
 ANTENNADIFFAREA                          0.218 LAYER ME2 ;
 ANTENNADIFFAREA                          0.218 LAYER ME3 ;
 ANTENNADIFFAREA                          0.218 LAYER ME4 ;
 ANTENNAMAXAREACAR                       13.984 LAYER ME1 ;
 ANTENNAMAXAREACAR                       16.784 LAYER ME2 ;
 ANTENNAMAXAREACAR                       19.584 LAYER ME3 ;
 ANTENNAMAXAREACAR                       22.384 LAYER ME4 ;
END DI2
PIN DO2
  DIRECTION OUTPUT ;
 PORT
  LAYER ME4 ;
  RECT 22.644 0.000 22.924 0.720 ;
  LAYER ME3 ;
  RECT 22.644 0.000 22.924 0.720 ;
  LAYER ME2 ;
  RECT 22.644 0.000 22.924 0.720 ;
  LAYER ME1 ;
  RECT 22.644 0.000 22.924 0.720 ;
 END
 ANTENNAPARTIALMETALAREA                  2.030 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME3 ;
 ANTENNADIFFAREA                          1.293 LAYER ME4 ;
END DO2
PIN DI1
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 16.614 0.000 16.894 0.720 ;
  LAYER ME3 ;
  RECT 16.614 0.000 16.894 0.720 ;
  LAYER ME2 ;
  RECT 16.614 0.000 16.894 0.720 ;
  LAYER ME1 ;
  RECT 16.614 0.000 16.894 0.720 ;
 END
 ANTENNAPARTIALMETALAREA                  0.805 LAYER ME1 ;
 ANTENNAGATEAREA                          0.072 LAYER ME1 ;
 ANTENNAGATEAREA                          0.072 LAYER ME2 ;
 ANTENNAGATEAREA                          0.072 LAYER ME3 ;
 ANTENNAGATEAREA                          0.072 LAYER ME4 ;
 ANTENNADIFFAREA                          0.218 LAYER ME1 ;
 ANTENNADIFFAREA                          0.218 LAYER ME2 ;
 ANTENNADIFFAREA                          0.218 LAYER ME3 ;
 ANTENNADIFFAREA                          0.218 LAYER ME4 ;
 ANTENNAMAXAREACAR                       13.984 LAYER ME1 ;
 ANTENNAMAXAREACAR                       16.784 LAYER ME2 ;
 ANTENNAMAXAREACAR                       19.584 LAYER ME3 ;
 ANTENNAMAXAREACAR                       22.384 LAYER ME4 ;
END DI1
PIN DO1
  DIRECTION OUTPUT ;
 PORT
  LAYER ME4 ;
  RECT 14.636 0.000 14.916 0.720 ;
  LAYER ME3 ;
  RECT 14.636 0.000 14.916 0.720 ;
  LAYER ME2 ;
  RECT 14.636 0.000 14.916 0.720 ;
  LAYER ME1 ;
  RECT 14.636 0.000 14.916 0.720 ;
 END
 ANTENNAPARTIALMETALAREA                  2.030 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME3 ;
 ANTENNADIFFAREA                          1.293 LAYER ME4 ;
END DO1
PIN DI0
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 8.606 0.000 8.886 0.720 ;
  LAYER ME3 ;
  RECT 8.606 0.000 8.886 0.720 ;
  LAYER ME2 ;
  RECT 8.606 0.000 8.886 0.720 ;
  LAYER ME1 ;
  RECT 8.606 0.000 8.886 0.720 ;
 END
 ANTENNAPARTIALMETALAREA                  0.522 LAYER ME1 ;
 ANTENNAGATEAREA                          0.072 LAYER ME1 ;
 ANTENNAGATEAREA                          0.072 LAYER ME2 ;
 ANTENNAGATEAREA                          0.072 LAYER ME3 ;
 ANTENNAGATEAREA                          0.072 LAYER ME4 ;
 ANTENNADIFFAREA                          0.218 LAYER ME1 ;
 ANTENNADIFFAREA                          0.218 LAYER ME2 ;
 ANTENNADIFFAREA                          0.218 LAYER ME3 ;
 ANTENNADIFFAREA                          0.218 LAYER ME4 ;
 ANTENNAMAXAREACAR                       10.048 LAYER ME1 ;
 ANTENNAMAXAREACAR                       12.848 LAYER ME2 ;
 ANTENNAMAXAREACAR                       15.648 LAYER ME3 ;
 ANTENNAMAXAREACAR                       18.448 LAYER ME4 ;
END DI0
PIN DO0
  DIRECTION OUTPUT ;
 PORT
  LAYER ME4 ;
  RECT 6.548 0.000 6.828 0.720 ;
  LAYER ME3 ;
  RECT 6.548 0.000 6.828 0.720 ;
  LAYER ME2 ;
  RECT 6.548 0.000 6.828 0.720 ;
  LAYER ME1 ;
  RECT 6.548 0.000 6.828 0.720 ;
 END
 ANTENNAPARTIALMETALAREA                  2.030 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME3 ;
 ANTENNADIFFAREA                          1.293 LAYER ME4 ;
END DO0
PIN WEB0
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 7.028 0.000 7.308 0.720 ;
  LAYER ME3 ;
  RECT 7.028 0.000 7.308 0.720 ;
  LAYER ME2 ;
  RECT 7.028 0.000 7.308 0.720 ;
  LAYER ME1 ;
  RECT 7.028 0.000 7.308 0.720 ;
 END
 ANTENNAPARTIALMETALAREA                  0.436 LAYER ME2 ;
 ANTENNAGATEAREA                          0.288 LAYER ME2 ;
 ANTENNAGATEAREA                          0.288 LAYER ME3 ;
 ANTENNAGATEAREA                          0.288 LAYER ME4 ;
 ANTENNADIFFAREA                          0.218 LAYER ME2 ;
 ANTENNADIFFAREA                          0.218 LAYER ME3 ;
 ANTENNADIFFAREA                          0.218 LAYER ME4 ;
 ANTENNAMAXAREACAR                        4.602 LAYER ME2 ;
 ANTENNAMAXAREACAR                        5.302 LAYER ME3 ;
 ANTENNAMAXAREACAR                        6.002 LAYER ME4 ;
END WEB0
PIN A2
  DIRECTION INPUT ;
 PORT
  LAYER ME3 ;
  RECT 307.172 0.000 307.492 0.600 ;
  LAYER ME2 ;
  RECT 307.172 0.000 307.492 0.600 ;
  LAYER ME1 ;
  RECT 307.172 0.000 307.492 0.600 ;
 END
 ANTENNAPARTIALMETALAREA                  1.067 LAYER ME2 ;
 ANTENNAGATEAREA                          0.144 LAYER ME2 ;
 ANTENNAGATEAREA                          0.144 LAYER ME3 ;
 ANTENNADIFFAREA                          0.218 LAYER ME2 ;
 ANTENNADIFFAREA                          0.218 LAYER ME3 ;
 ANTENNAMAXAREACAR                        9.746 LAYER ME2 ;
 ANTENNAMAXAREACAR                       11.079 LAYER ME3 ;
END A2
PIN A3
  DIRECTION INPUT ;
 PORT
  LAYER ME3 ;
  RECT 307.759 0.000 308.079 0.600 ;
  LAYER ME2 ;
  RECT 307.759 0.000 308.079 0.600 ;
  LAYER ME1 ;
  RECT 307.759 0.000 308.079 0.600 ;
 END
 ANTENNAPARTIALMETALAREA                  1.188 LAYER ME2 ;
 ANTENNAGATEAREA                          0.144 LAYER ME2 ;
 ANTENNAGATEAREA                          0.144 LAYER ME3 ;
 ANTENNADIFFAREA                          0.218 LAYER ME2 ;
 ANTENNADIFFAREA                          0.218 LAYER ME3 ;
 ANTENNAMAXAREACAR                       10.582 LAYER ME2 ;
 ANTENNAMAXAREACAR                       11.915 LAYER ME3 ;
END A3
PIN A4
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 300.920 0.000 301.240 0.600 ;
  LAYER ME3 ;
  RECT 300.920 0.000 301.240 0.600 ;
  LAYER ME2 ;
  RECT 300.920 0.000 301.240 0.600 ;
  LAYER ME1 ;
  RECT 300.920 0.000 301.240 0.600 ;
 END
 ANTENNAPARTIALMETALAREA                  1.910 LAYER ME2 ;
 ANTENNAGATEAREA                          0.180 LAYER ME2 ;
 ANTENNAGATEAREA                          0.180 LAYER ME3 ;
 ANTENNAGATEAREA                          0.180 LAYER ME4 ;
 ANTENNADIFFAREA                          0.218 LAYER ME2 ;
 ANTENNADIFFAREA                          0.218 LAYER ME3 ;
 ANTENNADIFFAREA                          0.218 LAYER ME4 ;
 ANTENNAMAXAREACAR                       13.456 LAYER ME2 ;
 ANTENNAMAXAREACAR                       14.522 LAYER ME3 ;
 ANTENNAMAXAREACAR                       15.589 LAYER ME4 ;
END A4
PIN A5
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 300.300 0.000 300.620 0.600 ;
  LAYER ME3 ;
  RECT 300.300 0.000 300.620 0.600 ;
  LAYER ME2 ;
  RECT 300.300 0.000 300.620 0.600 ;
  LAYER ME1 ;
  RECT 300.300 0.000 300.620 0.600 ;
 END
 ANTENNAPARTIALMETALAREA                  1.447 LAYER ME2 ;
 ANTENNAGATEAREA                          0.180 LAYER ME2 ;
 ANTENNAGATEAREA                          0.180 LAYER ME3 ;
 ANTENNAGATEAREA                          0.180 LAYER ME4 ;
 ANTENNADIFFAREA                          0.218 LAYER ME2 ;
 ANTENNADIFFAREA                          0.218 LAYER ME3 ;
 ANTENNADIFFAREA                          0.218 LAYER ME4 ;
 ANTENNAMAXAREACAR                       12.818 LAYER ME2 ;
 ANTENNAMAXAREACAR                       13.884 LAYER ME3 ;
 ANTENNAMAXAREACAR                       14.951 LAYER ME4 ;
END A5
PIN A6
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 296.760 0.000 297.080 0.600 ;
  LAYER ME3 ;
  RECT 296.760 0.000 297.080 0.600 ;
  LAYER ME2 ;
  RECT 296.760 0.000 297.080 0.600 ;
  LAYER ME1 ;
  RECT 296.760 0.000 297.080 0.600 ;
 END
 ANTENNAPARTIALMETALAREA                  1.910 LAYER ME2 ;
 ANTENNAGATEAREA                          0.180 LAYER ME2 ;
 ANTENNAGATEAREA                          0.180 LAYER ME3 ;
 ANTENNAGATEAREA                          0.180 LAYER ME4 ;
 ANTENNADIFFAREA                          0.218 LAYER ME2 ;
 ANTENNADIFFAREA                          0.218 LAYER ME3 ;
 ANTENNADIFFAREA                          0.218 LAYER ME4 ;
 ANTENNAMAXAREACAR                       13.456 LAYER ME2 ;
 ANTENNAMAXAREACAR                       14.522 LAYER ME3 ;
 ANTENNAMAXAREACAR                       15.589 LAYER ME4 ;
END A6
PIN A7
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 296.140 0.000 296.460 0.600 ;
  LAYER ME3 ;
  RECT 296.140 0.000 296.460 0.600 ;
  LAYER ME2 ;
  RECT 296.140 0.000 296.460 0.600 ;
  LAYER ME1 ;
  RECT 296.140 0.000 296.460 0.600 ;
 END
 ANTENNAPARTIALMETALAREA                  1.447 LAYER ME2 ;
 ANTENNAGATEAREA                          0.180 LAYER ME2 ;
 ANTENNAGATEAREA                          0.180 LAYER ME3 ;
 ANTENNAGATEAREA                          0.180 LAYER ME4 ;
 ANTENNADIFFAREA                          0.218 LAYER ME2 ;
 ANTENNADIFFAREA                          0.218 LAYER ME3 ;
 ANTENNADIFFAREA                          0.218 LAYER ME4 ;
 ANTENNAMAXAREACAR                       12.818 LAYER ME2 ;
 ANTENNAMAXAREACAR                       13.884 LAYER ME3 ;
 ANTENNAMAXAREACAR                       14.951 LAYER ME4 ;
END A7
PIN A1
  DIRECTION INPUT ;
 PORT
  LAYER ME3 ;
  RECT 312.045 0.000 312.365 0.712 ;
  LAYER ME2 ;
  RECT 312.045 0.000 312.365 0.712 ;
  LAYER ME1 ;
  RECT 312.045 0.000 312.365 0.712 ;
 END
 ANTENNAPARTIALMETALAREA                  3.219 LAYER ME2 ;
 ANTENNAGATEAREA                          0.108 LAYER ME2 ;
 ANTENNAGATEAREA                          0.108 LAYER ME3 ;
 ANTENNADIFFAREA                          0.218 LAYER ME2 ;
 ANTENNADIFFAREA                          0.218 LAYER ME3 ;
 ANTENNAMAXAREACAR                       33.245 LAYER ME2 ;
 ANTENNAMAXAREACAR                       35.355 LAYER ME3 ;
END A1
PIN A0
  DIRECTION INPUT ;
 PORT
  LAYER ME3 ;
  RECT 315.274 0.000 315.594 0.712 ;
  LAYER ME2 ;
  RECT 315.274 0.000 315.594 0.712 ;
  LAYER ME1 ;
  RECT 315.274 0.000 315.594 0.712 ;
 END
 ANTENNAPARTIALMETALAREA                  3.457 LAYER ME2 ;
 ANTENNAGATEAREA                          0.108 LAYER ME2 ;
 ANTENNAGATEAREA                          0.108 LAYER ME3 ;
 ANTENNADIFFAREA                          0.218 LAYER ME2 ;
 ANTENNADIFFAREA                          0.218 LAYER ME3 ;
 ANTENNAMAXAREACAR                       35.986 LAYER ME2 ;
 ANTENNAMAXAREACAR                       38.095 LAYER ME3 ;
END A0
PIN DVSE
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 327.865 0.000 328.185 0.717 ;
  LAYER ME3 ;
  RECT 327.865 0.000 328.185 0.717 ;
  LAYER ME3 ;
  RECT 327.865 0.000 328.185 0.717 ;
  LAYER ME2 ;
  RECT 327.865 0.000 328.185 0.717 ;
  LAYER ME2 ;
  RECT 327.865 0.000 328.185 0.717 ;
  LAYER ME1 ;
  RECT 327.865 0.000 328.185 0.717 ;
  LAYER ME1 ;
  RECT 327.865 0.000 328.185 0.717 ;
 END
 ANTENNAPARTIALMETALAREA                  5.305 LAYER ME2 ;
 ANTENNAGATEAREA                          0.612 LAYER ME2 ;
 ANTENNAGATEAREA                          0.612 LAYER ME3 ;
 ANTENNAGATEAREA                          0.612 LAYER ME4 ;
 ANTENNADIFFAREA                          0.218 LAYER ME2 ;
 ANTENNADIFFAREA                          0.218 LAYER ME3 ;
 ANTENNADIFFAREA                          0.218 LAYER ME4 ;
 ANTENNAMAXAREACAR                       53.132 LAYER ME2 ;
 ANTENNAMAXAREACAR                       55.256 LAYER ME3 ;
 ANTENNAMAXAREACAR                       57.381 LAYER ME4 ;
END DVSE
PIN DVS3
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 327.345 0.000 327.665 0.717 ;
  LAYER ME3 ;
  RECT 327.345 0.000 327.665 0.717 ;
  LAYER ME3 ;
  RECT 327.345 0.000 327.665 0.717 ;
  LAYER ME2 ;
  RECT 327.345 0.000 327.665 0.717 ;
  LAYER ME2 ;
  RECT 327.345 0.000 327.665 0.717 ;
  LAYER ME1 ;
  RECT 327.345 0.000 327.665 0.717 ;
  LAYER ME1 ;
  RECT 327.345 0.000 327.665 0.717 ;
 END
 ANTENNAPARTIALMETALAREA                  3.675 LAYER ME2 ;
 ANTENNAGATEAREA                          0.108 LAYER ME2 ;
 ANTENNAGATEAREA                          0.108 LAYER ME3 ;
 ANTENNAGATEAREA                          0.108 LAYER ME4 ;
 ANTENNADIFFAREA                          0.218 LAYER ME2 ;
 ANTENNADIFFAREA                          0.218 LAYER ME3 ;
 ANTENNADIFFAREA                          0.218 LAYER ME4 ;
 ANTENNAMAXAREACAR                       45.625 LAYER ME2 ;
 ANTENNAMAXAREACAR                       47.749 LAYER ME3 ;
 ANTENNAMAXAREACAR                       49.874 LAYER ME4 ;
END DVS3
PIN DVS2
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 328.385 0.000 328.705 0.717 ;
  LAYER ME3 ;
  RECT 328.385 0.000 328.705 0.717 ;
  LAYER ME3 ;
  RECT 328.385 0.000 328.705 0.717 ;
  LAYER ME2 ;
  RECT 328.385 0.000 328.705 0.717 ;
  LAYER ME2 ;
  RECT 328.385 0.000 328.705 0.717 ;
  LAYER ME1 ;
  RECT 328.385 0.000 328.705 0.717 ;
  LAYER ME1 ;
  RECT 328.385 0.000 328.705 0.717 ;
 END
 ANTENNAPARTIALMETALAREA                  5.371 LAYER ME2 ;
 ANTENNAGATEAREA                          0.108 LAYER ME2 ;
 ANTENNAGATEAREA                          0.108 LAYER ME3 ;
 ANTENNAGATEAREA                          0.108 LAYER ME4 ;
 ANTENNADIFFAREA                          0.218 LAYER ME2 ;
 ANTENNADIFFAREA                          0.218 LAYER ME3 ;
 ANTENNADIFFAREA                          0.218 LAYER ME4 ;
 ANTENNAMAXAREACAR                       60.060 LAYER ME2 ;
 ANTENNAMAXAREACAR                       62.184 LAYER ME3 ;
 ANTENNAMAXAREACAR                       64.309 LAYER ME4 ;
END DVS2
PIN DVS1
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 326.825 0.000 327.145 0.717 ;
  LAYER ME3 ;
  RECT 326.825 0.000 327.145 0.717 ;
  LAYER ME3 ;
  RECT 326.825 0.000 327.145 0.717 ;
  LAYER ME2 ;
  RECT 326.825 0.000 327.145 0.717 ;
  LAYER ME2 ;
  RECT 326.825 0.000 327.145 0.717 ;
  LAYER ME1 ;
  RECT 326.825 0.000 327.145 0.717 ;
  LAYER ME1 ;
  RECT 326.825 0.000 327.145 0.717 ;
 END
 ANTENNAPARTIALMETALAREA                  3.307 LAYER ME2 ;
 ANTENNAGATEAREA                          0.108 LAYER ME2 ;
 ANTENNAGATEAREA                          0.108 LAYER ME3 ;
 ANTENNAGATEAREA                          0.108 LAYER ME4 ;
 ANTENNADIFFAREA                          0.218 LAYER ME2 ;
 ANTENNADIFFAREA                          0.218 LAYER ME3 ;
 ANTENNADIFFAREA                          0.218 LAYER ME4 ;
 ANTENNAMAXAREACAR                       42.063 LAYER ME2 ;
 ANTENNAMAXAREACAR                       44.188 LAYER ME3 ;
 ANTENNAMAXAREACAR                       46.312 LAYER ME4 ;
END DVS1
PIN DVS0
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 328.905 0.000 329.225 0.693 ;
  LAYER ME3 ;
  RECT 328.905 0.000 329.225 0.693 ;
  LAYER ME3 ;
  RECT 328.905 0.000 329.225 0.693 ;
  LAYER ME2 ;
  RECT 328.905 0.000 329.225 0.693 ;
  LAYER ME2 ;
  RECT 328.905 0.000 329.225 0.693 ;
  LAYER ME1 ;
  RECT 328.905 0.000 329.225 0.693 ;
  LAYER ME1 ;
  RECT 328.905 0.000 329.225 0.693 ;
 END
 ANTENNAPARTIALMETALAREA                  4.376 LAYER ME2 ;
 ANTENNAGATEAREA                          0.108 LAYER ME2 ;
 ANTENNAGATEAREA                          0.108 LAYER ME3 ;
 ANTENNAGATEAREA                          0.108 LAYER ME4 ;
 ANTENNADIFFAREA                          0.218 LAYER ME2 ;
 ANTENNADIFFAREA                          0.218 LAYER ME3 ;
 ANTENNADIFFAREA                          0.218 LAYER ME4 ;
 ANTENNAMAXAREACAR                       53.260 LAYER ME2 ;
 ANTENNAMAXAREACAR                       55.313 LAYER ME3 ;
 ANTENNAMAXAREACAR                       57.367 LAYER ME4 ;
END DVS0
PIN CK
  DIRECTION INPUT ;
 PORT
  LAYER ME3 ;
  RECT 320.341 0.000 320.661 0.713 ;
  LAYER ME2 ;
  RECT 320.341 0.000 320.661 0.713 ;
  LAYER ME1 ;
  RECT 320.341 0.000 320.661 0.713 ;
 END
 ANTENNAPARTIALMETALAREA                  2.392 LAYER ME2 ;
 ANTENNAPARTIALMETALAREA                  7.363 LAYER ME3 ;
 ANTENNAGATEAREA                          0.072 LAYER ME2 ;
 ANTENNAGATEAREA                          1.260 LAYER ME3 ;
 ANTENNADIFFAREA                          0.218 LAYER ME2 ;
 ANTENNADIFFAREA                          0.218 LAYER ME3 ;
 ANTENNAMAXAREACAR                       46.148 LAYER ME2 ;
 ANTENNAMAXAREACAR                      151.587 LAYER ME3 ;
END CK
PIN CSB
  DIRECTION INPUT ;
 PORT
  LAYER ME3 ;
  RECT 313.553 0.000 313.873 0.712 ;
  LAYER ME2 ;
  RECT 313.553 0.000 313.873 0.712 ;
  LAYER ME1 ;
  RECT 313.553 0.000 313.873 0.712 ;
 END
 ANTENNAPARTIALMETALAREA                  3.350 LAYER ME2 ;
 ANTENNAPARTIALMETALAREA                  7.235 LAYER ME3 ;
 ANTENNAGATEAREA                          2.244 LAYER ME2 ;
 ANTENNAGATEAREA                          3.216 LAYER ME3 ;
 ANTENNADIFFAREA                          0.218 LAYER ME2 ;
 ANTENNADIFFAREA                          0.218 LAYER ME3 ;
 ANTENNAMAXAREACAR                       17.231 LAYER ME2 ;
 ANTENNAMAXAREACAR                       51.784 LAYER ME3 ;
END CSB
PIN DI71
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 614.851 0.000 615.131 0.720 ;
  LAYER ME3 ;
  RECT 614.851 0.000 615.131 0.720 ;
  LAYER ME2 ;
  RECT 614.851 0.000 615.131 0.720 ;
  LAYER ME1 ;
  RECT 614.851 0.000 615.131 0.720 ;
 END
 ANTENNAPARTIALMETALAREA                  0.805 LAYER ME1 ;
 ANTENNAGATEAREA                          0.072 LAYER ME1 ;
 ANTENNAGATEAREA                          0.072 LAYER ME2 ;
 ANTENNAGATEAREA                          0.072 LAYER ME3 ;
 ANTENNAGATEAREA                          0.072 LAYER ME4 ;
 ANTENNADIFFAREA                          0.218 LAYER ME1 ;
 ANTENNADIFFAREA                          0.218 LAYER ME2 ;
 ANTENNADIFFAREA                          0.218 LAYER ME3 ;
 ANTENNADIFFAREA                          0.218 LAYER ME4 ;
 ANTENNAMAXAREACAR                       13.984 LAYER ME1 ;
 ANTENNAMAXAREACAR                       16.784 LAYER ME2 ;
 ANTENNAMAXAREACAR                       19.584 LAYER ME3 ;
 ANTENNAMAXAREACAR                       22.384 LAYER ME4 ;
END DI71
PIN DO71
  DIRECTION OUTPUT ;
 PORT
  LAYER ME4 ;
  RECT 612.873 0.000 613.153 0.720 ;
  LAYER ME3 ;
  RECT 612.873 0.000 613.153 0.720 ;
  LAYER ME2 ;
  RECT 612.873 0.000 613.153 0.720 ;
  LAYER ME1 ;
  RECT 612.873 0.000 613.153 0.720 ;
 END
 ANTENNAPARTIALMETALAREA                  2.030 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME3 ;
 ANTENNADIFFAREA                          1.293 LAYER ME4 ;
END DO71
PIN DI70
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 606.843 0.000 607.123 0.720 ;
  LAYER ME3 ;
  RECT 606.843 0.000 607.123 0.720 ;
  LAYER ME2 ;
  RECT 606.843 0.000 607.123 0.720 ;
  LAYER ME1 ;
  RECT 606.843 0.000 607.123 0.720 ;
 END
 ANTENNAPARTIALMETALAREA                  0.805 LAYER ME1 ;
 ANTENNAGATEAREA                          0.072 LAYER ME1 ;
 ANTENNAGATEAREA                          0.072 LAYER ME2 ;
 ANTENNAGATEAREA                          0.072 LAYER ME3 ;
 ANTENNAGATEAREA                          0.072 LAYER ME4 ;
 ANTENNADIFFAREA                          0.218 LAYER ME1 ;
 ANTENNADIFFAREA                          0.218 LAYER ME2 ;
 ANTENNADIFFAREA                          0.218 LAYER ME3 ;
 ANTENNADIFFAREA                          0.218 LAYER ME4 ;
 ANTENNAMAXAREACAR                       13.984 LAYER ME1 ;
 ANTENNAMAXAREACAR                       16.784 LAYER ME2 ;
 ANTENNAMAXAREACAR                       19.584 LAYER ME3 ;
 ANTENNAMAXAREACAR                       22.384 LAYER ME4 ;
END DI70
PIN DO70
  DIRECTION OUTPUT ;
 PORT
  LAYER ME4 ;
  RECT 604.865 0.000 605.145 0.720 ;
  LAYER ME3 ;
  RECT 604.865 0.000 605.145 0.720 ;
  LAYER ME2 ;
  RECT 604.865 0.000 605.145 0.720 ;
  LAYER ME1 ;
  RECT 604.865 0.000 605.145 0.720 ;
 END
 ANTENNAPARTIALMETALAREA                  2.030 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME3 ;
 ANTENNADIFFAREA                          1.293 LAYER ME4 ;
END DO70
PIN DI69
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 598.835 0.000 599.115 0.720 ;
  LAYER ME3 ;
  RECT 598.835 0.000 599.115 0.720 ;
  LAYER ME2 ;
  RECT 598.835 0.000 599.115 0.720 ;
  LAYER ME1 ;
  RECT 598.835 0.000 599.115 0.720 ;
 END
 ANTENNAPARTIALMETALAREA                  0.805 LAYER ME1 ;
 ANTENNAGATEAREA                          0.072 LAYER ME1 ;
 ANTENNAGATEAREA                          0.072 LAYER ME2 ;
 ANTENNAGATEAREA                          0.072 LAYER ME3 ;
 ANTENNAGATEAREA                          0.072 LAYER ME4 ;
 ANTENNADIFFAREA                          0.218 LAYER ME1 ;
 ANTENNADIFFAREA                          0.218 LAYER ME2 ;
 ANTENNADIFFAREA                          0.218 LAYER ME3 ;
 ANTENNADIFFAREA                          0.218 LAYER ME4 ;
 ANTENNAMAXAREACAR                       13.984 LAYER ME1 ;
 ANTENNAMAXAREACAR                       16.784 LAYER ME2 ;
 ANTENNAMAXAREACAR                       19.584 LAYER ME3 ;
 ANTENNAMAXAREACAR                       22.384 LAYER ME4 ;
END DI69
PIN DO69
  DIRECTION OUTPUT ;
 PORT
  LAYER ME4 ;
  RECT 596.857 0.000 597.137 0.720 ;
  LAYER ME3 ;
  RECT 596.857 0.000 597.137 0.720 ;
  LAYER ME2 ;
  RECT 596.857 0.000 597.137 0.720 ;
  LAYER ME1 ;
  RECT 596.857 0.000 597.137 0.720 ;
 END
 ANTENNAPARTIALMETALAREA                  2.030 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME3 ;
 ANTENNADIFFAREA                          1.293 LAYER ME4 ;
END DO69
PIN DI68
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 590.827 0.000 591.107 0.720 ;
  LAYER ME3 ;
  RECT 590.827 0.000 591.107 0.720 ;
  LAYER ME2 ;
  RECT 590.827 0.000 591.107 0.720 ;
  LAYER ME1 ;
  RECT 590.827 0.000 591.107 0.720 ;
 END
 ANTENNAPARTIALMETALAREA                  0.805 LAYER ME1 ;
 ANTENNAGATEAREA                          0.072 LAYER ME1 ;
 ANTENNAGATEAREA                          0.072 LAYER ME2 ;
 ANTENNAGATEAREA                          0.072 LAYER ME3 ;
 ANTENNAGATEAREA                          0.072 LAYER ME4 ;
 ANTENNADIFFAREA                          0.218 LAYER ME1 ;
 ANTENNADIFFAREA                          0.218 LAYER ME2 ;
 ANTENNADIFFAREA                          0.218 LAYER ME3 ;
 ANTENNADIFFAREA                          0.218 LAYER ME4 ;
 ANTENNAMAXAREACAR                       13.984 LAYER ME1 ;
 ANTENNAMAXAREACAR                       16.784 LAYER ME2 ;
 ANTENNAMAXAREACAR                       19.584 LAYER ME3 ;
 ANTENNAMAXAREACAR                       22.384 LAYER ME4 ;
END DI68
PIN DO68
  DIRECTION OUTPUT ;
 PORT
  LAYER ME4 ;
  RECT 588.849 0.000 589.129 0.720 ;
  LAYER ME3 ;
  RECT 588.849 0.000 589.129 0.720 ;
  LAYER ME2 ;
  RECT 588.849 0.000 589.129 0.720 ;
  LAYER ME1 ;
  RECT 588.849 0.000 589.129 0.720 ;
 END
 ANTENNAPARTIALMETALAREA                  2.030 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME3 ;
 ANTENNADIFFAREA                          1.293 LAYER ME4 ;
END DO68
PIN DI67
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 582.819 0.000 583.099 0.720 ;
  LAYER ME3 ;
  RECT 582.819 0.000 583.099 0.720 ;
  LAYER ME2 ;
  RECT 582.819 0.000 583.099 0.720 ;
  LAYER ME1 ;
  RECT 582.819 0.000 583.099 0.720 ;
 END
 ANTENNAPARTIALMETALAREA                  0.805 LAYER ME1 ;
 ANTENNAGATEAREA                          0.072 LAYER ME1 ;
 ANTENNAGATEAREA                          0.072 LAYER ME2 ;
 ANTENNAGATEAREA                          0.072 LAYER ME3 ;
 ANTENNAGATEAREA                          0.072 LAYER ME4 ;
 ANTENNADIFFAREA                          0.218 LAYER ME1 ;
 ANTENNADIFFAREA                          0.218 LAYER ME2 ;
 ANTENNADIFFAREA                          0.218 LAYER ME3 ;
 ANTENNADIFFAREA                          0.218 LAYER ME4 ;
 ANTENNAMAXAREACAR                       13.984 LAYER ME1 ;
 ANTENNAMAXAREACAR                       16.784 LAYER ME2 ;
 ANTENNAMAXAREACAR                       19.584 LAYER ME3 ;
 ANTENNAMAXAREACAR                       22.384 LAYER ME4 ;
END DI67
PIN DO67
  DIRECTION OUTPUT ;
 PORT
  LAYER ME4 ;
  RECT 580.841 0.000 581.121 0.720 ;
  LAYER ME3 ;
  RECT 580.841 0.000 581.121 0.720 ;
  LAYER ME2 ;
  RECT 580.841 0.000 581.121 0.720 ;
  LAYER ME1 ;
  RECT 580.841 0.000 581.121 0.720 ;
 END
 ANTENNAPARTIALMETALAREA                  2.030 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME3 ;
 ANTENNADIFFAREA                          1.293 LAYER ME4 ;
END DO67
PIN DI66
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 574.811 0.000 575.091 0.720 ;
  LAYER ME3 ;
  RECT 574.811 0.000 575.091 0.720 ;
  LAYER ME2 ;
  RECT 574.811 0.000 575.091 0.720 ;
  LAYER ME1 ;
  RECT 574.811 0.000 575.091 0.720 ;
 END
 ANTENNAPARTIALMETALAREA                  0.805 LAYER ME1 ;
 ANTENNAGATEAREA                          0.072 LAYER ME1 ;
 ANTENNAGATEAREA                          0.072 LAYER ME2 ;
 ANTENNAGATEAREA                          0.072 LAYER ME3 ;
 ANTENNAGATEAREA                          0.072 LAYER ME4 ;
 ANTENNADIFFAREA                          0.218 LAYER ME1 ;
 ANTENNADIFFAREA                          0.218 LAYER ME2 ;
 ANTENNADIFFAREA                          0.218 LAYER ME3 ;
 ANTENNADIFFAREA                          0.218 LAYER ME4 ;
 ANTENNAMAXAREACAR                       13.984 LAYER ME1 ;
 ANTENNAMAXAREACAR                       16.784 LAYER ME2 ;
 ANTENNAMAXAREACAR                       19.584 LAYER ME3 ;
 ANTENNAMAXAREACAR                       22.384 LAYER ME4 ;
END DI66
PIN DO66
  DIRECTION OUTPUT ;
 PORT
  LAYER ME4 ;
  RECT 572.833 0.000 573.113 0.720 ;
  LAYER ME3 ;
  RECT 572.833 0.000 573.113 0.720 ;
  LAYER ME2 ;
  RECT 572.833 0.000 573.113 0.720 ;
  LAYER ME1 ;
  RECT 572.833 0.000 573.113 0.720 ;
 END
 ANTENNAPARTIALMETALAREA                  2.030 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME3 ;
 ANTENNADIFFAREA                          1.293 LAYER ME4 ;
END DO66
PIN DI65
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 566.803 0.000 567.083 0.720 ;
  LAYER ME3 ;
  RECT 566.803 0.000 567.083 0.720 ;
  LAYER ME2 ;
  RECT 566.803 0.000 567.083 0.720 ;
  LAYER ME1 ;
  RECT 566.803 0.000 567.083 0.720 ;
 END
 ANTENNAPARTIALMETALAREA                  0.805 LAYER ME1 ;
 ANTENNAGATEAREA                          0.072 LAYER ME1 ;
 ANTENNAGATEAREA                          0.072 LAYER ME2 ;
 ANTENNAGATEAREA                          0.072 LAYER ME3 ;
 ANTENNAGATEAREA                          0.072 LAYER ME4 ;
 ANTENNADIFFAREA                          0.218 LAYER ME1 ;
 ANTENNADIFFAREA                          0.218 LAYER ME2 ;
 ANTENNADIFFAREA                          0.218 LAYER ME3 ;
 ANTENNADIFFAREA                          0.218 LAYER ME4 ;
 ANTENNAMAXAREACAR                       13.984 LAYER ME1 ;
 ANTENNAMAXAREACAR                       16.784 LAYER ME2 ;
 ANTENNAMAXAREACAR                       19.584 LAYER ME3 ;
 ANTENNAMAXAREACAR                       22.384 LAYER ME4 ;
END DI65
PIN DO65
  DIRECTION OUTPUT ;
 PORT
  LAYER ME4 ;
  RECT 564.825 0.000 565.105 0.720 ;
  LAYER ME3 ;
  RECT 564.825 0.000 565.105 0.720 ;
  LAYER ME2 ;
  RECT 564.825 0.000 565.105 0.720 ;
  LAYER ME1 ;
  RECT 564.825 0.000 565.105 0.720 ;
 END
 ANTENNAPARTIALMETALAREA                  2.030 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME3 ;
 ANTENNADIFFAREA                          1.293 LAYER ME4 ;
END DO65
PIN DI64
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 558.795 0.000 559.075 0.720 ;
  LAYER ME3 ;
  RECT 558.795 0.000 559.075 0.720 ;
  LAYER ME2 ;
  RECT 558.795 0.000 559.075 0.720 ;
  LAYER ME1 ;
  RECT 558.795 0.000 559.075 0.720 ;
 END
 ANTENNAPARTIALMETALAREA                  0.805 LAYER ME1 ;
 ANTENNAGATEAREA                          0.072 LAYER ME1 ;
 ANTENNAGATEAREA                          0.072 LAYER ME2 ;
 ANTENNAGATEAREA                          0.072 LAYER ME3 ;
 ANTENNAGATEAREA                          0.072 LAYER ME4 ;
 ANTENNADIFFAREA                          0.218 LAYER ME1 ;
 ANTENNADIFFAREA                          0.218 LAYER ME2 ;
 ANTENNADIFFAREA                          0.218 LAYER ME3 ;
 ANTENNADIFFAREA                          0.218 LAYER ME4 ;
 ANTENNAMAXAREACAR                       13.984 LAYER ME1 ;
 ANTENNAMAXAREACAR                       16.784 LAYER ME2 ;
 ANTENNAMAXAREACAR                       19.584 LAYER ME3 ;
 ANTENNAMAXAREACAR                       22.384 LAYER ME4 ;
END DI64
PIN DO64
  DIRECTION OUTPUT ;
 PORT
  LAYER ME4 ;
  RECT 556.817 0.000 557.097 0.720 ;
  LAYER ME3 ;
  RECT 556.817 0.000 557.097 0.720 ;
  LAYER ME2 ;
  RECT 556.817 0.000 557.097 0.720 ;
  LAYER ME1 ;
  RECT 556.817 0.000 557.097 0.720 ;
 END
 ANTENNAPARTIALMETALAREA                  2.030 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME3 ;
 ANTENNADIFFAREA                          1.293 LAYER ME4 ;
END DO64
PIN DI63
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 550.787 0.000 551.067 0.720 ;
  LAYER ME3 ;
  RECT 550.787 0.000 551.067 0.720 ;
  LAYER ME2 ;
  RECT 550.787 0.000 551.067 0.720 ;
  LAYER ME1 ;
  RECT 550.787 0.000 551.067 0.720 ;
 END
 ANTENNAPARTIALMETALAREA                  0.522 LAYER ME1 ;
 ANTENNAGATEAREA                          0.072 LAYER ME1 ;
 ANTENNAGATEAREA                          0.072 LAYER ME2 ;
 ANTENNAGATEAREA                          0.072 LAYER ME3 ;
 ANTENNAGATEAREA                          0.072 LAYER ME4 ;
 ANTENNADIFFAREA                          0.218 LAYER ME1 ;
 ANTENNADIFFAREA                          0.218 LAYER ME2 ;
 ANTENNADIFFAREA                          0.218 LAYER ME3 ;
 ANTENNADIFFAREA                          0.218 LAYER ME4 ;
 ANTENNAMAXAREACAR                       10.048 LAYER ME1 ;
 ANTENNAMAXAREACAR                       12.848 LAYER ME2 ;
 ANTENNAMAXAREACAR                       15.648 LAYER ME3 ;
 ANTENNAMAXAREACAR                       18.448 LAYER ME4 ;
END DI63
PIN DO63
  DIRECTION OUTPUT ;
 PORT
  LAYER ME4 ;
  RECT 548.729 0.000 549.009 0.720 ;
  LAYER ME3 ;
  RECT 548.729 0.000 549.009 0.720 ;
  LAYER ME2 ;
  RECT 548.729 0.000 549.009 0.720 ;
  LAYER ME1 ;
  RECT 548.729 0.000 549.009 0.720 ;
 END
 ANTENNAPARTIALMETALAREA                  2.030 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME3 ;
 ANTENNADIFFAREA                          1.293 LAYER ME4 ;
END DO63
PIN WEB7
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 549.209 0.000 549.489 0.720 ;
  LAYER ME3 ;
  RECT 549.209 0.000 549.489 0.720 ;
  LAYER ME2 ;
  RECT 549.209 0.000 549.489 0.720 ;
  LAYER ME1 ;
  RECT 549.209 0.000 549.489 0.720 ;
 END
 ANTENNAPARTIALMETALAREA                  0.436 LAYER ME2 ;
 ANTENNAGATEAREA                          0.288 LAYER ME2 ;
 ANTENNAGATEAREA                          0.288 LAYER ME3 ;
 ANTENNAGATEAREA                          0.288 LAYER ME4 ;
 ANTENNADIFFAREA                          0.218 LAYER ME2 ;
 ANTENNADIFFAREA                          0.218 LAYER ME3 ;
 ANTENNADIFFAREA                          0.218 LAYER ME4 ;
 ANTENNAMAXAREACAR                        4.602 LAYER ME2 ;
 ANTENNAMAXAREACAR                        5.302 LAYER ME3 ;
 ANTENNAMAXAREACAR                        6.002 LAYER ME4 ;
END WEB7
PIN DI62
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 542.779 0.000 543.059 0.720 ;
  LAYER ME3 ;
  RECT 542.779 0.000 543.059 0.720 ;
  LAYER ME2 ;
  RECT 542.779 0.000 543.059 0.720 ;
  LAYER ME1 ;
  RECT 542.779 0.000 543.059 0.720 ;
 END
 ANTENNAPARTIALMETALAREA                  0.805 LAYER ME1 ;
 ANTENNAGATEAREA                          0.072 LAYER ME1 ;
 ANTENNAGATEAREA                          0.072 LAYER ME2 ;
 ANTENNAGATEAREA                          0.072 LAYER ME3 ;
 ANTENNAGATEAREA                          0.072 LAYER ME4 ;
 ANTENNADIFFAREA                          0.218 LAYER ME1 ;
 ANTENNADIFFAREA                          0.218 LAYER ME2 ;
 ANTENNADIFFAREA                          0.218 LAYER ME3 ;
 ANTENNADIFFAREA                          0.218 LAYER ME4 ;
 ANTENNAMAXAREACAR                       13.984 LAYER ME1 ;
 ANTENNAMAXAREACAR                       16.784 LAYER ME2 ;
 ANTENNAMAXAREACAR                       19.584 LAYER ME3 ;
 ANTENNAMAXAREACAR                       22.384 LAYER ME4 ;
END DI62
PIN DO62
  DIRECTION OUTPUT ;
 PORT
  LAYER ME4 ;
  RECT 540.801 0.000 541.081 0.720 ;
  LAYER ME3 ;
  RECT 540.801 0.000 541.081 0.720 ;
  LAYER ME2 ;
  RECT 540.801 0.000 541.081 0.720 ;
  LAYER ME1 ;
  RECT 540.801 0.000 541.081 0.720 ;
 END
 ANTENNAPARTIALMETALAREA                  2.030 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME3 ;
 ANTENNADIFFAREA                          1.293 LAYER ME4 ;
END DO62
PIN DI61
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 534.771 0.000 535.051 0.720 ;
  LAYER ME3 ;
  RECT 534.771 0.000 535.051 0.720 ;
  LAYER ME2 ;
  RECT 534.771 0.000 535.051 0.720 ;
  LAYER ME1 ;
  RECT 534.771 0.000 535.051 0.720 ;
 END
 ANTENNAPARTIALMETALAREA                  0.805 LAYER ME1 ;
 ANTENNAGATEAREA                          0.072 LAYER ME1 ;
 ANTENNAGATEAREA                          0.072 LAYER ME2 ;
 ANTENNAGATEAREA                          0.072 LAYER ME3 ;
 ANTENNAGATEAREA                          0.072 LAYER ME4 ;
 ANTENNADIFFAREA                          0.218 LAYER ME1 ;
 ANTENNADIFFAREA                          0.218 LAYER ME2 ;
 ANTENNADIFFAREA                          0.218 LAYER ME3 ;
 ANTENNADIFFAREA                          0.218 LAYER ME4 ;
 ANTENNAMAXAREACAR                       13.984 LAYER ME1 ;
 ANTENNAMAXAREACAR                       16.784 LAYER ME2 ;
 ANTENNAMAXAREACAR                       19.584 LAYER ME3 ;
 ANTENNAMAXAREACAR                       22.384 LAYER ME4 ;
END DI61
PIN DO61
  DIRECTION OUTPUT ;
 PORT
  LAYER ME4 ;
  RECT 532.793 0.000 533.073 0.720 ;
  LAYER ME3 ;
  RECT 532.793 0.000 533.073 0.720 ;
  LAYER ME2 ;
  RECT 532.793 0.000 533.073 0.720 ;
  LAYER ME1 ;
  RECT 532.793 0.000 533.073 0.720 ;
 END
 ANTENNAPARTIALMETALAREA                  2.030 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME3 ;
 ANTENNADIFFAREA                          1.293 LAYER ME4 ;
END DO61
PIN DI60
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 526.763 0.000 527.043 0.720 ;
  LAYER ME3 ;
  RECT 526.763 0.000 527.043 0.720 ;
  LAYER ME2 ;
  RECT 526.763 0.000 527.043 0.720 ;
  LAYER ME1 ;
  RECT 526.763 0.000 527.043 0.720 ;
 END
 ANTENNAPARTIALMETALAREA                  0.805 LAYER ME1 ;
 ANTENNAGATEAREA                          0.072 LAYER ME1 ;
 ANTENNAGATEAREA                          0.072 LAYER ME2 ;
 ANTENNAGATEAREA                          0.072 LAYER ME3 ;
 ANTENNAGATEAREA                          0.072 LAYER ME4 ;
 ANTENNADIFFAREA                          0.218 LAYER ME1 ;
 ANTENNADIFFAREA                          0.218 LAYER ME2 ;
 ANTENNADIFFAREA                          0.218 LAYER ME3 ;
 ANTENNADIFFAREA                          0.218 LAYER ME4 ;
 ANTENNAMAXAREACAR                       13.984 LAYER ME1 ;
 ANTENNAMAXAREACAR                       16.784 LAYER ME2 ;
 ANTENNAMAXAREACAR                       19.584 LAYER ME3 ;
 ANTENNAMAXAREACAR                       22.384 LAYER ME4 ;
END DI60
PIN DO60
  DIRECTION OUTPUT ;
 PORT
  LAYER ME4 ;
  RECT 524.785 0.000 525.065 0.720 ;
  LAYER ME3 ;
  RECT 524.785 0.000 525.065 0.720 ;
  LAYER ME2 ;
  RECT 524.785 0.000 525.065 0.720 ;
  LAYER ME1 ;
  RECT 524.785 0.000 525.065 0.720 ;
 END
 ANTENNAPARTIALMETALAREA                  2.030 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME3 ;
 ANTENNADIFFAREA                          1.293 LAYER ME4 ;
END DO60
PIN DI59
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 518.755 0.000 519.035 0.720 ;
  LAYER ME3 ;
  RECT 518.755 0.000 519.035 0.720 ;
  LAYER ME2 ;
  RECT 518.755 0.000 519.035 0.720 ;
  LAYER ME1 ;
  RECT 518.755 0.000 519.035 0.720 ;
 END
 ANTENNAPARTIALMETALAREA                  0.805 LAYER ME1 ;
 ANTENNAGATEAREA                          0.072 LAYER ME1 ;
 ANTENNAGATEAREA                          0.072 LAYER ME2 ;
 ANTENNAGATEAREA                          0.072 LAYER ME3 ;
 ANTENNAGATEAREA                          0.072 LAYER ME4 ;
 ANTENNADIFFAREA                          0.218 LAYER ME1 ;
 ANTENNADIFFAREA                          0.218 LAYER ME2 ;
 ANTENNADIFFAREA                          0.218 LAYER ME3 ;
 ANTENNADIFFAREA                          0.218 LAYER ME4 ;
 ANTENNAMAXAREACAR                       13.984 LAYER ME1 ;
 ANTENNAMAXAREACAR                       16.784 LAYER ME2 ;
 ANTENNAMAXAREACAR                       19.584 LAYER ME3 ;
 ANTENNAMAXAREACAR                       22.384 LAYER ME4 ;
END DI59
PIN DO59
  DIRECTION OUTPUT ;
 PORT
  LAYER ME4 ;
  RECT 516.777 0.000 517.057 0.720 ;
  LAYER ME3 ;
  RECT 516.777 0.000 517.057 0.720 ;
  LAYER ME2 ;
  RECT 516.777 0.000 517.057 0.720 ;
  LAYER ME1 ;
  RECT 516.777 0.000 517.057 0.720 ;
 END
 ANTENNAPARTIALMETALAREA                  2.030 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME3 ;
 ANTENNADIFFAREA                          1.293 LAYER ME4 ;
END DO59
PIN DI58
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 510.747 0.000 511.027 0.720 ;
  LAYER ME3 ;
  RECT 510.747 0.000 511.027 0.720 ;
  LAYER ME2 ;
  RECT 510.747 0.000 511.027 0.720 ;
  LAYER ME1 ;
  RECT 510.747 0.000 511.027 0.720 ;
 END
 ANTENNAPARTIALMETALAREA                  0.805 LAYER ME1 ;
 ANTENNAGATEAREA                          0.072 LAYER ME1 ;
 ANTENNAGATEAREA                          0.072 LAYER ME2 ;
 ANTENNAGATEAREA                          0.072 LAYER ME3 ;
 ANTENNAGATEAREA                          0.072 LAYER ME4 ;
 ANTENNADIFFAREA                          0.218 LAYER ME1 ;
 ANTENNADIFFAREA                          0.218 LAYER ME2 ;
 ANTENNADIFFAREA                          0.218 LAYER ME3 ;
 ANTENNADIFFAREA                          0.218 LAYER ME4 ;
 ANTENNAMAXAREACAR                       13.984 LAYER ME1 ;
 ANTENNAMAXAREACAR                       16.784 LAYER ME2 ;
 ANTENNAMAXAREACAR                       19.584 LAYER ME3 ;
 ANTENNAMAXAREACAR                       22.384 LAYER ME4 ;
END DI58
PIN DO58
  DIRECTION OUTPUT ;
 PORT
  LAYER ME4 ;
  RECT 508.769 0.000 509.049 0.720 ;
  LAYER ME3 ;
  RECT 508.769 0.000 509.049 0.720 ;
  LAYER ME2 ;
  RECT 508.769 0.000 509.049 0.720 ;
  LAYER ME1 ;
  RECT 508.769 0.000 509.049 0.720 ;
 END
 ANTENNAPARTIALMETALAREA                  2.030 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME3 ;
 ANTENNADIFFAREA                          1.293 LAYER ME4 ;
END DO58
PIN DI57
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 502.739 0.000 503.019 0.720 ;
  LAYER ME3 ;
  RECT 502.739 0.000 503.019 0.720 ;
  LAYER ME2 ;
  RECT 502.739 0.000 503.019 0.720 ;
  LAYER ME1 ;
  RECT 502.739 0.000 503.019 0.720 ;
 END
 ANTENNAPARTIALMETALAREA                  0.805 LAYER ME1 ;
 ANTENNAGATEAREA                          0.072 LAYER ME1 ;
 ANTENNAGATEAREA                          0.072 LAYER ME2 ;
 ANTENNAGATEAREA                          0.072 LAYER ME3 ;
 ANTENNAGATEAREA                          0.072 LAYER ME4 ;
 ANTENNADIFFAREA                          0.218 LAYER ME1 ;
 ANTENNADIFFAREA                          0.218 LAYER ME2 ;
 ANTENNADIFFAREA                          0.218 LAYER ME3 ;
 ANTENNADIFFAREA                          0.218 LAYER ME4 ;
 ANTENNAMAXAREACAR                       13.984 LAYER ME1 ;
 ANTENNAMAXAREACAR                       16.784 LAYER ME2 ;
 ANTENNAMAXAREACAR                       19.584 LAYER ME3 ;
 ANTENNAMAXAREACAR                       22.384 LAYER ME4 ;
END DI57
PIN DO57
  DIRECTION OUTPUT ;
 PORT
  LAYER ME4 ;
  RECT 500.761 0.000 501.041 0.720 ;
  LAYER ME3 ;
  RECT 500.761 0.000 501.041 0.720 ;
  LAYER ME2 ;
  RECT 500.761 0.000 501.041 0.720 ;
  LAYER ME1 ;
  RECT 500.761 0.000 501.041 0.720 ;
 END
 ANTENNAPARTIALMETALAREA                  2.030 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME3 ;
 ANTENNADIFFAREA                          1.293 LAYER ME4 ;
END DO57
PIN DI56
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 494.731 0.000 495.011 0.720 ;
  LAYER ME3 ;
  RECT 494.731 0.000 495.011 0.720 ;
  LAYER ME2 ;
  RECT 494.731 0.000 495.011 0.720 ;
  LAYER ME1 ;
  RECT 494.731 0.000 495.011 0.720 ;
 END
 ANTENNAPARTIALMETALAREA                  0.805 LAYER ME1 ;
 ANTENNAGATEAREA                          0.072 LAYER ME1 ;
 ANTENNAGATEAREA                          0.072 LAYER ME2 ;
 ANTENNAGATEAREA                          0.072 LAYER ME3 ;
 ANTENNAGATEAREA                          0.072 LAYER ME4 ;
 ANTENNADIFFAREA                          0.218 LAYER ME1 ;
 ANTENNADIFFAREA                          0.218 LAYER ME2 ;
 ANTENNADIFFAREA                          0.218 LAYER ME3 ;
 ANTENNADIFFAREA                          0.218 LAYER ME4 ;
 ANTENNAMAXAREACAR                       13.984 LAYER ME1 ;
 ANTENNAMAXAREACAR                       16.784 LAYER ME2 ;
 ANTENNAMAXAREACAR                       19.584 LAYER ME3 ;
 ANTENNAMAXAREACAR                       22.384 LAYER ME4 ;
END DI56
PIN DO56
  DIRECTION OUTPUT ;
 PORT
  LAYER ME4 ;
  RECT 492.753 0.000 493.033 0.720 ;
  LAYER ME3 ;
  RECT 492.753 0.000 493.033 0.720 ;
  LAYER ME2 ;
  RECT 492.753 0.000 493.033 0.720 ;
  LAYER ME1 ;
  RECT 492.753 0.000 493.033 0.720 ;
 END
 ANTENNAPARTIALMETALAREA                  2.030 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME3 ;
 ANTENNADIFFAREA                          1.293 LAYER ME4 ;
END DO56
PIN DI55
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 486.723 0.000 487.003 0.720 ;
  LAYER ME3 ;
  RECT 486.723 0.000 487.003 0.720 ;
  LAYER ME2 ;
  RECT 486.723 0.000 487.003 0.720 ;
  LAYER ME1 ;
  RECT 486.723 0.000 487.003 0.720 ;
 END
 ANTENNAPARTIALMETALAREA                  0.805 LAYER ME1 ;
 ANTENNAGATEAREA                          0.072 LAYER ME1 ;
 ANTENNAGATEAREA                          0.072 LAYER ME2 ;
 ANTENNAGATEAREA                          0.072 LAYER ME3 ;
 ANTENNAGATEAREA                          0.072 LAYER ME4 ;
 ANTENNADIFFAREA                          0.218 LAYER ME1 ;
 ANTENNADIFFAREA                          0.218 LAYER ME2 ;
 ANTENNADIFFAREA                          0.218 LAYER ME3 ;
 ANTENNADIFFAREA                          0.218 LAYER ME4 ;
 ANTENNAMAXAREACAR                       13.984 LAYER ME1 ;
 ANTENNAMAXAREACAR                       16.784 LAYER ME2 ;
 ANTENNAMAXAREACAR                       19.584 LAYER ME3 ;
 ANTENNAMAXAREACAR                       22.384 LAYER ME4 ;
END DI55
PIN DO55
  DIRECTION OUTPUT ;
 PORT
  LAYER ME4 ;
  RECT 484.745 0.000 485.025 0.720 ;
  LAYER ME3 ;
  RECT 484.745 0.000 485.025 0.720 ;
  LAYER ME2 ;
  RECT 484.745 0.000 485.025 0.720 ;
  LAYER ME1 ;
  RECT 484.745 0.000 485.025 0.720 ;
 END
 ANTENNAPARTIALMETALAREA                  2.030 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME3 ;
 ANTENNADIFFAREA                          1.293 LAYER ME4 ;
END DO55
PIN DI54
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 478.715 0.000 478.995 0.720 ;
  LAYER ME3 ;
  RECT 478.715 0.000 478.995 0.720 ;
  LAYER ME2 ;
  RECT 478.715 0.000 478.995 0.720 ;
  LAYER ME1 ;
  RECT 478.715 0.000 478.995 0.720 ;
 END
 ANTENNAPARTIALMETALAREA                  0.522 LAYER ME1 ;
 ANTENNAGATEAREA                          0.072 LAYER ME1 ;
 ANTENNAGATEAREA                          0.072 LAYER ME2 ;
 ANTENNAGATEAREA                          0.072 LAYER ME3 ;
 ANTENNAGATEAREA                          0.072 LAYER ME4 ;
 ANTENNADIFFAREA                          0.218 LAYER ME1 ;
 ANTENNADIFFAREA                          0.218 LAYER ME2 ;
 ANTENNADIFFAREA                          0.218 LAYER ME3 ;
 ANTENNADIFFAREA                          0.218 LAYER ME4 ;
 ANTENNAMAXAREACAR                       10.048 LAYER ME1 ;
 ANTENNAMAXAREACAR                       12.848 LAYER ME2 ;
 ANTENNAMAXAREACAR                       15.648 LAYER ME3 ;
 ANTENNAMAXAREACAR                       18.448 LAYER ME4 ;
END DI54
PIN DO54
  DIRECTION OUTPUT ;
 PORT
  LAYER ME4 ;
  RECT 476.657 0.000 476.937 0.720 ;
  LAYER ME3 ;
  RECT 476.657 0.000 476.937 0.720 ;
  LAYER ME2 ;
  RECT 476.657 0.000 476.937 0.720 ;
  LAYER ME1 ;
  RECT 476.657 0.000 476.937 0.720 ;
 END
 ANTENNAPARTIALMETALAREA                  2.030 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME3 ;
 ANTENNADIFFAREA                          1.293 LAYER ME4 ;
END DO54
PIN WEB6
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 477.137 0.000 477.417 0.720 ;
  LAYER ME3 ;
  RECT 477.137 0.000 477.417 0.720 ;
  LAYER ME2 ;
  RECT 477.137 0.000 477.417 0.720 ;
  LAYER ME1 ;
  RECT 477.137 0.000 477.417 0.720 ;
 END
 ANTENNAPARTIALMETALAREA                  0.436 LAYER ME2 ;
 ANTENNAGATEAREA                          0.288 LAYER ME2 ;
 ANTENNAGATEAREA                          0.288 LAYER ME3 ;
 ANTENNAGATEAREA                          0.288 LAYER ME4 ;
 ANTENNADIFFAREA                          0.218 LAYER ME2 ;
 ANTENNADIFFAREA                          0.218 LAYER ME3 ;
 ANTENNADIFFAREA                          0.218 LAYER ME4 ;
 ANTENNAMAXAREACAR                        4.602 LAYER ME2 ;
 ANTENNAMAXAREACAR                        5.302 LAYER ME3 ;
 ANTENNAMAXAREACAR                        6.002 LAYER ME4 ;
END WEB6
PIN DI53
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 470.707 0.000 470.987 0.720 ;
  LAYER ME3 ;
  RECT 470.707 0.000 470.987 0.720 ;
  LAYER ME2 ;
  RECT 470.707 0.000 470.987 0.720 ;
  LAYER ME1 ;
  RECT 470.707 0.000 470.987 0.720 ;
 END
 ANTENNAPARTIALMETALAREA                  0.805 LAYER ME1 ;
 ANTENNAGATEAREA                          0.072 LAYER ME1 ;
 ANTENNAGATEAREA                          0.072 LAYER ME2 ;
 ANTENNAGATEAREA                          0.072 LAYER ME3 ;
 ANTENNAGATEAREA                          0.072 LAYER ME4 ;
 ANTENNADIFFAREA                          0.218 LAYER ME1 ;
 ANTENNADIFFAREA                          0.218 LAYER ME2 ;
 ANTENNADIFFAREA                          0.218 LAYER ME3 ;
 ANTENNADIFFAREA                          0.218 LAYER ME4 ;
 ANTENNAMAXAREACAR                       13.984 LAYER ME1 ;
 ANTENNAMAXAREACAR                       16.784 LAYER ME2 ;
 ANTENNAMAXAREACAR                       19.584 LAYER ME3 ;
 ANTENNAMAXAREACAR                       22.384 LAYER ME4 ;
END DI53
PIN DO53
  DIRECTION OUTPUT ;
 PORT
  LAYER ME4 ;
  RECT 468.729 0.000 469.009 0.720 ;
  LAYER ME3 ;
  RECT 468.729 0.000 469.009 0.720 ;
  LAYER ME2 ;
  RECT 468.729 0.000 469.009 0.720 ;
  LAYER ME1 ;
  RECT 468.729 0.000 469.009 0.720 ;
 END
 ANTENNAPARTIALMETALAREA                  2.030 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME3 ;
 ANTENNADIFFAREA                          1.293 LAYER ME4 ;
END DO53
PIN DI52
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 462.699 0.000 462.979 0.720 ;
  LAYER ME3 ;
  RECT 462.699 0.000 462.979 0.720 ;
  LAYER ME2 ;
  RECT 462.699 0.000 462.979 0.720 ;
  LAYER ME1 ;
  RECT 462.699 0.000 462.979 0.720 ;
 END
 ANTENNAPARTIALMETALAREA                  0.805 LAYER ME1 ;
 ANTENNAGATEAREA                          0.072 LAYER ME1 ;
 ANTENNAGATEAREA                          0.072 LAYER ME2 ;
 ANTENNAGATEAREA                          0.072 LAYER ME3 ;
 ANTENNAGATEAREA                          0.072 LAYER ME4 ;
 ANTENNADIFFAREA                          0.218 LAYER ME1 ;
 ANTENNADIFFAREA                          0.218 LAYER ME2 ;
 ANTENNADIFFAREA                          0.218 LAYER ME3 ;
 ANTENNADIFFAREA                          0.218 LAYER ME4 ;
 ANTENNAMAXAREACAR                       13.984 LAYER ME1 ;
 ANTENNAMAXAREACAR                       16.784 LAYER ME2 ;
 ANTENNAMAXAREACAR                       19.584 LAYER ME3 ;
 ANTENNAMAXAREACAR                       22.384 LAYER ME4 ;
END DI52
PIN DO52
  DIRECTION OUTPUT ;
 PORT
  LAYER ME4 ;
  RECT 460.721 0.000 461.001 0.720 ;
  LAYER ME3 ;
  RECT 460.721 0.000 461.001 0.720 ;
  LAYER ME2 ;
  RECT 460.721 0.000 461.001 0.720 ;
  LAYER ME1 ;
  RECT 460.721 0.000 461.001 0.720 ;
 END
 ANTENNAPARTIALMETALAREA                  2.030 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME3 ;
 ANTENNADIFFAREA                          1.293 LAYER ME4 ;
END DO52
PIN DI51
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 454.691 0.000 454.971 0.720 ;
  LAYER ME3 ;
  RECT 454.691 0.000 454.971 0.720 ;
  LAYER ME2 ;
  RECT 454.691 0.000 454.971 0.720 ;
  LAYER ME1 ;
  RECT 454.691 0.000 454.971 0.720 ;
 END
 ANTENNAPARTIALMETALAREA                  0.805 LAYER ME1 ;
 ANTENNAGATEAREA                          0.072 LAYER ME1 ;
 ANTENNAGATEAREA                          0.072 LAYER ME2 ;
 ANTENNAGATEAREA                          0.072 LAYER ME3 ;
 ANTENNAGATEAREA                          0.072 LAYER ME4 ;
 ANTENNADIFFAREA                          0.218 LAYER ME1 ;
 ANTENNADIFFAREA                          0.218 LAYER ME2 ;
 ANTENNADIFFAREA                          0.218 LAYER ME3 ;
 ANTENNADIFFAREA                          0.218 LAYER ME4 ;
 ANTENNAMAXAREACAR                       13.984 LAYER ME1 ;
 ANTENNAMAXAREACAR                       16.784 LAYER ME2 ;
 ANTENNAMAXAREACAR                       19.584 LAYER ME3 ;
 ANTENNAMAXAREACAR                       22.384 LAYER ME4 ;
END DI51
PIN DO51
  DIRECTION OUTPUT ;
 PORT
  LAYER ME4 ;
  RECT 452.713 0.000 452.993 0.720 ;
  LAYER ME3 ;
  RECT 452.713 0.000 452.993 0.720 ;
  LAYER ME2 ;
  RECT 452.713 0.000 452.993 0.720 ;
  LAYER ME1 ;
  RECT 452.713 0.000 452.993 0.720 ;
 END
 ANTENNAPARTIALMETALAREA                  2.030 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME3 ;
 ANTENNADIFFAREA                          1.293 LAYER ME4 ;
END DO51
PIN DI50
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 446.683 0.000 446.963 0.720 ;
  LAYER ME3 ;
  RECT 446.683 0.000 446.963 0.720 ;
  LAYER ME2 ;
  RECT 446.683 0.000 446.963 0.720 ;
  LAYER ME1 ;
  RECT 446.683 0.000 446.963 0.720 ;
 END
 ANTENNAPARTIALMETALAREA                  0.805 LAYER ME1 ;
 ANTENNAGATEAREA                          0.072 LAYER ME1 ;
 ANTENNAGATEAREA                          0.072 LAYER ME2 ;
 ANTENNAGATEAREA                          0.072 LAYER ME3 ;
 ANTENNAGATEAREA                          0.072 LAYER ME4 ;
 ANTENNADIFFAREA                          0.218 LAYER ME1 ;
 ANTENNADIFFAREA                          0.218 LAYER ME2 ;
 ANTENNADIFFAREA                          0.218 LAYER ME3 ;
 ANTENNADIFFAREA                          0.218 LAYER ME4 ;
 ANTENNAMAXAREACAR                       13.984 LAYER ME1 ;
 ANTENNAMAXAREACAR                       16.784 LAYER ME2 ;
 ANTENNAMAXAREACAR                       19.584 LAYER ME3 ;
 ANTENNAMAXAREACAR                       22.384 LAYER ME4 ;
END DI50
PIN DO50
  DIRECTION OUTPUT ;
 PORT
  LAYER ME4 ;
  RECT 444.705 0.000 444.985 0.720 ;
  LAYER ME3 ;
  RECT 444.705 0.000 444.985 0.720 ;
  LAYER ME2 ;
  RECT 444.705 0.000 444.985 0.720 ;
  LAYER ME1 ;
  RECT 444.705 0.000 444.985 0.720 ;
 END
 ANTENNAPARTIALMETALAREA                  2.030 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME3 ;
 ANTENNADIFFAREA                          1.293 LAYER ME4 ;
END DO50
PIN DI49
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 438.675 0.000 438.955 0.720 ;
  LAYER ME3 ;
  RECT 438.675 0.000 438.955 0.720 ;
  LAYER ME2 ;
  RECT 438.675 0.000 438.955 0.720 ;
  LAYER ME1 ;
  RECT 438.675 0.000 438.955 0.720 ;
 END
 ANTENNAPARTIALMETALAREA                  0.805 LAYER ME1 ;
 ANTENNAGATEAREA                          0.072 LAYER ME1 ;
 ANTENNAGATEAREA                          0.072 LAYER ME2 ;
 ANTENNAGATEAREA                          0.072 LAYER ME3 ;
 ANTENNAGATEAREA                          0.072 LAYER ME4 ;
 ANTENNADIFFAREA                          0.218 LAYER ME1 ;
 ANTENNADIFFAREA                          0.218 LAYER ME2 ;
 ANTENNADIFFAREA                          0.218 LAYER ME3 ;
 ANTENNADIFFAREA                          0.218 LAYER ME4 ;
 ANTENNAMAXAREACAR                       13.984 LAYER ME1 ;
 ANTENNAMAXAREACAR                       16.784 LAYER ME2 ;
 ANTENNAMAXAREACAR                       19.584 LAYER ME3 ;
 ANTENNAMAXAREACAR                       22.384 LAYER ME4 ;
END DI49
PIN DO49
  DIRECTION OUTPUT ;
 PORT
  LAYER ME4 ;
  RECT 436.697 0.000 436.977 0.720 ;
  LAYER ME3 ;
  RECT 436.697 0.000 436.977 0.720 ;
  LAYER ME2 ;
  RECT 436.697 0.000 436.977 0.720 ;
  LAYER ME1 ;
  RECT 436.697 0.000 436.977 0.720 ;
 END
 ANTENNAPARTIALMETALAREA                  2.030 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME3 ;
 ANTENNADIFFAREA                          1.293 LAYER ME4 ;
END DO49
PIN DI48
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 430.667 0.000 430.947 0.720 ;
  LAYER ME3 ;
  RECT 430.667 0.000 430.947 0.720 ;
  LAYER ME2 ;
  RECT 430.667 0.000 430.947 0.720 ;
  LAYER ME1 ;
  RECT 430.667 0.000 430.947 0.720 ;
 END
 ANTENNAPARTIALMETALAREA                  0.805 LAYER ME1 ;
 ANTENNAGATEAREA                          0.072 LAYER ME1 ;
 ANTENNAGATEAREA                          0.072 LAYER ME2 ;
 ANTENNAGATEAREA                          0.072 LAYER ME3 ;
 ANTENNAGATEAREA                          0.072 LAYER ME4 ;
 ANTENNADIFFAREA                          0.218 LAYER ME1 ;
 ANTENNADIFFAREA                          0.218 LAYER ME2 ;
 ANTENNADIFFAREA                          0.218 LAYER ME3 ;
 ANTENNADIFFAREA                          0.218 LAYER ME4 ;
 ANTENNAMAXAREACAR                       13.984 LAYER ME1 ;
 ANTENNAMAXAREACAR                       16.784 LAYER ME2 ;
 ANTENNAMAXAREACAR                       19.584 LAYER ME3 ;
 ANTENNAMAXAREACAR                       22.384 LAYER ME4 ;
END DI48
PIN DO48
  DIRECTION OUTPUT ;
 PORT
  LAYER ME4 ;
  RECT 428.689 0.000 428.969 0.720 ;
  LAYER ME3 ;
  RECT 428.689 0.000 428.969 0.720 ;
  LAYER ME2 ;
  RECT 428.689 0.000 428.969 0.720 ;
  LAYER ME1 ;
  RECT 428.689 0.000 428.969 0.720 ;
 END
 ANTENNAPARTIALMETALAREA                  2.030 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME3 ;
 ANTENNADIFFAREA                          1.293 LAYER ME4 ;
END DO48
PIN DI47
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 422.659 0.000 422.939 0.720 ;
  LAYER ME3 ;
  RECT 422.659 0.000 422.939 0.720 ;
  LAYER ME2 ;
  RECT 422.659 0.000 422.939 0.720 ;
  LAYER ME1 ;
  RECT 422.659 0.000 422.939 0.720 ;
 END
 ANTENNAPARTIALMETALAREA                  0.805 LAYER ME1 ;
 ANTENNAGATEAREA                          0.072 LAYER ME1 ;
 ANTENNAGATEAREA                          0.072 LAYER ME2 ;
 ANTENNAGATEAREA                          0.072 LAYER ME3 ;
 ANTENNAGATEAREA                          0.072 LAYER ME4 ;
 ANTENNADIFFAREA                          0.218 LAYER ME1 ;
 ANTENNADIFFAREA                          0.218 LAYER ME2 ;
 ANTENNADIFFAREA                          0.218 LAYER ME3 ;
 ANTENNADIFFAREA                          0.218 LAYER ME4 ;
 ANTENNAMAXAREACAR                       13.984 LAYER ME1 ;
 ANTENNAMAXAREACAR                       16.784 LAYER ME2 ;
 ANTENNAMAXAREACAR                       19.584 LAYER ME3 ;
 ANTENNAMAXAREACAR                       22.384 LAYER ME4 ;
END DI47
PIN DO47
  DIRECTION OUTPUT ;
 PORT
  LAYER ME4 ;
  RECT 420.681 0.000 420.961 0.720 ;
  LAYER ME3 ;
  RECT 420.681 0.000 420.961 0.720 ;
  LAYER ME2 ;
  RECT 420.681 0.000 420.961 0.720 ;
  LAYER ME1 ;
  RECT 420.681 0.000 420.961 0.720 ;
 END
 ANTENNAPARTIALMETALAREA                  2.030 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME3 ;
 ANTENNADIFFAREA                          1.293 LAYER ME4 ;
END DO47
PIN DI46
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 414.651 0.000 414.931 0.720 ;
  LAYER ME3 ;
  RECT 414.651 0.000 414.931 0.720 ;
  LAYER ME2 ;
  RECT 414.651 0.000 414.931 0.720 ;
  LAYER ME1 ;
  RECT 414.651 0.000 414.931 0.720 ;
 END
 ANTENNAPARTIALMETALAREA                  0.805 LAYER ME1 ;
 ANTENNAGATEAREA                          0.072 LAYER ME1 ;
 ANTENNAGATEAREA                          0.072 LAYER ME2 ;
 ANTENNAGATEAREA                          0.072 LAYER ME3 ;
 ANTENNAGATEAREA                          0.072 LAYER ME4 ;
 ANTENNADIFFAREA                          0.218 LAYER ME1 ;
 ANTENNADIFFAREA                          0.218 LAYER ME2 ;
 ANTENNADIFFAREA                          0.218 LAYER ME3 ;
 ANTENNADIFFAREA                          0.218 LAYER ME4 ;
 ANTENNAMAXAREACAR                       13.984 LAYER ME1 ;
 ANTENNAMAXAREACAR                       16.784 LAYER ME2 ;
 ANTENNAMAXAREACAR                       19.584 LAYER ME3 ;
 ANTENNAMAXAREACAR                       22.384 LAYER ME4 ;
END DI46
PIN DO46
  DIRECTION OUTPUT ;
 PORT
  LAYER ME4 ;
  RECT 412.673 0.000 412.953 0.720 ;
  LAYER ME3 ;
  RECT 412.673 0.000 412.953 0.720 ;
  LAYER ME2 ;
  RECT 412.673 0.000 412.953 0.720 ;
  LAYER ME1 ;
  RECT 412.673 0.000 412.953 0.720 ;
 END
 ANTENNAPARTIALMETALAREA                  2.030 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME3 ;
 ANTENNADIFFAREA                          1.293 LAYER ME4 ;
END DO46
PIN DI45
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 406.643 0.000 406.923 0.720 ;
  LAYER ME3 ;
  RECT 406.643 0.000 406.923 0.720 ;
  LAYER ME2 ;
  RECT 406.643 0.000 406.923 0.720 ;
  LAYER ME1 ;
  RECT 406.643 0.000 406.923 0.720 ;
 END
 ANTENNAPARTIALMETALAREA                  0.522 LAYER ME1 ;
 ANTENNAGATEAREA                          0.072 LAYER ME1 ;
 ANTENNAGATEAREA                          0.072 LAYER ME2 ;
 ANTENNAGATEAREA                          0.072 LAYER ME3 ;
 ANTENNAGATEAREA                          0.072 LAYER ME4 ;
 ANTENNADIFFAREA                          0.218 LAYER ME1 ;
 ANTENNADIFFAREA                          0.218 LAYER ME2 ;
 ANTENNADIFFAREA                          0.218 LAYER ME3 ;
 ANTENNADIFFAREA                          0.218 LAYER ME4 ;
 ANTENNAMAXAREACAR                       10.048 LAYER ME1 ;
 ANTENNAMAXAREACAR                       12.848 LAYER ME2 ;
 ANTENNAMAXAREACAR                       15.648 LAYER ME3 ;
 ANTENNAMAXAREACAR                       18.448 LAYER ME4 ;
END DI45
PIN DO45
  DIRECTION OUTPUT ;
 PORT
  LAYER ME4 ;
  RECT 404.585 0.000 404.865 0.720 ;
  LAYER ME3 ;
  RECT 404.585 0.000 404.865 0.720 ;
  LAYER ME2 ;
  RECT 404.585 0.000 404.865 0.720 ;
  LAYER ME1 ;
  RECT 404.585 0.000 404.865 0.720 ;
 END
 ANTENNAPARTIALMETALAREA                  2.030 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME3 ;
 ANTENNADIFFAREA                          1.293 LAYER ME4 ;
END DO45
PIN WEB5
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 405.065 0.000 405.345 0.720 ;
  LAYER ME3 ;
  RECT 405.065 0.000 405.345 0.720 ;
  LAYER ME2 ;
  RECT 405.065 0.000 405.345 0.720 ;
  LAYER ME1 ;
  RECT 405.065 0.000 405.345 0.720 ;
 END
 ANTENNAPARTIALMETALAREA                  0.436 LAYER ME2 ;
 ANTENNAGATEAREA                          0.288 LAYER ME2 ;
 ANTENNAGATEAREA                          0.288 LAYER ME3 ;
 ANTENNAGATEAREA                          0.288 LAYER ME4 ;
 ANTENNADIFFAREA                          0.218 LAYER ME2 ;
 ANTENNADIFFAREA                          0.218 LAYER ME3 ;
 ANTENNADIFFAREA                          0.218 LAYER ME4 ;
 ANTENNAMAXAREACAR                        4.602 LAYER ME2 ;
 ANTENNAMAXAREACAR                        5.302 LAYER ME3 ;
 ANTENNAMAXAREACAR                        6.002 LAYER ME4 ;
END WEB5
PIN DI44
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 398.635 0.000 398.915 0.720 ;
  LAYER ME3 ;
  RECT 398.635 0.000 398.915 0.720 ;
  LAYER ME2 ;
  RECT 398.635 0.000 398.915 0.720 ;
  LAYER ME1 ;
  RECT 398.635 0.000 398.915 0.720 ;
 END
 ANTENNAPARTIALMETALAREA                  0.805 LAYER ME1 ;
 ANTENNAGATEAREA                          0.072 LAYER ME1 ;
 ANTENNAGATEAREA                          0.072 LAYER ME2 ;
 ANTENNAGATEAREA                          0.072 LAYER ME3 ;
 ANTENNAGATEAREA                          0.072 LAYER ME4 ;
 ANTENNADIFFAREA                          0.218 LAYER ME1 ;
 ANTENNADIFFAREA                          0.218 LAYER ME2 ;
 ANTENNADIFFAREA                          0.218 LAYER ME3 ;
 ANTENNADIFFAREA                          0.218 LAYER ME4 ;
 ANTENNAMAXAREACAR                       13.984 LAYER ME1 ;
 ANTENNAMAXAREACAR                       16.784 LAYER ME2 ;
 ANTENNAMAXAREACAR                       19.584 LAYER ME3 ;
 ANTENNAMAXAREACAR                       22.384 LAYER ME4 ;
END DI44
PIN DO44
  DIRECTION OUTPUT ;
 PORT
  LAYER ME4 ;
  RECT 396.657 0.000 396.937 0.720 ;
  LAYER ME3 ;
  RECT 396.657 0.000 396.937 0.720 ;
  LAYER ME2 ;
  RECT 396.657 0.000 396.937 0.720 ;
  LAYER ME1 ;
  RECT 396.657 0.000 396.937 0.720 ;
 END
 ANTENNAPARTIALMETALAREA                  2.030 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME3 ;
 ANTENNADIFFAREA                          1.293 LAYER ME4 ;
END DO44
PIN DI43
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 390.627 0.000 390.907 0.720 ;
  LAYER ME3 ;
  RECT 390.627 0.000 390.907 0.720 ;
  LAYER ME2 ;
  RECT 390.627 0.000 390.907 0.720 ;
  LAYER ME1 ;
  RECT 390.627 0.000 390.907 0.720 ;
 END
 ANTENNAPARTIALMETALAREA                  0.805 LAYER ME1 ;
 ANTENNAGATEAREA                          0.072 LAYER ME1 ;
 ANTENNAGATEAREA                          0.072 LAYER ME2 ;
 ANTENNAGATEAREA                          0.072 LAYER ME3 ;
 ANTENNAGATEAREA                          0.072 LAYER ME4 ;
 ANTENNADIFFAREA                          0.218 LAYER ME1 ;
 ANTENNADIFFAREA                          0.218 LAYER ME2 ;
 ANTENNADIFFAREA                          0.218 LAYER ME3 ;
 ANTENNADIFFAREA                          0.218 LAYER ME4 ;
 ANTENNAMAXAREACAR                       13.984 LAYER ME1 ;
 ANTENNAMAXAREACAR                       16.784 LAYER ME2 ;
 ANTENNAMAXAREACAR                       19.584 LAYER ME3 ;
 ANTENNAMAXAREACAR                       22.384 LAYER ME4 ;
END DI43
PIN DO43
  DIRECTION OUTPUT ;
 PORT
  LAYER ME4 ;
  RECT 388.649 0.000 388.929 0.720 ;
  LAYER ME3 ;
  RECT 388.649 0.000 388.929 0.720 ;
  LAYER ME2 ;
  RECT 388.649 0.000 388.929 0.720 ;
  LAYER ME1 ;
  RECT 388.649 0.000 388.929 0.720 ;
 END
 ANTENNAPARTIALMETALAREA                  2.030 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME3 ;
 ANTENNADIFFAREA                          1.293 LAYER ME4 ;
END DO43
PIN DI42
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 382.619 0.000 382.899 0.720 ;
  LAYER ME3 ;
  RECT 382.619 0.000 382.899 0.720 ;
  LAYER ME2 ;
  RECT 382.619 0.000 382.899 0.720 ;
  LAYER ME1 ;
  RECT 382.619 0.000 382.899 0.720 ;
 END
 ANTENNAPARTIALMETALAREA                  0.805 LAYER ME1 ;
 ANTENNAGATEAREA                          0.072 LAYER ME1 ;
 ANTENNAGATEAREA                          0.072 LAYER ME2 ;
 ANTENNAGATEAREA                          0.072 LAYER ME3 ;
 ANTENNAGATEAREA                          0.072 LAYER ME4 ;
 ANTENNADIFFAREA                          0.218 LAYER ME1 ;
 ANTENNADIFFAREA                          0.218 LAYER ME2 ;
 ANTENNADIFFAREA                          0.218 LAYER ME3 ;
 ANTENNADIFFAREA                          0.218 LAYER ME4 ;
 ANTENNAMAXAREACAR                       13.984 LAYER ME1 ;
 ANTENNAMAXAREACAR                       16.784 LAYER ME2 ;
 ANTENNAMAXAREACAR                       19.584 LAYER ME3 ;
 ANTENNAMAXAREACAR                       22.384 LAYER ME4 ;
END DI42
PIN DO42
  DIRECTION OUTPUT ;
 PORT
  LAYER ME4 ;
  RECT 380.641 0.000 380.921 0.720 ;
  LAYER ME3 ;
  RECT 380.641 0.000 380.921 0.720 ;
  LAYER ME2 ;
  RECT 380.641 0.000 380.921 0.720 ;
  LAYER ME1 ;
  RECT 380.641 0.000 380.921 0.720 ;
 END
 ANTENNAPARTIALMETALAREA                  2.030 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME3 ;
 ANTENNADIFFAREA                          1.293 LAYER ME4 ;
END DO42
PIN DI41
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 374.611 0.000 374.891 0.720 ;
  LAYER ME3 ;
  RECT 374.611 0.000 374.891 0.720 ;
  LAYER ME2 ;
  RECT 374.611 0.000 374.891 0.720 ;
  LAYER ME1 ;
  RECT 374.611 0.000 374.891 0.720 ;
 END
 ANTENNAPARTIALMETALAREA                  0.805 LAYER ME1 ;
 ANTENNAGATEAREA                          0.072 LAYER ME1 ;
 ANTENNAGATEAREA                          0.072 LAYER ME2 ;
 ANTENNAGATEAREA                          0.072 LAYER ME3 ;
 ANTENNAGATEAREA                          0.072 LAYER ME4 ;
 ANTENNADIFFAREA                          0.218 LAYER ME1 ;
 ANTENNADIFFAREA                          0.218 LAYER ME2 ;
 ANTENNADIFFAREA                          0.218 LAYER ME3 ;
 ANTENNADIFFAREA                          0.218 LAYER ME4 ;
 ANTENNAMAXAREACAR                       13.984 LAYER ME1 ;
 ANTENNAMAXAREACAR                       16.784 LAYER ME2 ;
 ANTENNAMAXAREACAR                       19.584 LAYER ME3 ;
 ANTENNAMAXAREACAR                       22.384 LAYER ME4 ;
END DI41
PIN DO41
  DIRECTION OUTPUT ;
 PORT
  LAYER ME4 ;
  RECT 372.633 0.000 372.913 0.720 ;
  LAYER ME3 ;
  RECT 372.633 0.000 372.913 0.720 ;
  LAYER ME2 ;
  RECT 372.633 0.000 372.913 0.720 ;
  LAYER ME1 ;
  RECT 372.633 0.000 372.913 0.720 ;
 END
 ANTENNAPARTIALMETALAREA                  2.030 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME3 ;
 ANTENNADIFFAREA                          1.293 LAYER ME4 ;
END DO41
PIN DI40
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 366.603 0.000 366.883 0.720 ;
  LAYER ME3 ;
  RECT 366.603 0.000 366.883 0.720 ;
  LAYER ME2 ;
  RECT 366.603 0.000 366.883 0.720 ;
  LAYER ME1 ;
  RECT 366.603 0.000 366.883 0.720 ;
 END
 ANTENNAPARTIALMETALAREA                  0.805 LAYER ME1 ;
 ANTENNAGATEAREA                          0.072 LAYER ME1 ;
 ANTENNAGATEAREA                          0.072 LAYER ME2 ;
 ANTENNAGATEAREA                          0.072 LAYER ME3 ;
 ANTENNAGATEAREA                          0.072 LAYER ME4 ;
 ANTENNADIFFAREA                          0.218 LAYER ME1 ;
 ANTENNADIFFAREA                          0.218 LAYER ME2 ;
 ANTENNADIFFAREA                          0.218 LAYER ME3 ;
 ANTENNADIFFAREA                          0.218 LAYER ME4 ;
 ANTENNAMAXAREACAR                       13.984 LAYER ME1 ;
 ANTENNAMAXAREACAR                       16.784 LAYER ME2 ;
 ANTENNAMAXAREACAR                       19.584 LAYER ME3 ;
 ANTENNAMAXAREACAR                       22.384 LAYER ME4 ;
END DI40
PIN DO40
  DIRECTION OUTPUT ;
 PORT
  LAYER ME4 ;
  RECT 364.625 0.000 364.905 0.720 ;
  LAYER ME3 ;
  RECT 364.625 0.000 364.905 0.720 ;
  LAYER ME2 ;
  RECT 364.625 0.000 364.905 0.720 ;
  LAYER ME1 ;
  RECT 364.625 0.000 364.905 0.720 ;
 END
 ANTENNAPARTIALMETALAREA                  2.030 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME3 ;
 ANTENNADIFFAREA                          1.293 LAYER ME4 ;
END DO40
PIN DI39
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 358.595 0.000 358.875 0.720 ;
  LAYER ME3 ;
  RECT 358.595 0.000 358.875 0.720 ;
  LAYER ME2 ;
  RECT 358.595 0.000 358.875 0.720 ;
  LAYER ME1 ;
  RECT 358.595 0.000 358.875 0.720 ;
 END
 ANTENNAPARTIALMETALAREA                  0.805 LAYER ME1 ;
 ANTENNAGATEAREA                          0.072 LAYER ME1 ;
 ANTENNAGATEAREA                          0.072 LAYER ME2 ;
 ANTENNAGATEAREA                          0.072 LAYER ME3 ;
 ANTENNAGATEAREA                          0.072 LAYER ME4 ;
 ANTENNADIFFAREA                          0.218 LAYER ME1 ;
 ANTENNADIFFAREA                          0.218 LAYER ME2 ;
 ANTENNADIFFAREA                          0.218 LAYER ME3 ;
 ANTENNADIFFAREA                          0.218 LAYER ME4 ;
 ANTENNAMAXAREACAR                       13.984 LAYER ME1 ;
 ANTENNAMAXAREACAR                       16.784 LAYER ME2 ;
 ANTENNAMAXAREACAR                       19.584 LAYER ME3 ;
 ANTENNAMAXAREACAR                       22.384 LAYER ME4 ;
END DI39
PIN DO39
  DIRECTION OUTPUT ;
 PORT
  LAYER ME4 ;
  RECT 356.617 0.000 356.897 0.720 ;
  LAYER ME3 ;
  RECT 356.617 0.000 356.897 0.720 ;
  LAYER ME2 ;
  RECT 356.617 0.000 356.897 0.720 ;
  LAYER ME1 ;
  RECT 356.617 0.000 356.897 0.720 ;
 END
 ANTENNAPARTIALMETALAREA                  2.030 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME3 ;
 ANTENNADIFFAREA                          1.293 LAYER ME4 ;
END DO39
PIN DI38
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 350.587 0.000 350.867 0.720 ;
  LAYER ME3 ;
  RECT 350.587 0.000 350.867 0.720 ;
  LAYER ME2 ;
  RECT 350.587 0.000 350.867 0.720 ;
  LAYER ME1 ;
  RECT 350.587 0.000 350.867 0.720 ;
 END
 ANTENNAPARTIALMETALAREA                  0.805 LAYER ME1 ;
 ANTENNAGATEAREA                          0.072 LAYER ME1 ;
 ANTENNAGATEAREA                          0.072 LAYER ME2 ;
 ANTENNAGATEAREA                          0.072 LAYER ME3 ;
 ANTENNAGATEAREA                          0.072 LAYER ME4 ;
 ANTENNADIFFAREA                          0.218 LAYER ME1 ;
 ANTENNADIFFAREA                          0.218 LAYER ME2 ;
 ANTENNADIFFAREA                          0.218 LAYER ME3 ;
 ANTENNADIFFAREA                          0.218 LAYER ME4 ;
 ANTENNAMAXAREACAR                       13.984 LAYER ME1 ;
 ANTENNAMAXAREACAR                       16.784 LAYER ME2 ;
 ANTENNAMAXAREACAR                       19.584 LAYER ME3 ;
 ANTENNAMAXAREACAR                       22.384 LAYER ME4 ;
END DI38
PIN DO38
  DIRECTION OUTPUT ;
 PORT
  LAYER ME4 ;
  RECT 348.609 0.000 348.889 0.720 ;
  LAYER ME3 ;
  RECT 348.609 0.000 348.889 0.720 ;
  LAYER ME2 ;
  RECT 348.609 0.000 348.889 0.720 ;
  LAYER ME1 ;
  RECT 348.609 0.000 348.889 0.720 ;
 END
 ANTENNAPARTIALMETALAREA                  2.030 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME3 ;
 ANTENNADIFFAREA                          1.293 LAYER ME4 ;
END DO38
PIN DI37
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 342.579 0.000 342.859 0.720 ;
  LAYER ME3 ;
  RECT 342.579 0.000 342.859 0.720 ;
  LAYER ME2 ;
  RECT 342.579 0.000 342.859 0.720 ;
  LAYER ME1 ;
  RECT 342.579 0.000 342.859 0.720 ;
 END
 ANTENNAPARTIALMETALAREA                  0.805 LAYER ME1 ;
 ANTENNAGATEAREA                          0.072 LAYER ME1 ;
 ANTENNAGATEAREA                          0.072 LAYER ME2 ;
 ANTENNAGATEAREA                          0.072 LAYER ME3 ;
 ANTENNAGATEAREA                          0.072 LAYER ME4 ;
 ANTENNADIFFAREA                          0.218 LAYER ME1 ;
 ANTENNADIFFAREA                          0.218 LAYER ME2 ;
 ANTENNADIFFAREA                          0.218 LAYER ME3 ;
 ANTENNADIFFAREA                          0.218 LAYER ME4 ;
 ANTENNAMAXAREACAR                       13.984 LAYER ME1 ;
 ANTENNAMAXAREACAR                       16.784 LAYER ME2 ;
 ANTENNAMAXAREACAR                       19.584 LAYER ME3 ;
 ANTENNAMAXAREACAR                       22.384 LAYER ME4 ;
END DI37
PIN DO37
  DIRECTION OUTPUT ;
 PORT
  LAYER ME4 ;
  RECT 340.601 0.000 340.881 0.720 ;
  LAYER ME3 ;
  RECT 340.601 0.000 340.881 0.720 ;
  LAYER ME2 ;
  RECT 340.601 0.000 340.881 0.720 ;
  LAYER ME1 ;
  RECT 340.601 0.000 340.881 0.720 ;
 END
 ANTENNAPARTIALMETALAREA                  2.030 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME3 ;
 ANTENNADIFFAREA                          1.293 LAYER ME4 ;
END DO37
PIN DI36
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 334.571 0.000 334.851 0.720 ;
  LAYER ME3 ;
  RECT 334.571 0.000 334.851 0.720 ;
  LAYER ME2 ;
  RECT 334.571 0.000 334.851 0.720 ;
  LAYER ME1 ;
  RECT 334.571 0.000 334.851 0.720 ;
 END
 ANTENNAPARTIALMETALAREA                  0.522 LAYER ME1 ;
 ANTENNAGATEAREA                          0.072 LAYER ME1 ;
 ANTENNAGATEAREA                          0.072 LAYER ME2 ;
 ANTENNAGATEAREA                          0.072 LAYER ME3 ;
 ANTENNAGATEAREA                          0.072 LAYER ME4 ;
 ANTENNADIFFAREA                          0.218 LAYER ME1 ;
 ANTENNADIFFAREA                          0.218 LAYER ME2 ;
 ANTENNADIFFAREA                          0.218 LAYER ME3 ;
 ANTENNADIFFAREA                          0.218 LAYER ME4 ;
 ANTENNAMAXAREACAR                       10.048 LAYER ME1 ;
 ANTENNAMAXAREACAR                       12.848 LAYER ME2 ;
 ANTENNAMAXAREACAR                       15.648 LAYER ME3 ;
 ANTENNAMAXAREACAR                       18.448 LAYER ME4 ;
END DI36
PIN DO36
  DIRECTION OUTPUT ;
 PORT
  LAYER ME4 ;
  RECT 332.513 0.000 332.793 0.720 ;
  LAYER ME3 ;
  RECT 332.513 0.000 332.793 0.720 ;
  LAYER ME2 ;
  RECT 332.513 0.000 332.793 0.720 ;
  LAYER ME1 ;
  RECT 332.513 0.000 332.793 0.720 ;
 END
 ANTENNAPARTIALMETALAREA                  2.030 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME3 ;
 ANTENNADIFFAREA                          1.293 LAYER ME4 ;
END DO36
PIN WEB4
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 332.993 0.000 333.273 0.720 ;
  LAYER ME3 ;
  RECT 332.993 0.000 333.273 0.720 ;
  LAYER ME2 ;
  RECT 332.993 0.000 333.273 0.720 ;
  LAYER ME1 ;
  RECT 332.993 0.000 333.273 0.720 ;
 END
 ANTENNAPARTIALMETALAREA                  0.436 LAYER ME2 ;
 ANTENNAGATEAREA                          0.288 LAYER ME2 ;
 ANTENNAGATEAREA                          0.288 LAYER ME3 ;
 ANTENNAGATEAREA                          0.288 LAYER ME4 ;
 ANTENNADIFFAREA                          0.218 LAYER ME2 ;
 ANTENNADIFFAREA                          0.218 LAYER ME3 ;
 ANTENNADIFFAREA                          0.218 LAYER ME4 ;
 ANTENNAMAXAREACAR                        4.602 LAYER ME2 ;
 ANTENNAMAXAREACAR                        5.302 LAYER ME3 ;
 ANTENNAMAXAREACAR                        6.002 LAYER ME4 ;
END WEB4
OBS
  LAYER ME3 SPACING 0.260 ;
  RECT 0.000 0.000 620.075 98.967 ;
  LAYER ME2 SPACING 0.260 ;
  RECT 0.000 0.000 620.075 98.967 ;
  LAYER ME1 SPACING 0.260 ;
  RECT 0.000 0.000 620.075 98.967 ;
  LAYER ME4 SPACING 0.260 ;
  RECT 0.000 0.000 304.030 98.967 ;
  LAYER ME4 SPACING 0.260 ;
  RECT 305.684 0.000 306.804 98.967 ;
  LAYER ME4 SPACING 0.260 ;
  RECT 308.399 0.000 309.119 98.967 ;
  LAYER ME4 SPACING 0.260 ;
  RECT 309.849 0.000 310.569 98.967 ;
  LAYER ME4 SPACING 0.260 ;
  RECT 312.629 0.000 313.229 98.967 ;
  LAYER ME4 SPACING 0.260 ;
  RECT 315.843 0.000 317.529 98.967 ;
  LAYER ME4 SPACING 0.260 ;
  RECT 318.919 0.000 320.039 98.967 ;
  LAYER ME4 SPACING 0.260 ;
  RECT 321.314 0.000 322.034 98.967 ;
  LAYER ME4 SPACING 0.260 ;
  RECT 323.029 0.000 323.749 98.967 ;
  LAYER ME4 SPACING 0.260 ;
  RECT 324.949 0.000 620.075 98.967 ;
END
END SYKB110_256X9X8CM4
END LIBRARY





