# ________________________________________________________________________________________________
# 
# 
#             Synchronous One-Port Register File Compiler
# 
#                 UMC 0.11um LL AE Logic Process
# 
# ________________________________________________________________________________________________
# 
#               
#         Copyright (C) 2024 Faraday Technology Corporation. All Rights Reserved.       
#                
#         This source code is an unpublished work belongs to Faraday Technology Corporation       
#         It is considered a trade secret and is not to be divulged or       
#         used by parties who have not received written authorization from       
#         Faraday Technology Corporation       
#                
#         Faraday's home page can be found at: http://www.faraday-tech.com/       
#                
# ________________________________________________________________________________________________
# 
#        IP Name            :  FSR0K_B_SY                
#        IP Version         :  1.4.0                     
#        IP Release Status  :  Active                    
#        Word               :  64                        
#        Bit                :  12                        
#        Byte               :  8                         
#        Mux                :  2                         
#        Output Loading     :  0.01                      
#        Clock Input Slew   :  0.016                     
#        Data Input Slew    :  0.016                     
#        Ring Type          :  Ringless Model            
#        Ring Width         :  0                         
#        Bus Format         :  0                         
#        Memaker Path       :  /home/mem/Desktop/memlib  
#        GUI Version        :  m20230904                 
#        Date               :  2024/09/07 14:44:15       
# ________________________________________________________________________________________________
# 

VERSION 5.5 ;
NAMESCASESENSITIVE ON ;
MACRO SYKB110_64X12X8CM2
CLASS BLOCK ;
FOREIGN SYKB110_64X12X8CM2 0.000 0.000 ;
ORIGIN 0.000 0.000 ;
SIZE 427.883 BY 80.703 ;
SYMMETRY x y r90 ;
SITE core ;
PIN GND
  DIRECTION INOUT ;
  USE GROUND ;
 PORT
  LAYER ME4 ;
  RECT 236.614 1.781 236.954 80.703 ;
 END
 PORT
  LAYER ME4 ;
  RECT 232.610 1.781 232.950 80.703 ;
 END
 PORT
  LAYER ME4 ;
  RECT 234.612 1.781 234.952 80.703 ;
 END
 PORT
  LAYER ME4 ;
  RECT 235.423 0.000 236.143 44.094 ;
 END
 PORT
  LAYER ME4 ;
  RECT 240.618 1.781 240.958 80.703 ;
 END
 PORT
  LAYER ME4 ;
  RECT 238.616 1.781 238.956 80.703 ;
 END
 PORT
  LAYER ME4 ;
  RECT 239.427 0.000 240.147 44.094 ;
 END
 PORT
  LAYER ME4 ;
  RECT 244.622 1.781 244.962 80.703 ;
 END
 PORT
  LAYER ME4 ;
  RECT 242.620 1.781 242.960 80.703 ;
 END
 PORT
  LAYER ME4 ;
  RECT 243.431 0.000 244.151 44.094 ;
 END
 PORT
  LAYER ME4 ;
  RECT 248.626 1.781 248.966 80.703 ;
 END
 PORT
  LAYER ME4 ;
  RECT 246.624 1.781 246.964 80.703 ;
 END
 PORT
  LAYER ME4 ;
  RECT 247.435 0.000 248.155 44.094 ;
 END
 PORT
  LAYER ME4 ;
  RECT 252.630 1.781 252.970 80.703 ;
 END
 PORT
  LAYER ME4 ;
  RECT 250.628 1.781 250.968 80.703 ;
 END
 PORT
  LAYER ME4 ;
  RECT 251.439 0.000 252.159 44.094 ;
 END
 PORT
  LAYER ME4 ;
  RECT 256.634 1.781 256.974 80.703 ;
 END
 PORT
  LAYER ME4 ;
  RECT 254.632 1.781 254.972 80.703 ;
 END
 PORT
  LAYER ME4 ;
  RECT 255.443 0.000 256.163 44.094 ;
 END
 PORT
  LAYER ME4 ;
  RECT 260.638 1.781 260.978 80.703 ;
 END
 PORT
  LAYER ME4 ;
  RECT 258.636 1.781 258.976 80.703 ;
 END
 PORT
  LAYER ME4 ;
  RECT 259.447 0.000 260.167 44.094 ;
 END
 PORT
  LAYER ME4 ;
  RECT 264.642 1.781 264.982 80.703 ;
 END
 PORT
  LAYER ME4 ;
  RECT 262.640 1.781 262.980 80.703 ;
 END
 PORT
  LAYER ME4 ;
  RECT 263.451 0.000 264.171 44.094 ;
 END
 PORT
  LAYER ME4 ;
  RECT 268.646 1.781 268.986 80.703 ;
 END
 PORT
  LAYER ME4 ;
  RECT 266.644 1.781 266.984 80.703 ;
 END
 PORT
  LAYER ME4 ;
  RECT 267.455 0.000 268.175 44.094 ;
 END
 PORT
  LAYER ME4 ;
  RECT 272.650 1.781 272.990 80.703 ;
 END
 PORT
  LAYER ME4 ;
  RECT 270.648 1.781 270.988 80.703 ;
 END
 PORT
  LAYER ME4 ;
  RECT 271.459 0.000 272.179 44.094 ;
 END
 PORT
  LAYER ME4 ;
  RECT 276.654 1.781 276.994 80.703 ;
 END
 PORT
  LAYER ME4 ;
  RECT 274.652 1.781 274.992 80.703 ;
 END
 PORT
  LAYER ME4 ;
  RECT 275.463 0.000 276.183 44.094 ;
 END
 PORT
  LAYER ME4 ;
  RECT 280.658 1.781 280.998 80.703 ;
 END
 PORT
  LAYER ME4 ;
  RECT 278.656 1.781 278.996 80.703 ;
 END
 PORT
  LAYER ME4 ;
  RECT 279.467 0.000 280.187 44.094 ;
 END
 PORT
  LAYER ME4 ;
  RECT 284.662 1.781 285.002 80.703 ;
 END
 PORT
  LAYER ME4 ;
  RECT 282.660 1.781 283.000 80.703 ;
 END
 PORT
  LAYER ME4 ;
  RECT 283.471 0.000 284.191 44.094 ;
 END
 PORT
  LAYER ME4 ;
  RECT 288.666 1.781 289.006 80.703 ;
 END
 PORT
  LAYER ME4 ;
  RECT 286.664 1.781 287.004 80.703 ;
 END
 PORT
  LAYER ME4 ;
  RECT 287.475 0.000 288.195 44.094 ;
 END
 PORT
  LAYER ME4 ;
  RECT 292.670 1.781 293.010 80.703 ;
 END
 PORT
  LAYER ME4 ;
  RECT 290.668 1.781 291.008 80.703 ;
 END
 PORT
  LAYER ME4 ;
  RECT 291.479 0.000 292.199 44.094 ;
 END
 PORT
  LAYER ME4 ;
  RECT 296.674 1.781 297.014 80.703 ;
 END
 PORT
  LAYER ME4 ;
  RECT 294.672 1.781 295.012 80.703 ;
 END
 PORT
  LAYER ME4 ;
  RECT 295.483 0.000 296.203 44.094 ;
 END
 PORT
  LAYER ME4 ;
  RECT 300.678 1.781 301.018 80.703 ;
 END
 PORT
  LAYER ME4 ;
  RECT 298.676 1.781 299.016 80.703 ;
 END
 PORT
  LAYER ME4 ;
  RECT 299.487 0.000 300.207 44.094 ;
 END
 PORT
  LAYER ME4 ;
  RECT 304.682 1.781 305.022 80.703 ;
 END
 PORT
  LAYER ME4 ;
  RECT 302.680 1.781 303.020 80.703 ;
 END
 PORT
  LAYER ME4 ;
  RECT 303.491 0.000 304.211 44.094 ;
 END
 PORT
  LAYER ME4 ;
  RECT 308.686 1.781 309.026 80.703 ;
 END
 PORT
  LAYER ME4 ;
  RECT 306.684 1.781 307.024 80.703 ;
 END
 PORT
  LAYER ME4 ;
  RECT 307.495 0.000 308.215 44.094 ;
 END
 PORT
  LAYER ME4 ;
  RECT 312.690 1.781 313.030 80.703 ;
 END
 PORT
  LAYER ME4 ;
  RECT 310.688 1.781 311.028 80.703 ;
 END
 PORT
  LAYER ME4 ;
  RECT 311.499 0.000 312.219 44.094 ;
 END
 PORT
  LAYER ME4 ;
  RECT 316.694 1.781 317.034 80.703 ;
 END
 PORT
  LAYER ME4 ;
  RECT 314.692 1.781 315.032 80.703 ;
 END
 PORT
  LAYER ME4 ;
  RECT 315.503 0.000 316.223 44.094 ;
 END
 PORT
  LAYER ME4 ;
  RECT 320.698 1.781 321.038 80.703 ;
 END
 PORT
  LAYER ME4 ;
  RECT 318.696 1.781 319.036 80.703 ;
 END
 PORT
  LAYER ME4 ;
  RECT 319.507 0.000 320.227 44.094 ;
 END
 PORT
  LAYER ME4 ;
  RECT 324.702 1.781 325.042 80.703 ;
 END
 PORT
  LAYER ME4 ;
  RECT 322.700 1.781 323.040 80.703 ;
 END
 PORT
  LAYER ME4 ;
  RECT 323.511 0.000 324.231 44.094 ;
 END
 PORT
  LAYER ME4 ;
  RECT 328.706 1.781 329.046 80.703 ;
 END
 PORT
  LAYER ME4 ;
  RECT 326.704 1.781 327.044 80.703 ;
 END
 PORT
  LAYER ME4 ;
  RECT 327.515 0.000 328.235 44.094 ;
 END
 PORT
  LAYER ME4 ;
  RECT 332.710 1.781 333.050 80.703 ;
 END
 PORT
  LAYER ME4 ;
  RECT 330.708 1.781 331.048 80.703 ;
 END
 PORT
  LAYER ME4 ;
  RECT 331.519 0.000 332.239 44.094 ;
 END
 PORT
  LAYER ME4 ;
  RECT 336.714 1.781 337.054 80.703 ;
 END
 PORT
  LAYER ME4 ;
  RECT 334.712 1.781 335.052 80.703 ;
 END
 PORT
  LAYER ME4 ;
  RECT 335.523 0.000 336.243 44.094 ;
 END
 PORT
  LAYER ME4 ;
  RECT 340.718 1.781 341.058 80.703 ;
 END
 PORT
  LAYER ME4 ;
  RECT 338.716 1.781 339.056 80.703 ;
 END
 PORT
  LAYER ME4 ;
  RECT 339.527 0.000 340.247 44.094 ;
 END
 PORT
  LAYER ME4 ;
  RECT 344.722 1.781 345.062 80.703 ;
 END
 PORT
  LAYER ME4 ;
  RECT 342.720 1.781 343.060 80.703 ;
 END
 PORT
  LAYER ME4 ;
  RECT 343.531 0.000 344.251 44.094 ;
 END
 PORT
  LAYER ME4 ;
  RECT 348.726 1.781 349.066 80.703 ;
 END
 PORT
  LAYER ME4 ;
  RECT 346.724 1.781 347.064 80.703 ;
 END
 PORT
  LAYER ME4 ;
  RECT 347.535 0.000 348.255 44.094 ;
 END
 PORT
  LAYER ME4 ;
  RECT 352.730 1.781 353.070 80.703 ;
 END
 PORT
  LAYER ME4 ;
  RECT 350.728 1.781 351.068 80.703 ;
 END
 PORT
  LAYER ME4 ;
  RECT 351.539 0.000 352.259 44.094 ;
 END
 PORT
  LAYER ME4 ;
  RECT 356.734 1.781 357.074 80.703 ;
 END
 PORT
  LAYER ME4 ;
  RECT 354.732 1.781 355.072 80.703 ;
 END
 PORT
  LAYER ME4 ;
  RECT 355.543 0.000 356.263 44.094 ;
 END
 PORT
  LAYER ME4 ;
  RECT 360.738 1.781 361.078 80.703 ;
 END
 PORT
  LAYER ME4 ;
  RECT 358.736 1.781 359.076 80.703 ;
 END
 PORT
  LAYER ME4 ;
  RECT 359.547 0.000 360.267 44.094 ;
 END
 PORT
  LAYER ME4 ;
  RECT 364.742 1.781 365.082 80.703 ;
 END
 PORT
  LAYER ME4 ;
  RECT 362.740 1.781 363.080 80.703 ;
 END
 PORT
  LAYER ME4 ;
  RECT 363.551 0.000 364.271 44.094 ;
 END
 PORT
  LAYER ME4 ;
  RECT 368.746 1.781 369.086 80.703 ;
 END
 PORT
  LAYER ME4 ;
  RECT 366.744 1.781 367.084 80.703 ;
 END
 PORT
  LAYER ME4 ;
  RECT 367.555 0.000 368.275 44.094 ;
 END
 PORT
  LAYER ME4 ;
  RECT 372.750 1.781 373.090 80.703 ;
 END
 PORT
  LAYER ME4 ;
  RECT 370.748 1.781 371.088 80.703 ;
 END
 PORT
  LAYER ME4 ;
  RECT 371.559 0.000 372.279 44.094 ;
 END
 PORT
  LAYER ME4 ;
  RECT 376.754 1.781 377.094 80.703 ;
 END
 PORT
  LAYER ME4 ;
  RECT 374.752 1.781 375.092 80.703 ;
 END
 PORT
  LAYER ME4 ;
  RECT 375.563 0.000 376.283 44.094 ;
 END
 PORT
  LAYER ME4 ;
  RECT 380.758 1.781 381.098 80.703 ;
 END
 PORT
  LAYER ME4 ;
  RECT 378.756 1.781 379.096 80.703 ;
 END
 PORT
  LAYER ME4 ;
  RECT 379.567 0.000 380.287 44.094 ;
 END
 PORT
  LAYER ME4 ;
  RECT 384.762 1.781 385.102 80.703 ;
 END
 PORT
  LAYER ME4 ;
  RECT 382.760 1.781 383.100 80.703 ;
 END
 PORT
  LAYER ME4 ;
  RECT 383.571 0.000 384.291 44.094 ;
 END
 PORT
  LAYER ME4 ;
  RECT 388.766 1.781 389.106 80.703 ;
 END
 PORT
  LAYER ME4 ;
  RECT 386.764 1.781 387.104 80.703 ;
 END
 PORT
  LAYER ME4 ;
  RECT 387.575 0.000 388.295 44.094 ;
 END
 PORT
  LAYER ME4 ;
  RECT 392.770 1.781 393.110 80.703 ;
 END
 PORT
  LAYER ME4 ;
  RECT 390.768 1.781 391.108 80.703 ;
 END
 PORT
  LAYER ME4 ;
  RECT 391.579 0.000 392.299 44.094 ;
 END
 PORT
  LAYER ME4 ;
  RECT 396.774 1.781 397.114 80.703 ;
 END
 PORT
  LAYER ME4 ;
  RECT 394.772 1.781 395.112 80.703 ;
 END
 PORT
  LAYER ME4 ;
  RECT 395.583 0.000 396.303 44.094 ;
 END
 PORT
  LAYER ME4 ;
  RECT 400.778 1.781 401.118 80.703 ;
 END
 PORT
  LAYER ME4 ;
  RECT 398.776 1.781 399.116 80.703 ;
 END
 PORT
  LAYER ME4 ;
  RECT 399.587 0.000 400.307 44.094 ;
 END
 PORT
  LAYER ME4 ;
  RECT 404.782 1.781 405.122 80.703 ;
 END
 PORT
  LAYER ME4 ;
  RECT 402.780 1.781 403.120 80.703 ;
 END
 PORT
  LAYER ME4 ;
  RECT 403.591 0.000 404.311 44.094 ;
 END
 PORT
  LAYER ME4 ;
  RECT 408.786 1.781 409.126 80.703 ;
 END
 PORT
  LAYER ME4 ;
  RECT 406.784 1.781 407.124 80.703 ;
 END
 PORT
  LAYER ME4 ;
  RECT 407.595 0.000 408.315 44.094 ;
 END
 PORT
  LAYER ME4 ;
  RECT 412.790 1.781 413.130 80.703 ;
 END
 PORT
  LAYER ME4 ;
  RECT 410.788 1.781 411.128 80.703 ;
 END
 PORT
  LAYER ME4 ;
  RECT 411.599 0.000 412.319 44.094 ;
 END
 PORT
  LAYER ME4 ;
  RECT 416.794 1.781 417.134 80.703 ;
 END
 PORT
  LAYER ME4 ;
  RECT 414.792 1.781 415.132 80.703 ;
 END
 PORT
  LAYER ME4 ;
  RECT 415.603 0.000 416.323 44.094 ;
 END
 PORT
  LAYER ME4 ;
  RECT 420.798 1.781 421.138 80.703 ;
 END
 PORT
  LAYER ME4 ;
  RECT 418.796 1.781 419.136 80.703 ;
 END
 PORT
  LAYER ME4 ;
  RECT 419.607 0.000 420.327 44.094 ;
 END
 PORT
  LAYER ME4 ;
  RECT 424.802 1.781 425.142 80.703 ;
 END
 PORT
  LAYER ME4 ;
  RECT 422.800 1.781 423.140 80.703 ;
 END
 PORT
  LAYER ME4 ;
  RECT 423.611 0.000 424.331 44.094 ;
 END
 PORT
  LAYER ME4 ;
  RECT 425.803 0.000 426.143 80.703 ;
 END
 PORT
  LAYER ME4 ;
  RECT 213.753 0.000 214.473 80.703 ;
 END
 PORT
  LAYER ME4 ;
  RECT 219.747 0.000 220.467 80.703 ;
 END
 PORT
  LAYER ME4 ;
  RECT 225.218 0.000 225.938 80.703 ;
 END
 PORT
  LAYER ME4 ;
  RECT 226.933 0.000 227.653 80.703 ;
 END
 PORT
  LAYER ME4 ;
  RECT 229.929 0.000 230.529 80.703 ;
 END
 PORT
  LAYER ME4 ;
  RECT 231.609 1.781 231.949 80.703 ;
 END
 PORT
  LAYER ME4 ;
  RECT 206.194 0.000 206.914 80.703 ;
 END
 PORT
  LAYER ME4 ;
  RECT 204.154 1.781 204.874 79.944 ;
 END
 PORT
  LAYER ME4 ;
  RECT 202.034 0.000 202.754 80.703 ;
 END
 PORT
  LAYER ME4 ;
  RECT 199.994 1.781 200.714 80.703 ;
 END
 PORT
  LAYER ME4 ;
  RECT 1.740 0.000 2.080 80.703 ;
 END
 PORT
  LAYER ME4 ;
  RECT 6.745 1.781 7.085 80.703 ;
 END
 PORT
  LAYER ME4 ;
  RECT 2.741 1.781 3.081 80.703 ;
 END
 PORT
  LAYER ME4 ;
  RECT 4.743 1.781 5.083 80.703 ;
 END
 PORT
  LAYER ME4 ;
  RECT 5.554 0.000 6.274 44.094 ;
 END
 PORT
  LAYER ME4 ;
  RECT 10.749 1.781 11.089 80.703 ;
 END
 PORT
  LAYER ME4 ;
  RECT 8.747 1.781 9.087 80.703 ;
 END
 PORT
  LAYER ME4 ;
  RECT 9.558 0.000 10.278 44.094 ;
 END
 PORT
  LAYER ME4 ;
  RECT 14.753 1.781 15.093 80.703 ;
 END
 PORT
  LAYER ME4 ;
  RECT 12.751 1.781 13.091 80.703 ;
 END
 PORT
  LAYER ME4 ;
  RECT 13.562 0.000 14.282 44.094 ;
 END
 PORT
  LAYER ME4 ;
  RECT 18.757 1.781 19.097 80.703 ;
 END
 PORT
  LAYER ME4 ;
  RECT 16.755 1.781 17.095 80.703 ;
 END
 PORT
  LAYER ME4 ;
  RECT 17.566 0.000 18.286 44.094 ;
 END
 PORT
  LAYER ME4 ;
  RECT 22.761 1.781 23.101 80.703 ;
 END
 PORT
  LAYER ME4 ;
  RECT 20.759 1.781 21.099 80.703 ;
 END
 PORT
  LAYER ME4 ;
  RECT 21.570 0.000 22.290 44.094 ;
 END
 PORT
  LAYER ME4 ;
  RECT 26.765 1.781 27.105 80.703 ;
 END
 PORT
  LAYER ME4 ;
  RECT 24.763 1.781 25.103 80.703 ;
 END
 PORT
  LAYER ME4 ;
  RECT 25.574 0.000 26.294 44.094 ;
 END
 PORT
  LAYER ME4 ;
  RECT 30.769 1.781 31.109 80.703 ;
 END
 PORT
  LAYER ME4 ;
  RECT 28.767 1.781 29.107 80.703 ;
 END
 PORT
  LAYER ME4 ;
  RECT 29.578 0.000 30.298 44.094 ;
 END
 PORT
  LAYER ME4 ;
  RECT 34.773 1.781 35.113 80.703 ;
 END
 PORT
  LAYER ME4 ;
  RECT 32.771 1.781 33.111 80.703 ;
 END
 PORT
  LAYER ME4 ;
  RECT 33.582 0.000 34.302 44.094 ;
 END
 PORT
  LAYER ME4 ;
  RECT 38.777 1.781 39.117 80.703 ;
 END
 PORT
  LAYER ME4 ;
  RECT 36.775 1.781 37.115 80.703 ;
 END
 PORT
  LAYER ME4 ;
  RECT 37.586 0.000 38.306 44.094 ;
 END
 PORT
  LAYER ME4 ;
  RECT 42.781 1.781 43.121 80.703 ;
 END
 PORT
  LAYER ME4 ;
  RECT 40.779 1.781 41.119 80.703 ;
 END
 PORT
  LAYER ME4 ;
  RECT 41.590 0.000 42.310 44.094 ;
 END
 PORT
  LAYER ME4 ;
  RECT 46.785 1.781 47.125 80.703 ;
 END
 PORT
  LAYER ME4 ;
  RECT 44.783 1.781 45.123 80.703 ;
 END
 PORT
  LAYER ME4 ;
  RECT 45.594 0.000 46.314 44.094 ;
 END
 PORT
  LAYER ME4 ;
  RECT 50.789 1.781 51.129 80.703 ;
 END
 PORT
  LAYER ME4 ;
  RECT 48.787 1.781 49.127 80.703 ;
 END
 PORT
  LAYER ME4 ;
  RECT 49.598 0.000 50.318 44.094 ;
 END
 PORT
  LAYER ME4 ;
  RECT 54.793 1.781 55.133 80.703 ;
 END
 PORT
  LAYER ME4 ;
  RECT 52.791 1.781 53.131 80.703 ;
 END
 PORT
  LAYER ME4 ;
  RECT 53.602 0.000 54.322 44.094 ;
 END
 PORT
  LAYER ME4 ;
  RECT 58.797 1.781 59.137 80.703 ;
 END
 PORT
  LAYER ME4 ;
  RECT 56.795 1.781 57.135 80.703 ;
 END
 PORT
  LAYER ME4 ;
  RECT 57.606 0.000 58.326 44.094 ;
 END
 PORT
  LAYER ME4 ;
  RECT 62.801 1.781 63.141 80.703 ;
 END
 PORT
  LAYER ME4 ;
  RECT 60.799 1.781 61.139 80.703 ;
 END
 PORT
  LAYER ME4 ;
  RECT 61.610 0.000 62.330 44.094 ;
 END
 PORT
  LAYER ME4 ;
  RECT 66.805 1.781 67.145 80.703 ;
 END
 PORT
  LAYER ME4 ;
  RECT 64.803 1.781 65.143 80.703 ;
 END
 PORT
  LAYER ME4 ;
  RECT 65.614 0.000 66.334 44.094 ;
 END
 PORT
  LAYER ME4 ;
  RECT 70.809 1.781 71.149 80.703 ;
 END
 PORT
  LAYER ME4 ;
  RECT 68.807 1.781 69.147 80.703 ;
 END
 PORT
  LAYER ME4 ;
  RECT 69.618 0.000 70.338 44.094 ;
 END
 PORT
  LAYER ME4 ;
  RECT 74.813 1.781 75.153 80.703 ;
 END
 PORT
  LAYER ME4 ;
  RECT 72.811 1.781 73.151 80.703 ;
 END
 PORT
  LAYER ME4 ;
  RECT 73.622 0.000 74.342 44.094 ;
 END
 PORT
  LAYER ME4 ;
  RECT 78.817 1.781 79.157 80.703 ;
 END
 PORT
  LAYER ME4 ;
  RECT 76.815 1.781 77.155 80.703 ;
 END
 PORT
  LAYER ME4 ;
  RECT 77.626 0.000 78.346 44.094 ;
 END
 PORT
  LAYER ME4 ;
  RECT 82.821 1.781 83.161 80.703 ;
 END
 PORT
  LAYER ME4 ;
  RECT 80.819 1.781 81.159 80.703 ;
 END
 PORT
  LAYER ME4 ;
  RECT 81.630 0.000 82.350 44.094 ;
 END
 PORT
  LAYER ME4 ;
  RECT 86.825 1.781 87.165 80.703 ;
 END
 PORT
  LAYER ME4 ;
  RECT 84.823 1.781 85.163 80.703 ;
 END
 PORT
  LAYER ME4 ;
  RECT 85.634 0.000 86.354 44.094 ;
 END
 PORT
  LAYER ME4 ;
  RECT 90.829 1.781 91.169 80.703 ;
 END
 PORT
  LAYER ME4 ;
  RECT 88.827 1.781 89.167 80.703 ;
 END
 PORT
  LAYER ME4 ;
  RECT 89.638 0.000 90.358 44.094 ;
 END
 PORT
  LAYER ME4 ;
  RECT 94.833 1.781 95.173 80.703 ;
 END
 PORT
  LAYER ME4 ;
  RECT 92.831 1.781 93.171 80.703 ;
 END
 PORT
  LAYER ME4 ;
  RECT 93.642 0.000 94.362 44.094 ;
 END
 PORT
  LAYER ME4 ;
  RECT 98.837 1.781 99.177 80.703 ;
 END
 PORT
  LAYER ME4 ;
  RECT 96.835 1.781 97.175 80.703 ;
 END
 PORT
  LAYER ME4 ;
  RECT 97.646 0.000 98.366 44.094 ;
 END
 PORT
  LAYER ME4 ;
  RECT 102.841 1.781 103.181 80.703 ;
 END
 PORT
  LAYER ME4 ;
  RECT 100.839 1.781 101.179 80.703 ;
 END
 PORT
  LAYER ME4 ;
  RECT 101.650 0.000 102.370 44.094 ;
 END
 PORT
  LAYER ME4 ;
  RECT 106.845 1.781 107.185 80.703 ;
 END
 PORT
  LAYER ME4 ;
  RECT 104.843 1.781 105.183 80.703 ;
 END
 PORT
  LAYER ME4 ;
  RECT 105.654 0.000 106.374 44.094 ;
 END
 PORT
  LAYER ME4 ;
  RECT 110.849 1.781 111.189 80.703 ;
 END
 PORT
  LAYER ME4 ;
  RECT 108.847 1.781 109.187 80.703 ;
 END
 PORT
  LAYER ME4 ;
  RECT 109.658 0.000 110.378 44.094 ;
 END
 PORT
  LAYER ME4 ;
  RECT 114.853 1.781 115.193 80.703 ;
 END
 PORT
  LAYER ME4 ;
  RECT 112.851 1.781 113.191 80.703 ;
 END
 PORT
  LAYER ME4 ;
  RECT 113.662 0.000 114.382 44.094 ;
 END
 PORT
  LAYER ME4 ;
  RECT 118.857 1.781 119.197 80.703 ;
 END
 PORT
  LAYER ME4 ;
  RECT 116.855 1.781 117.195 80.703 ;
 END
 PORT
  LAYER ME4 ;
  RECT 117.666 0.000 118.386 44.094 ;
 END
 PORT
  LAYER ME4 ;
  RECT 122.861 1.781 123.201 80.703 ;
 END
 PORT
  LAYER ME4 ;
  RECT 120.859 1.781 121.199 80.703 ;
 END
 PORT
  LAYER ME4 ;
  RECT 121.670 0.000 122.390 44.094 ;
 END
 PORT
  LAYER ME4 ;
  RECT 126.865 1.781 127.205 80.703 ;
 END
 PORT
  LAYER ME4 ;
  RECT 124.863 1.781 125.203 80.703 ;
 END
 PORT
  LAYER ME4 ;
  RECT 125.674 0.000 126.394 44.094 ;
 END
 PORT
  LAYER ME4 ;
  RECT 130.869 1.781 131.209 80.703 ;
 END
 PORT
  LAYER ME4 ;
  RECT 128.867 1.781 129.207 80.703 ;
 END
 PORT
  LAYER ME4 ;
  RECT 129.678 0.000 130.398 44.094 ;
 END
 PORT
  LAYER ME4 ;
  RECT 134.873 1.781 135.213 80.703 ;
 END
 PORT
  LAYER ME4 ;
  RECT 132.871 1.781 133.211 80.703 ;
 END
 PORT
  LAYER ME4 ;
  RECT 133.682 0.000 134.402 44.094 ;
 END
 PORT
  LAYER ME4 ;
  RECT 138.877 1.781 139.217 80.703 ;
 END
 PORT
  LAYER ME4 ;
  RECT 136.875 1.781 137.215 80.703 ;
 END
 PORT
  LAYER ME4 ;
  RECT 137.686 0.000 138.406 44.094 ;
 END
 PORT
  LAYER ME4 ;
  RECT 142.881 1.781 143.221 80.703 ;
 END
 PORT
  LAYER ME4 ;
  RECT 140.879 1.781 141.219 80.703 ;
 END
 PORT
  LAYER ME4 ;
  RECT 141.690 0.000 142.410 44.094 ;
 END
 PORT
  LAYER ME4 ;
  RECT 146.885 1.781 147.225 80.703 ;
 END
 PORT
  LAYER ME4 ;
  RECT 144.883 1.781 145.223 80.703 ;
 END
 PORT
  LAYER ME4 ;
  RECT 145.694 0.000 146.414 44.094 ;
 END
 PORT
  LAYER ME4 ;
  RECT 150.889 1.781 151.229 80.703 ;
 END
 PORT
  LAYER ME4 ;
  RECT 148.887 1.781 149.227 80.703 ;
 END
 PORT
  LAYER ME4 ;
  RECT 149.698 0.000 150.418 44.094 ;
 END
 PORT
  LAYER ME4 ;
  RECT 154.893 1.781 155.233 80.703 ;
 END
 PORT
  LAYER ME4 ;
  RECT 152.891 1.781 153.231 80.703 ;
 END
 PORT
  LAYER ME4 ;
  RECT 153.702 0.000 154.422 44.094 ;
 END
 PORT
  LAYER ME4 ;
  RECT 158.897 1.781 159.237 80.703 ;
 END
 PORT
  LAYER ME4 ;
  RECT 156.895 1.781 157.235 80.703 ;
 END
 PORT
  LAYER ME4 ;
  RECT 157.706 0.000 158.426 44.094 ;
 END
 PORT
  LAYER ME4 ;
  RECT 162.901 1.781 163.241 80.703 ;
 END
 PORT
  LAYER ME4 ;
  RECT 160.899 1.781 161.239 80.703 ;
 END
 PORT
  LAYER ME4 ;
  RECT 161.710 0.000 162.430 44.094 ;
 END
 PORT
  LAYER ME4 ;
  RECT 166.905 1.781 167.245 80.703 ;
 END
 PORT
  LAYER ME4 ;
  RECT 164.903 1.781 165.243 80.703 ;
 END
 PORT
  LAYER ME4 ;
  RECT 165.714 0.000 166.434 44.094 ;
 END
 PORT
  LAYER ME4 ;
  RECT 170.909 1.781 171.249 80.703 ;
 END
 PORT
  LAYER ME4 ;
  RECT 168.907 1.781 169.247 80.703 ;
 END
 PORT
  LAYER ME4 ;
  RECT 169.718 0.000 170.438 44.094 ;
 END
 PORT
  LAYER ME4 ;
  RECT 174.913 1.781 175.253 80.703 ;
 END
 PORT
  LAYER ME4 ;
  RECT 172.911 1.781 173.251 80.703 ;
 END
 PORT
  LAYER ME4 ;
  RECT 173.722 0.000 174.442 44.094 ;
 END
 PORT
  LAYER ME4 ;
  RECT 178.917 1.781 179.257 80.703 ;
 END
 PORT
  LAYER ME4 ;
  RECT 176.915 1.781 177.255 80.703 ;
 END
 PORT
  LAYER ME4 ;
  RECT 177.726 0.000 178.446 44.094 ;
 END
 PORT
  LAYER ME4 ;
  RECT 182.921 1.781 183.261 80.703 ;
 END
 PORT
  LAYER ME4 ;
  RECT 180.919 1.781 181.259 80.703 ;
 END
 PORT
  LAYER ME4 ;
  RECT 181.730 0.000 182.450 44.094 ;
 END
 PORT
  LAYER ME4 ;
  RECT 186.925 1.781 187.265 80.703 ;
 END
 PORT
  LAYER ME4 ;
  RECT 184.923 1.781 185.263 80.703 ;
 END
 PORT
  LAYER ME4 ;
  RECT 185.734 0.000 186.454 44.094 ;
 END
 PORT
  LAYER ME4 ;
  RECT 190.929 1.781 191.269 80.703 ;
 END
 PORT
  LAYER ME4 ;
  RECT 188.927 1.781 189.267 80.703 ;
 END
 PORT
  LAYER ME4 ;
  RECT 189.738 0.000 190.458 44.094 ;
 END
 PORT
  LAYER ME4 ;
  RECT 194.933 1.781 195.273 80.703 ;
 END
 PORT
  LAYER ME4 ;
  RECT 192.931 1.781 193.271 80.703 ;
 END
 PORT
  LAYER ME4 ;
  RECT 193.742 0.000 194.462 44.094 ;
 END
 PORT
  LAYER ME4 ;
  RECT 197.874 0.000 198.594 80.703 ;
 END
 PORT
  LAYER ME4 ;
  RECT 195.934 0.000 196.274 80.703 ;
 END
END GND
PIN VCC
  DIRECTION INOUT ;
  USE POWER ;
 PORT
  LAYER ME4 ;
  RECT 235.613 45.394 235.953 80.703 ;
 END
 PORT
  LAYER ME4 ;
  RECT 233.421 0.000 234.141 46.394 ;
 END
 PORT
  LAYER ME4 ;
  RECT 239.617 45.394 239.957 80.703 ;
 END
 PORT
  LAYER ME4 ;
  RECT 237.425 0.000 238.145 46.394 ;
 END
 PORT
  LAYER ME4 ;
  RECT 243.621 45.394 243.961 80.703 ;
 END
 PORT
  LAYER ME4 ;
  RECT 241.429 0.000 242.149 46.394 ;
 END
 PORT
  LAYER ME4 ;
  RECT 247.625 45.394 247.965 80.703 ;
 END
 PORT
  LAYER ME4 ;
  RECT 245.433 0.000 246.153 46.394 ;
 END
 PORT
  LAYER ME4 ;
  RECT 251.629 45.394 251.969 80.703 ;
 END
 PORT
  LAYER ME4 ;
  RECT 249.437 0.000 250.157 46.394 ;
 END
 PORT
  LAYER ME4 ;
  RECT 255.633 45.394 255.973 80.703 ;
 END
 PORT
  LAYER ME4 ;
  RECT 253.441 0.000 254.161 46.394 ;
 END
 PORT
  LAYER ME4 ;
  RECT 259.637 45.394 259.977 80.703 ;
 END
 PORT
  LAYER ME4 ;
  RECT 257.445 0.000 258.165 46.394 ;
 END
 PORT
  LAYER ME4 ;
  RECT 263.641 45.394 263.981 80.703 ;
 END
 PORT
  LAYER ME4 ;
  RECT 261.449 0.000 262.169 46.394 ;
 END
 PORT
  LAYER ME4 ;
  RECT 267.645 45.394 267.985 80.703 ;
 END
 PORT
  LAYER ME4 ;
  RECT 265.453 0.000 266.173 46.394 ;
 END
 PORT
  LAYER ME4 ;
  RECT 271.649 45.394 271.989 80.703 ;
 END
 PORT
  LAYER ME4 ;
  RECT 269.457 0.000 270.177 46.394 ;
 END
 PORT
  LAYER ME4 ;
  RECT 275.653 45.394 275.993 80.703 ;
 END
 PORT
  LAYER ME4 ;
  RECT 273.461 0.000 274.181 46.394 ;
 END
 PORT
  LAYER ME4 ;
  RECT 279.657 45.394 279.997 80.703 ;
 END
 PORT
  LAYER ME4 ;
  RECT 277.465 0.000 278.185 46.394 ;
 END
 PORT
  LAYER ME4 ;
  RECT 283.661 45.394 284.001 80.703 ;
 END
 PORT
  LAYER ME4 ;
  RECT 281.469 0.000 282.189 46.394 ;
 END
 PORT
  LAYER ME4 ;
  RECT 287.665 45.394 288.005 80.703 ;
 END
 PORT
  LAYER ME4 ;
  RECT 285.473 0.000 286.193 46.394 ;
 END
 PORT
  LAYER ME4 ;
  RECT 291.669 45.394 292.009 80.703 ;
 END
 PORT
  LAYER ME4 ;
  RECT 289.477 0.000 290.197 46.394 ;
 END
 PORT
  LAYER ME4 ;
  RECT 295.673 45.394 296.013 80.703 ;
 END
 PORT
  LAYER ME4 ;
  RECT 293.481 0.000 294.201 46.394 ;
 END
 PORT
  LAYER ME4 ;
  RECT 299.677 45.394 300.017 80.703 ;
 END
 PORT
  LAYER ME4 ;
  RECT 297.485 0.000 298.205 46.394 ;
 END
 PORT
  LAYER ME4 ;
  RECT 303.681 45.394 304.021 80.703 ;
 END
 PORT
  LAYER ME4 ;
  RECT 301.489 0.000 302.209 46.394 ;
 END
 PORT
  LAYER ME4 ;
  RECT 307.685 45.394 308.025 80.703 ;
 END
 PORT
  LAYER ME4 ;
  RECT 305.493 0.000 306.213 46.394 ;
 END
 PORT
  LAYER ME4 ;
  RECT 311.689 45.394 312.029 80.703 ;
 END
 PORT
  LAYER ME4 ;
  RECT 309.497 0.000 310.217 46.394 ;
 END
 PORT
  LAYER ME4 ;
  RECT 315.693 45.394 316.033 80.703 ;
 END
 PORT
  LAYER ME4 ;
  RECT 313.501 0.000 314.221 46.394 ;
 END
 PORT
  LAYER ME4 ;
  RECT 319.697 45.394 320.037 80.703 ;
 END
 PORT
  LAYER ME4 ;
  RECT 317.505 0.000 318.225 46.394 ;
 END
 PORT
  LAYER ME4 ;
  RECT 323.701 45.394 324.041 80.703 ;
 END
 PORT
  LAYER ME4 ;
  RECT 321.509 0.000 322.229 46.394 ;
 END
 PORT
  LAYER ME4 ;
  RECT 327.705 45.394 328.045 80.703 ;
 END
 PORT
  LAYER ME4 ;
  RECT 325.513 0.000 326.233 46.394 ;
 END
 PORT
  LAYER ME4 ;
  RECT 331.709 45.394 332.049 80.703 ;
 END
 PORT
  LAYER ME4 ;
  RECT 329.517 0.000 330.237 46.394 ;
 END
 PORT
  LAYER ME4 ;
  RECT 335.713 45.394 336.053 80.703 ;
 END
 PORT
  LAYER ME4 ;
  RECT 333.521 0.000 334.241 46.394 ;
 END
 PORT
  LAYER ME4 ;
  RECT 339.717 45.394 340.057 80.703 ;
 END
 PORT
  LAYER ME4 ;
  RECT 337.525 0.000 338.245 46.394 ;
 END
 PORT
  LAYER ME4 ;
  RECT 343.721 45.394 344.061 80.703 ;
 END
 PORT
  LAYER ME4 ;
  RECT 341.529 0.000 342.249 46.394 ;
 END
 PORT
  LAYER ME4 ;
  RECT 347.725 45.394 348.065 80.703 ;
 END
 PORT
  LAYER ME4 ;
  RECT 345.533 0.000 346.253 46.394 ;
 END
 PORT
  LAYER ME4 ;
  RECT 351.729 45.394 352.069 80.703 ;
 END
 PORT
  LAYER ME4 ;
  RECT 349.537 0.000 350.257 46.394 ;
 END
 PORT
  LAYER ME4 ;
  RECT 355.733 45.394 356.073 80.703 ;
 END
 PORT
  LAYER ME4 ;
  RECT 353.541 0.000 354.261 46.394 ;
 END
 PORT
  LAYER ME4 ;
  RECT 359.737 45.394 360.077 80.703 ;
 END
 PORT
  LAYER ME4 ;
  RECT 357.545 0.000 358.265 46.394 ;
 END
 PORT
  LAYER ME4 ;
  RECT 363.741 45.394 364.081 80.703 ;
 END
 PORT
  LAYER ME4 ;
  RECT 361.549 0.000 362.269 46.394 ;
 END
 PORT
  LAYER ME4 ;
  RECT 367.745 45.394 368.085 80.703 ;
 END
 PORT
  LAYER ME4 ;
  RECT 365.553 0.000 366.273 46.394 ;
 END
 PORT
  LAYER ME4 ;
  RECT 371.749 45.394 372.089 80.703 ;
 END
 PORT
  LAYER ME4 ;
  RECT 369.557 0.000 370.277 46.394 ;
 END
 PORT
  LAYER ME4 ;
  RECT 375.753 45.394 376.093 80.703 ;
 END
 PORT
  LAYER ME4 ;
  RECT 373.561 0.000 374.281 46.394 ;
 END
 PORT
  LAYER ME4 ;
  RECT 379.757 45.394 380.097 80.703 ;
 END
 PORT
  LAYER ME4 ;
  RECT 377.565 0.000 378.285 46.394 ;
 END
 PORT
  LAYER ME4 ;
  RECT 383.761 45.394 384.101 80.703 ;
 END
 PORT
  LAYER ME4 ;
  RECT 381.569 0.000 382.289 46.394 ;
 END
 PORT
  LAYER ME4 ;
  RECT 387.765 45.394 388.105 80.703 ;
 END
 PORT
  LAYER ME4 ;
  RECT 385.573 0.000 386.293 46.394 ;
 END
 PORT
  LAYER ME4 ;
  RECT 391.769 45.394 392.109 80.703 ;
 END
 PORT
  LAYER ME4 ;
  RECT 389.577 0.000 390.297 46.394 ;
 END
 PORT
  LAYER ME4 ;
  RECT 395.773 45.394 396.113 80.703 ;
 END
 PORT
  LAYER ME4 ;
  RECT 393.581 0.000 394.301 46.394 ;
 END
 PORT
  LAYER ME4 ;
  RECT 399.777 45.394 400.117 80.703 ;
 END
 PORT
  LAYER ME4 ;
  RECT 397.585 0.000 398.305 46.394 ;
 END
 PORT
  LAYER ME4 ;
  RECT 403.781 45.394 404.121 80.703 ;
 END
 PORT
  LAYER ME4 ;
  RECT 401.589 0.000 402.309 46.394 ;
 END
 PORT
  LAYER ME4 ;
  RECT 407.785 45.394 408.125 80.703 ;
 END
 PORT
  LAYER ME4 ;
  RECT 405.593 0.000 406.313 46.394 ;
 END
 PORT
  LAYER ME4 ;
  RECT 411.789 45.394 412.129 80.703 ;
 END
 PORT
  LAYER ME4 ;
  RECT 409.597 0.000 410.317 46.394 ;
 END
 PORT
  LAYER ME4 ;
  RECT 415.793 45.394 416.133 80.703 ;
 END
 PORT
  LAYER ME4 ;
  RECT 413.601 0.000 414.321 46.394 ;
 END
 PORT
  LAYER ME4 ;
  RECT 419.797 45.394 420.137 80.703 ;
 END
 PORT
  LAYER ME4 ;
  RECT 417.605 0.000 418.325 46.394 ;
 END
 PORT
  LAYER ME4 ;
  RECT 423.801 45.394 424.141 80.703 ;
 END
 PORT
  LAYER ME4 ;
  RECT 421.609 0.000 422.329 46.394 ;
 END
 PORT
  LAYER ME4 ;
  RECT 426.583 0.000 426.963 80.703 ;
 END
 PORT
  LAYER ME4 ;
  RECT 216.533 0.000 217.133 80.703 ;
 END
 PORT
  LAYER ME4 ;
  RECT 220.713 0.000 221.433 80.703 ;
 END
 PORT
  LAYER ME4 ;
  RECT 222.823 0.000 223.943 80.703 ;
 END
 PORT
  LAYER ME4 ;
  RECT 228.853 0.000 229.573 80.703 ;
 END
 PORT
  LAYER ME4 ;
  RECT 230.789 1.781 231.169 80.703 ;
 END
 PORT
  LAYER ME4 ;
  RECT 212.303 0.000 213.023 80.703 ;
 END
 PORT
  LAYER ME4 ;
  RECT 209.588 0.000 210.708 80.703 ;
 END
 PORT
  LAYER ME4 ;
  RECT 207.214 0.000 207.934 79.944 ;
 END
 PORT
  LAYER ME4 ;
  RECT 205.174 1.781 205.894 80.703 ;
 END
 PORT
  LAYER ME4 ;
  RECT 203.054 0.000 203.774 80.703 ;
 END
 PORT
  LAYER ME4 ;
  RECT 201.014 1.781 201.734 80.703 ;
 END
 PORT
  LAYER ME4 ;
  RECT 0.920 0.000 1.300 80.703 ;
 END
 PORT
  LAYER ME4 ;
  RECT 5.744 45.394 6.084 80.703 ;
 END
 PORT
  LAYER ME4 ;
  RECT 3.552 0.000 4.272 46.394 ;
 END
 PORT
  LAYER ME4 ;
  RECT 9.748 45.394 10.088 80.703 ;
 END
 PORT
  LAYER ME4 ;
  RECT 7.556 0.000 8.276 46.394 ;
 END
 PORT
  LAYER ME4 ;
  RECT 13.752 45.394 14.092 80.703 ;
 END
 PORT
  LAYER ME4 ;
  RECT 11.560 0.000 12.280 46.394 ;
 END
 PORT
  LAYER ME4 ;
  RECT 17.756 45.394 18.096 80.703 ;
 END
 PORT
  LAYER ME4 ;
  RECT 15.564 0.000 16.284 46.394 ;
 END
 PORT
  LAYER ME4 ;
  RECT 21.760 45.394 22.100 80.703 ;
 END
 PORT
  LAYER ME4 ;
  RECT 19.568 0.000 20.288 46.394 ;
 END
 PORT
  LAYER ME4 ;
  RECT 25.764 45.394 26.104 80.703 ;
 END
 PORT
  LAYER ME4 ;
  RECT 23.572 0.000 24.292 46.394 ;
 END
 PORT
  LAYER ME4 ;
  RECT 29.768 45.394 30.108 80.703 ;
 END
 PORT
  LAYER ME4 ;
  RECT 27.576 0.000 28.296 46.394 ;
 END
 PORT
  LAYER ME4 ;
  RECT 33.772 45.394 34.112 80.703 ;
 END
 PORT
  LAYER ME4 ;
  RECT 31.580 0.000 32.300 46.394 ;
 END
 PORT
  LAYER ME4 ;
  RECT 37.776 45.394 38.116 80.703 ;
 END
 PORT
  LAYER ME4 ;
  RECT 35.584 0.000 36.304 46.394 ;
 END
 PORT
  LAYER ME4 ;
  RECT 41.780 45.394 42.120 80.703 ;
 END
 PORT
  LAYER ME4 ;
  RECT 39.588 0.000 40.308 46.394 ;
 END
 PORT
  LAYER ME4 ;
  RECT 45.784 45.394 46.124 80.703 ;
 END
 PORT
  LAYER ME4 ;
  RECT 43.592 0.000 44.312 46.394 ;
 END
 PORT
  LAYER ME4 ;
  RECT 49.788 45.394 50.128 80.703 ;
 END
 PORT
  LAYER ME4 ;
  RECT 47.596 0.000 48.316 46.394 ;
 END
 PORT
  LAYER ME4 ;
  RECT 53.792 45.394 54.132 80.703 ;
 END
 PORT
  LAYER ME4 ;
  RECT 51.600 0.000 52.320 46.394 ;
 END
 PORT
  LAYER ME4 ;
  RECT 57.796 45.394 58.136 80.703 ;
 END
 PORT
  LAYER ME4 ;
  RECT 55.604 0.000 56.324 46.394 ;
 END
 PORT
  LAYER ME4 ;
  RECT 61.800 45.394 62.140 80.703 ;
 END
 PORT
  LAYER ME4 ;
  RECT 59.608 0.000 60.328 46.394 ;
 END
 PORT
  LAYER ME4 ;
  RECT 65.804 45.394 66.144 80.703 ;
 END
 PORT
  LAYER ME4 ;
  RECT 63.612 0.000 64.332 46.394 ;
 END
 PORT
  LAYER ME4 ;
  RECT 69.808 45.394 70.148 80.703 ;
 END
 PORT
  LAYER ME4 ;
  RECT 67.616 0.000 68.336 46.394 ;
 END
 PORT
  LAYER ME4 ;
  RECT 73.812 45.394 74.152 80.703 ;
 END
 PORT
  LAYER ME4 ;
  RECT 71.620 0.000 72.340 46.394 ;
 END
 PORT
  LAYER ME4 ;
  RECT 77.816 45.394 78.156 80.703 ;
 END
 PORT
  LAYER ME4 ;
  RECT 75.624 0.000 76.344 46.394 ;
 END
 PORT
  LAYER ME4 ;
  RECT 81.820 45.394 82.160 80.703 ;
 END
 PORT
  LAYER ME4 ;
  RECT 79.628 0.000 80.348 46.394 ;
 END
 PORT
  LAYER ME4 ;
  RECT 85.824 45.394 86.164 80.703 ;
 END
 PORT
  LAYER ME4 ;
  RECT 83.632 0.000 84.352 46.394 ;
 END
 PORT
  LAYER ME4 ;
  RECT 89.828 45.394 90.168 80.703 ;
 END
 PORT
  LAYER ME4 ;
  RECT 87.636 0.000 88.356 46.394 ;
 END
 PORT
  LAYER ME4 ;
  RECT 93.832 45.394 94.172 80.703 ;
 END
 PORT
  LAYER ME4 ;
  RECT 91.640 0.000 92.360 46.394 ;
 END
 PORT
  LAYER ME4 ;
  RECT 97.836 45.394 98.176 80.703 ;
 END
 PORT
  LAYER ME4 ;
  RECT 95.644 0.000 96.364 46.394 ;
 END
 PORT
  LAYER ME4 ;
  RECT 101.840 45.394 102.180 80.703 ;
 END
 PORT
  LAYER ME4 ;
  RECT 99.648 0.000 100.368 46.394 ;
 END
 PORT
  LAYER ME4 ;
  RECT 105.844 45.394 106.184 80.703 ;
 END
 PORT
  LAYER ME4 ;
  RECT 103.652 0.000 104.372 46.394 ;
 END
 PORT
  LAYER ME4 ;
  RECT 109.848 45.394 110.188 80.703 ;
 END
 PORT
  LAYER ME4 ;
  RECT 107.656 0.000 108.376 46.394 ;
 END
 PORT
  LAYER ME4 ;
  RECT 113.852 45.394 114.192 80.703 ;
 END
 PORT
  LAYER ME4 ;
  RECT 111.660 0.000 112.380 46.394 ;
 END
 PORT
  LAYER ME4 ;
  RECT 117.856 45.394 118.196 80.703 ;
 END
 PORT
  LAYER ME4 ;
  RECT 115.664 0.000 116.384 46.394 ;
 END
 PORT
  LAYER ME4 ;
  RECT 121.860 45.394 122.200 80.703 ;
 END
 PORT
  LAYER ME4 ;
  RECT 119.668 0.000 120.388 46.394 ;
 END
 PORT
  LAYER ME4 ;
  RECT 125.864 45.394 126.204 80.703 ;
 END
 PORT
  LAYER ME4 ;
  RECT 123.672 0.000 124.392 46.394 ;
 END
 PORT
  LAYER ME4 ;
  RECT 129.868 45.394 130.208 80.703 ;
 END
 PORT
  LAYER ME4 ;
  RECT 127.676 0.000 128.396 46.394 ;
 END
 PORT
  LAYER ME4 ;
  RECT 133.872 45.394 134.212 80.703 ;
 END
 PORT
  LAYER ME4 ;
  RECT 131.680 0.000 132.400 46.394 ;
 END
 PORT
  LAYER ME4 ;
  RECT 137.876 45.394 138.216 80.703 ;
 END
 PORT
  LAYER ME4 ;
  RECT 135.684 0.000 136.404 46.394 ;
 END
 PORT
  LAYER ME4 ;
  RECT 141.880 45.394 142.220 80.703 ;
 END
 PORT
  LAYER ME4 ;
  RECT 139.688 0.000 140.408 46.394 ;
 END
 PORT
  LAYER ME4 ;
  RECT 145.884 45.394 146.224 80.703 ;
 END
 PORT
  LAYER ME4 ;
  RECT 143.692 0.000 144.412 46.394 ;
 END
 PORT
  LAYER ME4 ;
  RECT 149.888 45.394 150.228 80.703 ;
 END
 PORT
  LAYER ME4 ;
  RECT 147.696 0.000 148.416 46.394 ;
 END
 PORT
  LAYER ME4 ;
  RECT 153.892 45.394 154.232 80.703 ;
 END
 PORT
  LAYER ME4 ;
  RECT 151.700 0.000 152.420 46.394 ;
 END
 PORT
  LAYER ME4 ;
  RECT 157.896 45.394 158.236 80.703 ;
 END
 PORT
  LAYER ME4 ;
  RECT 155.704 0.000 156.424 46.394 ;
 END
 PORT
  LAYER ME4 ;
  RECT 161.900 45.394 162.240 80.703 ;
 END
 PORT
  LAYER ME4 ;
  RECT 159.708 0.000 160.428 46.394 ;
 END
 PORT
  LAYER ME4 ;
  RECT 165.904 45.394 166.244 80.703 ;
 END
 PORT
  LAYER ME4 ;
  RECT 163.712 0.000 164.432 46.394 ;
 END
 PORT
  LAYER ME4 ;
  RECT 169.908 45.394 170.248 80.703 ;
 END
 PORT
  LAYER ME4 ;
  RECT 167.716 0.000 168.436 46.394 ;
 END
 PORT
  LAYER ME4 ;
  RECT 173.912 45.394 174.252 80.703 ;
 END
 PORT
  LAYER ME4 ;
  RECT 171.720 0.000 172.440 46.394 ;
 END
 PORT
  LAYER ME4 ;
  RECT 177.916 45.394 178.256 80.703 ;
 END
 PORT
  LAYER ME4 ;
  RECT 175.724 0.000 176.444 46.394 ;
 END
 PORT
  LAYER ME4 ;
  RECT 181.920 45.394 182.260 80.703 ;
 END
 PORT
  LAYER ME4 ;
  RECT 179.728 0.000 180.448 46.394 ;
 END
 PORT
  LAYER ME4 ;
  RECT 185.924 45.394 186.264 80.703 ;
 END
 PORT
  LAYER ME4 ;
  RECT 183.732 0.000 184.452 46.394 ;
 END
 PORT
  LAYER ME4 ;
  RECT 189.928 45.394 190.268 80.703 ;
 END
 PORT
  LAYER ME4 ;
  RECT 187.736 0.000 188.456 46.394 ;
 END
 PORT
  LAYER ME4 ;
  RECT 193.932 45.394 194.272 80.703 ;
 END
 PORT
  LAYER ME4 ;
  RECT 191.740 0.000 192.460 46.394 ;
 END
 PORT
  LAYER ME4 ;
  RECT 198.894 0.000 199.614 80.703 ;
 END
 PORT
  LAYER ME4 ;
  RECT 196.714 0.000 197.094 80.703 ;
 END
 PORT
  LAYER ME4 ;
  RECT 233.611 47.744 233.951 80.703 ;
 END
 PORT
  LAYER ME4 ;
  RECT 237.615 47.744 237.955 80.703 ;
 END
 PORT
  LAYER ME4 ;
  RECT 241.619 47.744 241.959 80.703 ;
 END
 PORT
  LAYER ME4 ;
  RECT 245.623 47.744 245.963 80.703 ;
 END
 PORT
  LAYER ME4 ;
  RECT 249.627 47.744 249.967 80.703 ;
 END
 PORT
  LAYER ME4 ;
  RECT 253.631 47.744 253.971 80.703 ;
 END
 PORT
  LAYER ME4 ;
  RECT 257.635 47.744 257.975 80.703 ;
 END
 PORT
  LAYER ME4 ;
  RECT 261.639 47.744 261.979 80.703 ;
 END
 PORT
  LAYER ME4 ;
  RECT 265.643 47.744 265.983 80.703 ;
 END
 PORT
  LAYER ME4 ;
  RECT 269.647 47.744 269.987 80.703 ;
 END
 PORT
  LAYER ME4 ;
  RECT 273.651 47.744 273.991 80.703 ;
 END
 PORT
  LAYER ME4 ;
  RECT 277.655 47.744 277.995 80.703 ;
 END
 PORT
  LAYER ME4 ;
  RECT 281.659 47.744 281.999 80.703 ;
 END
 PORT
  LAYER ME4 ;
  RECT 285.663 47.744 286.003 80.703 ;
 END
 PORT
  LAYER ME4 ;
  RECT 289.667 47.744 290.007 80.703 ;
 END
 PORT
  LAYER ME4 ;
  RECT 293.671 47.744 294.011 80.703 ;
 END
 PORT
  LAYER ME4 ;
  RECT 297.675 47.744 298.015 80.703 ;
 END
 PORT
  LAYER ME4 ;
  RECT 301.679 47.744 302.019 80.703 ;
 END
 PORT
  LAYER ME4 ;
  RECT 305.683 47.744 306.023 80.703 ;
 END
 PORT
  LAYER ME4 ;
  RECT 309.687 47.744 310.027 80.703 ;
 END
 PORT
  LAYER ME4 ;
  RECT 313.691 47.744 314.031 80.703 ;
 END
 PORT
  LAYER ME4 ;
  RECT 317.695 47.744 318.035 80.703 ;
 END
 PORT
  LAYER ME4 ;
  RECT 321.699 47.744 322.039 80.703 ;
 END
 PORT
  LAYER ME4 ;
  RECT 325.703 47.744 326.043 80.703 ;
 END
 PORT
  LAYER ME4 ;
  RECT 329.707 47.744 330.047 80.703 ;
 END
 PORT
  LAYER ME4 ;
  RECT 333.711 47.744 334.051 80.703 ;
 END
 PORT
  LAYER ME4 ;
  RECT 337.715 47.744 338.055 80.703 ;
 END
 PORT
  LAYER ME4 ;
  RECT 341.719 47.744 342.059 80.703 ;
 END
 PORT
  LAYER ME4 ;
  RECT 345.723 47.744 346.063 80.703 ;
 END
 PORT
  LAYER ME4 ;
  RECT 349.727 47.744 350.067 80.703 ;
 END
 PORT
  LAYER ME4 ;
  RECT 353.731 47.744 354.071 80.703 ;
 END
 PORT
  LAYER ME4 ;
  RECT 357.735 47.744 358.075 80.703 ;
 END
 PORT
  LAYER ME4 ;
  RECT 361.739 47.744 362.079 80.703 ;
 END
 PORT
  LAYER ME4 ;
  RECT 365.743 47.744 366.083 80.703 ;
 END
 PORT
  LAYER ME4 ;
  RECT 369.747 47.744 370.087 80.703 ;
 END
 PORT
  LAYER ME4 ;
  RECT 373.751 47.744 374.091 80.703 ;
 END
 PORT
  LAYER ME4 ;
  RECT 377.755 47.744 378.095 80.703 ;
 END
 PORT
  LAYER ME4 ;
  RECT 381.759 47.744 382.099 80.703 ;
 END
 PORT
  LAYER ME4 ;
  RECT 385.763 47.744 386.103 80.703 ;
 END
 PORT
  LAYER ME4 ;
  RECT 389.767 47.744 390.107 80.703 ;
 END
 PORT
  LAYER ME4 ;
  RECT 393.771 47.744 394.111 80.703 ;
 END
 PORT
  LAYER ME4 ;
  RECT 397.775 47.744 398.115 80.703 ;
 END
 PORT
  LAYER ME4 ;
  RECT 401.779 47.744 402.119 80.703 ;
 END
 PORT
  LAYER ME4 ;
  RECT 405.783 47.744 406.123 80.703 ;
 END
 PORT
  LAYER ME4 ;
  RECT 409.787 47.744 410.127 80.703 ;
 END
 PORT
  LAYER ME4 ;
  RECT 413.791 47.744 414.131 80.703 ;
 END
 PORT
  LAYER ME4 ;
  RECT 417.795 47.744 418.135 80.703 ;
 END
 PORT
  LAYER ME4 ;
  RECT 421.799 47.744 422.139 80.703 ;
 END
 PORT
  LAYER ME4 ;
  RECT 3.742 47.744 4.082 80.703 ;
 END
 PORT
  LAYER ME4 ;
  RECT 7.746 47.744 8.086 80.703 ;
 END
 PORT
  LAYER ME4 ;
  RECT 11.750 47.744 12.090 80.703 ;
 END
 PORT
  LAYER ME4 ;
  RECT 15.754 47.744 16.094 80.703 ;
 END
 PORT
  LAYER ME4 ;
  RECT 19.758 47.744 20.098 80.703 ;
 END
 PORT
  LAYER ME4 ;
  RECT 23.762 47.744 24.102 80.703 ;
 END
 PORT
  LAYER ME4 ;
  RECT 27.766 47.744 28.106 80.703 ;
 END
 PORT
  LAYER ME4 ;
  RECT 31.770 47.744 32.110 80.703 ;
 END
 PORT
  LAYER ME4 ;
  RECT 35.774 47.744 36.114 80.703 ;
 END
 PORT
  LAYER ME4 ;
  RECT 39.778 47.744 40.118 80.703 ;
 END
 PORT
  LAYER ME4 ;
  RECT 43.782 47.744 44.122 80.703 ;
 END
 PORT
  LAYER ME4 ;
  RECT 47.786 47.744 48.126 80.703 ;
 END
 PORT
  LAYER ME4 ;
  RECT 51.790 47.744 52.130 80.703 ;
 END
 PORT
  LAYER ME4 ;
  RECT 55.794 47.744 56.134 80.703 ;
 END
 PORT
  LAYER ME4 ;
  RECT 59.798 47.744 60.138 80.703 ;
 END
 PORT
  LAYER ME4 ;
  RECT 63.802 47.744 64.142 80.703 ;
 END
 PORT
  LAYER ME4 ;
  RECT 67.806 47.744 68.146 80.703 ;
 END
 PORT
  LAYER ME4 ;
  RECT 71.810 47.744 72.150 80.703 ;
 END
 PORT
  LAYER ME4 ;
  RECT 75.814 47.744 76.154 80.703 ;
 END
 PORT
  LAYER ME4 ;
  RECT 79.818 47.744 80.158 80.703 ;
 END
 PORT
  LAYER ME4 ;
  RECT 83.822 47.744 84.162 80.703 ;
 END
 PORT
  LAYER ME4 ;
  RECT 87.826 47.744 88.166 80.703 ;
 END
 PORT
  LAYER ME4 ;
  RECT 91.830 47.744 92.170 80.703 ;
 END
 PORT
  LAYER ME4 ;
  RECT 95.834 47.744 96.174 80.703 ;
 END
 PORT
  LAYER ME4 ;
  RECT 99.838 47.744 100.178 80.703 ;
 END
 PORT
  LAYER ME4 ;
  RECT 103.842 47.744 104.182 80.703 ;
 END
 PORT
  LAYER ME4 ;
  RECT 107.846 47.744 108.186 80.703 ;
 END
 PORT
  LAYER ME4 ;
  RECT 111.850 47.744 112.190 80.703 ;
 END
 PORT
  LAYER ME4 ;
  RECT 115.854 47.744 116.194 80.703 ;
 END
 PORT
  LAYER ME4 ;
  RECT 119.858 47.744 120.198 80.703 ;
 END
 PORT
  LAYER ME4 ;
  RECT 123.862 47.744 124.202 80.703 ;
 END
 PORT
  LAYER ME4 ;
  RECT 127.866 47.744 128.206 80.703 ;
 END
 PORT
  LAYER ME4 ;
  RECT 131.870 47.744 132.210 80.703 ;
 END
 PORT
  LAYER ME4 ;
  RECT 135.874 47.744 136.214 80.703 ;
 END
 PORT
  LAYER ME4 ;
  RECT 139.878 47.744 140.218 80.703 ;
 END
 PORT
  LAYER ME4 ;
  RECT 143.882 47.744 144.222 80.703 ;
 END
 PORT
  LAYER ME4 ;
  RECT 147.886 47.744 148.226 80.703 ;
 END
 PORT
  LAYER ME4 ;
  RECT 151.890 47.744 152.230 80.703 ;
 END
 PORT
  LAYER ME4 ;
  RECT 155.894 47.744 156.234 80.703 ;
 END
 PORT
  LAYER ME4 ;
  RECT 159.898 47.744 160.238 80.703 ;
 END
 PORT
  LAYER ME4 ;
  RECT 163.902 47.744 164.242 80.703 ;
 END
 PORT
  LAYER ME4 ;
  RECT 167.906 47.744 168.246 80.703 ;
 END
 PORT
  LAYER ME4 ;
  RECT 171.910 47.744 172.250 80.703 ;
 END
 PORT
  LAYER ME4 ;
  RECT 175.914 47.744 176.254 80.703 ;
 END
 PORT
  LAYER ME4 ;
  RECT 179.918 47.744 180.258 80.703 ;
 END
 PORT
  LAYER ME4 ;
  RECT 183.922 47.744 184.262 80.703 ;
 END
 PORT
  LAYER ME4 ;
  RECT 187.926 47.744 188.266 80.703 ;
 END
 PORT
  LAYER ME4 ;
  RECT 191.930 47.744 192.270 80.703 ;
 END
END VCC
PIN DI47
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 193.222 0.000 193.542 0.600 ;
  LAYER ME3 ;
  RECT 193.222 0.000 193.542 0.600 ;
  LAYER ME2 ;
  RECT 193.222 0.000 193.542 0.600 ;
  LAYER ME1 ;
  RECT 193.222 0.000 193.542 0.600 ;
 END
 ANTENNAPARTIALMETALAREA                  1.058 LAYER ME2 ;
 ANTENNAGATEAREA                          0.072 LAYER ME2 ;
 ANTENNAGATEAREA                          0.072 LAYER ME3 ;
 ANTENNAGATEAREA                          0.072 LAYER ME4 ;
 ANTENNADIFFAREA                          0.160 LAYER ME2 ;
 ANTENNADIFFAREA                          0.160 LAYER ME3 ;
 ANTENNADIFFAREA                          0.160 LAYER ME4 ;
 ANTENNAMAXAREACAR                       21.782 LAYER ME2 ;
 ANTENNAMAXAREACAR                       24.449 LAYER ME3 ;
 ANTENNAMAXAREACAR                       27.116 LAYER ME4 ;
END DI47
PIN DO47
  DIRECTION OUTPUT ;
 PORT
  LAYER ME4 ;
  RECT 192.660 0.000 192.980 0.600 ;
  LAYER ME3 ;
  RECT 192.660 0.000 192.980 0.600 ;
  LAYER ME2 ;
  RECT 192.660 0.000 192.980 0.600 ;
  LAYER ME1 ;
  RECT 192.660 0.000 192.980 0.600 ;
 END
 ANTENNAPARTIALMETALAREA                  5.273 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME3 ;
 ANTENNADIFFAREA                          1.293 LAYER ME4 ;
END DO47
PIN DI46
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 189.218 0.000 189.538 0.600 ;
  LAYER ME3 ;
  RECT 189.218 0.000 189.538 0.600 ;
  LAYER ME2 ;
  RECT 189.218 0.000 189.538 0.600 ;
  LAYER ME1 ;
  RECT 189.218 0.000 189.538 0.600 ;
 END
 ANTENNAPARTIALMETALAREA                  1.058 LAYER ME2 ;
 ANTENNAGATEAREA                          0.072 LAYER ME2 ;
 ANTENNAGATEAREA                          0.072 LAYER ME3 ;
 ANTENNAGATEAREA                          0.072 LAYER ME4 ;
 ANTENNADIFFAREA                          0.160 LAYER ME2 ;
 ANTENNADIFFAREA                          0.160 LAYER ME3 ;
 ANTENNADIFFAREA                          0.160 LAYER ME4 ;
 ANTENNAMAXAREACAR                       21.782 LAYER ME2 ;
 ANTENNAMAXAREACAR                       24.449 LAYER ME3 ;
 ANTENNAMAXAREACAR                       27.116 LAYER ME4 ;
END DI46
PIN DO46
  DIRECTION OUTPUT ;
 PORT
  LAYER ME4 ;
  RECT 188.656 0.000 188.976 0.600 ;
  LAYER ME3 ;
  RECT 188.656 0.000 188.976 0.600 ;
  LAYER ME2 ;
  RECT 188.656 0.000 188.976 0.600 ;
  LAYER ME1 ;
  RECT 188.656 0.000 188.976 0.600 ;
 END
 ANTENNAPARTIALMETALAREA                  5.273 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME3 ;
 ANTENNADIFFAREA                          1.293 LAYER ME4 ;
END DO46
PIN DI45
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 185.214 0.000 185.534 0.600 ;
  LAYER ME3 ;
  RECT 185.214 0.000 185.534 0.600 ;
  LAYER ME2 ;
  RECT 185.214 0.000 185.534 0.600 ;
  LAYER ME1 ;
  RECT 185.214 0.000 185.534 0.600 ;
 END
 ANTENNAPARTIALMETALAREA                  1.058 LAYER ME2 ;
 ANTENNAGATEAREA                          0.072 LAYER ME2 ;
 ANTENNAGATEAREA                          0.072 LAYER ME3 ;
 ANTENNAGATEAREA                          0.072 LAYER ME4 ;
 ANTENNADIFFAREA                          0.160 LAYER ME2 ;
 ANTENNADIFFAREA                          0.160 LAYER ME3 ;
 ANTENNADIFFAREA                          0.160 LAYER ME4 ;
 ANTENNAMAXAREACAR                       21.782 LAYER ME2 ;
 ANTENNAMAXAREACAR                       24.449 LAYER ME3 ;
 ANTENNAMAXAREACAR                       27.116 LAYER ME4 ;
END DI45
PIN DO45
  DIRECTION OUTPUT ;
 PORT
  LAYER ME4 ;
  RECT 184.652 0.000 184.972 0.600 ;
  LAYER ME3 ;
  RECT 184.652 0.000 184.972 0.600 ;
  LAYER ME2 ;
  RECT 184.652 0.000 184.972 0.600 ;
  LAYER ME1 ;
  RECT 184.652 0.000 184.972 0.600 ;
 END
 ANTENNAPARTIALMETALAREA                  5.273 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME3 ;
 ANTENNADIFFAREA                          1.293 LAYER ME4 ;
END DO45
PIN DI44
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 181.210 0.000 181.530 0.600 ;
  LAYER ME3 ;
  RECT 181.210 0.000 181.530 0.600 ;
  LAYER ME2 ;
  RECT 181.210 0.000 181.530 0.600 ;
  LAYER ME1 ;
  RECT 181.210 0.000 181.530 0.600 ;
 END
 ANTENNAPARTIALMETALAREA                  1.058 LAYER ME2 ;
 ANTENNAGATEAREA                          0.072 LAYER ME2 ;
 ANTENNAGATEAREA                          0.072 LAYER ME3 ;
 ANTENNAGATEAREA                          0.072 LAYER ME4 ;
 ANTENNADIFFAREA                          0.160 LAYER ME2 ;
 ANTENNADIFFAREA                          0.160 LAYER ME3 ;
 ANTENNADIFFAREA                          0.160 LAYER ME4 ;
 ANTENNAMAXAREACAR                       21.782 LAYER ME2 ;
 ANTENNAMAXAREACAR                       24.449 LAYER ME3 ;
 ANTENNAMAXAREACAR                       27.116 LAYER ME4 ;
END DI44
PIN DO44
  DIRECTION OUTPUT ;
 PORT
  LAYER ME4 ;
  RECT 180.648 0.000 180.968 0.600 ;
  LAYER ME3 ;
  RECT 180.648 0.000 180.968 0.600 ;
  LAYER ME2 ;
  RECT 180.648 0.000 180.968 0.600 ;
  LAYER ME1 ;
  RECT 180.648 0.000 180.968 0.600 ;
 END
 ANTENNAPARTIALMETALAREA                  5.273 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME3 ;
 ANTENNADIFFAREA                          1.293 LAYER ME4 ;
END DO44
PIN DI43
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 177.206 0.000 177.526 0.600 ;
  LAYER ME3 ;
  RECT 177.206 0.000 177.526 0.600 ;
  LAYER ME2 ;
  RECT 177.206 0.000 177.526 0.600 ;
  LAYER ME1 ;
  RECT 177.206 0.000 177.526 0.600 ;
 END
 ANTENNAPARTIALMETALAREA                  1.058 LAYER ME2 ;
 ANTENNAGATEAREA                          0.072 LAYER ME2 ;
 ANTENNAGATEAREA                          0.072 LAYER ME3 ;
 ANTENNAGATEAREA                          0.072 LAYER ME4 ;
 ANTENNADIFFAREA                          0.160 LAYER ME2 ;
 ANTENNADIFFAREA                          0.160 LAYER ME3 ;
 ANTENNADIFFAREA                          0.160 LAYER ME4 ;
 ANTENNAMAXAREACAR                       21.782 LAYER ME2 ;
 ANTENNAMAXAREACAR                       24.449 LAYER ME3 ;
 ANTENNAMAXAREACAR                       27.116 LAYER ME4 ;
END DI43
PIN DO43
  DIRECTION OUTPUT ;
 PORT
  LAYER ME4 ;
  RECT 176.644 0.000 176.964 0.600 ;
  LAYER ME3 ;
  RECT 176.644 0.000 176.964 0.600 ;
  LAYER ME2 ;
  RECT 176.644 0.000 176.964 0.600 ;
  LAYER ME1 ;
  RECT 176.644 0.000 176.964 0.600 ;
 END
 ANTENNAPARTIALMETALAREA                  5.273 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME3 ;
 ANTENNADIFFAREA                          1.293 LAYER ME4 ;
END DO43
PIN DI42
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 173.202 0.000 173.522 0.600 ;
  LAYER ME3 ;
  RECT 173.202 0.000 173.522 0.600 ;
  LAYER ME2 ;
  RECT 173.202 0.000 173.522 0.600 ;
  LAYER ME1 ;
  RECT 173.202 0.000 173.522 0.600 ;
 END
 ANTENNAPARTIALMETALAREA                  1.058 LAYER ME2 ;
 ANTENNAGATEAREA                          0.072 LAYER ME2 ;
 ANTENNAGATEAREA                          0.072 LAYER ME3 ;
 ANTENNAGATEAREA                          0.072 LAYER ME4 ;
 ANTENNADIFFAREA                          0.160 LAYER ME2 ;
 ANTENNADIFFAREA                          0.160 LAYER ME3 ;
 ANTENNADIFFAREA                          0.160 LAYER ME4 ;
 ANTENNAMAXAREACAR                       21.782 LAYER ME2 ;
 ANTENNAMAXAREACAR                       24.449 LAYER ME3 ;
 ANTENNAMAXAREACAR                       27.116 LAYER ME4 ;
END DI42
PIN DO42
  DIRECTION OUTPUT ;
 PORT
  LAYER ME4 ;
  RECT 172.640 0.000 172.960 0.600 ;
  LAYER ME3 ;
  RECT 172.640 0.000 172.960 0.600 ;
  LAYER ME2 ;
  RECT 172.640 0.000 172.960 0.600 ;
  LAYER ME1 ;
  RECT 172.640 0.000 172.960 0.600 ;
 END
 ANTENNAPARTIALMETALAREA                  5.273 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME3 ;
 ANTENNADIFFAREA                          1.293 LAYER ME4 ;
END DO42
PIN DI41
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 169.198 0.000 169.518 0.600 ;
  LAYER ME3 ;
  RECT 169.198 0.000 169.518 0.600 ;
  LAYER ME2 ;
  RECT 169.198 0.000 169.518 0.600 ;
  LAYER ME1 ;
  RECT 169.198 0.000 169.518 0.600 ;
 END
 ANTENNAPARTIALMETALAREA                  1.058 LAYER ME2 ;
 ANTENNAGATEAREA                          0.072 LAYER ME2 ;
 ANTENNAGATEAREA                          0.072 LAYER ME3 ;
 ANTENNAGATEAREA                          0.072 LAYER ME4 ;
 ANTENNADIFFAREA                          0.160 LAYER ME2 ;
 ANTENNADIFFAREA                          0.160 LAYER ME3 ;
 ANTENNADIFFAREA                          0.160 LAYER ME4 ;
 ANTENNAMAXAREACAR                       21.782 LAYER ME2 ;
 ANTENNAMAXAREACAR                       24.449 LAYER ME3 ;
 ANTENNAMAXAREACAR                       27.116 LAYER ME4 ;
END DI41
PIN DO41
  DIRECTION OUTPUT ;
 PORT
  LAYER ME4 ;
  RECT 168.636 0.000 168.956 0.600 ;
  LAYER ME3 ;
  RECT 168.636 0.000 168.956 0.600 ;
  LAYER ME2 ;
  RECT 168.636 0.000 168.956 0.600 ;
  LAYER ME1 ;
  RECT 168.636 0.000 168.956 0.600 ;
 END
 ANTENNAPARTIALMETALAREA                  5.273 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME3 ;
 ANTENNADIFFAREA                          1.293 LAYER ME4 ;
END DO41
PIN DI40
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 165.194 0.000 165.514 0.600 ;
  LAYER ME3 ;
  RECT 165.194 0.000 165.514 0.600 ;
  LAYER ME2 ;
  RECT 165.194 0.000 165.514 0.600 ;
  LAYER ME1 ;
  RECT 165.194 0.000 165.514 0.600 ;
 END
 ANTENNAPARTIALMETALAREA                  1.058 LAYER ME2 ;
 ANTENNAGATEAREA                          0.072 LAYER ME2 ;
 ANTENNAGATEAREA                          0.072 LAYER ME3 ;
 ANTENNAGATEAREA                          0.072 LAYER ME4 ;
 ANTENNADIFFAREA                          0.160 LAYER ME2 ;
 ANTENNADIFFAREA                          0.160 LAYER ME3 ;
 ANTENNADIFFAREA                          0.160 LAYER ME4 ;
 ANTENNAMAXAREACAR                       21.782 LAYER ME2 ;
 ANTENNAMAXAREACAR                       24.449 LAYER ME3 ;
 ANTENNAMAXAREACAR                       27.116 LAYER ME4 ;
END DI40
PIN DO40
  DIRECTION OUTPUT ;
 PORT
  LAYER ME4 ;
  RECT 164.632 0.000 164.952 0.600 ;
  LAYER ME3 ;
  RECT 164.632 0.000 164.952 0.600 ;
  LAYER ME2 ;
  RECT 164.632 0.000 164.952 0.600 ;
  LAYER ME1 ;
  RECT 164.632 0.000 164.952 0.600 ;
 END
 ANTENNAPARTIALMETALAREA                  5.273 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME3 ;
 ANTENNADIFFAREA                          1.293 LAYER ME4 ;
END DO40
PIN DI39
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 161.190 0.000 161.510 0.600 ;
  LAYER ME3 ;
  RECT 161.190 0.000 161.510 0.600 ;
  LAYER ME2 ;
  RECT 161.190 0.000 161.510 0.600 ;
  LAYER ME1 ;
  RECT 161.190 0.000 161.510 0.600 ;
 END
 ANTENNAPARTIALMETALAREA                  1.058 LAYER ME2 ;
 ANTENNAGATEAREA                          0.072 LAYER ME2 ;
 ANTENNAGATEAREA                          0.072 LAYER ME3 ;
 ANTENNAGATEAREA                          0.072 LAYER ME4 ;
 ANTENNADIFFAREA                          0.160 LAYER ME2 ;
 ANTENNADIFFAREA                          0.160 LAYER ME3 ;
 ANTENNADIFFAREA                          0.160 LAYER ME4 ;
 ANTENNAMAXAREACAR                       21.782 LAYER ME2 ;
 ANTENNAMAXAREACAR                       24.449 LAYER ME3 ;
 ANTENNAMAXAREACAR                       27.116 LAYER ME4 ;
END DI39
PIN DO39
  DIRECTION OUTPUT ;
 PORT
  LAYER ME4 ;
  RECT 160.628 0.000 160.948 0.600 ;
  LAYER ME3 ;
  RECT 160.628 0.000 160.948 0.600 ;
  LAYER ME2 ;
  RECT 160.628 0.000 160.948 0.600 ;
  LAYER ME1 ;
  RECT 160.628 0.000 160.948 0.600 ;
 END
 ANTENNAPARTIALMETALAREA                  5.273 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME3 ;
 ANTENNADIFFAREA                          1.293 LAYER ME4 ;
END DO39
PIN DI38
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 157.186 0.000 157.506 0.600 ;
  LAYER ME3 ;
  RECT 157.186 0.000 157.506 0.600 ;
  LAYER ME2 ;
  RECT 157.186 0.000 157.506 0.600 ;
  LAYER ME1 ;
  RECT 157.186 0.000 157.506 0.600 ;
 END
 ANTENNAPARTIALMETALAREA                  1.058 LAYER ME2 ;
 ANTENNAGATEAREA                          0.072 LAYER ME2 ;
 ANTENNAGATEAREA                          0.072 LAYER ME3 ;
 ANTENNAGATEAREA                          0.072 LAYER ME4 ;
 ANTENNADIFFAREA                          0.160 LAYER ME2 ;
 ANTENNADIFFAREA                          0.160 LAYER ME3 ;
 ANTENNADIFFAREA                          0.160 LAYER ME4 ;
 ANTENNAMAXAREACAR                       21.782 LAYER ME2 ;
 ANTENNAMAXAREACAR                       24.449 LAYER ME3 ;
 ANTENNAMAXAREACAR                       27.116 LAYER ME4 ;
END DI38
PIN DO38
  DIRECTION OUTPUT ;
 PORT
  LAYER ME4 ;
  RECT 156.624 0.000 156.944 0.600 ;
  LAYER ME3 ;
  RECT 156.624 0.000 156.944 0.600 ;
  LAYER ME2 ;
  RECT 156.624 0.000 156.944 0.600 ;
  LAYER ME1 ;
  RECT 156.624 0.000 156.944 0.600 ;
 END
 ANTENNAPARTIALMETALAREA                  5.273 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME3 ;
 ANTENNADIFFAREA                          1.293 LAYER ME4 ;
END DO38
PIN DI37
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 153.182 0.000 153.502 0.600 ;
  LAYER ME3 ;
  RECT 153.182 0.000 153.502 0.600 ;
  LAYER ME2 ;
  RECT 153.182 0.000 153.502 0.600 ;
  LAYER ME1 ;
  RECT 153.182 0.000 153.502 0.600 ;
 END
 ANTENNAPARTIALMETALAREA                  1.058 LAYER ME2 ;
 ANTENNAGATEAREA                          0.072 LAYER ME2 ;
 ANTENNAGATEAREA                          0.072 LAYER ME3 ;
 ANTENNAGATEAREA                          0.072 LAYER ME4 ;
 ANTENNADIFFAREA                          0.160 LAYER ME2 ;
 ANTENNADIFFAREA                          0.160 LAYER ME3 ;
 ANTENNADIFFAREA                          0.160 LAYER ME4 ;
 ANTENNAMAXAREACAR                       21.782 LAYER ME2 ;
 ANTENNAMAXAREACAR                       24.449 LAYER ME3 ;
 ANTENNAMAXAREACAR                       27.116 LAYER ME4 ;
END DI37
PIN DO37
  DIRECTION OUTPUT ;
 PORT
  LAYER ME4 ;
  RECT 152.620 0.000 152.940 0.600 ;
  LAYER ME3 ;
  RECT 152.620 0.000 152.940 0.600 ;
  LAYER ME2 ;
  RECT 152.620 0.000 152.940 0.600 ;
  LAYER ME1 ;
  RECT 152.620 0.000 152.940 0.600 ;
 END
 ANTENNAPARTIALMETALAREA                  5.273 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME3 ;
 ANTENNADIFFAREA                          1.293 LAYER ME4 ;
END DO37
PIN DI36
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 148.616 0.000 148.936 0.600 ;
  LAYER ME3 ;
  RECT 148.616 0.000 148.936 0.600 ;
  LAYER ME2 ;
  RECT 148.616 0.000 148.936 0.600 ;
  LAYER ME1 ;
  RECT 148.616 0.000 148.936 0.600 ;
 END
 ANTENNAPARTIALMETALAREA                  0.346 LAYER ME1 ;
 ANTENNAPARTIALMETALAREA                  1.466 LAYER ME2 ;
 ANTENNAPARTIALMETALAREA                  0.508 LAYER ME3 ;
 ANTENNAGATEAREA                          0.072 LAYER ME3 ;
 ANTENNAGATEAREA                          0.072 LAYER ME4 ;
 ANTENNADIFFAREA                          0.218 LAYER ME1 ;
 ANTENNADIFFAREA                          0.218 LAYER ME2 ;
 ANTENNADIFFAREA                          0.218 LAYER ME3 ;
 ANTENNADIFFAREA                          0.218 LAYER ME4 ;
 ANTENNAMAXAREACAR                       17.267 LAYER ME3 ;
 ANTENNAMAXAREACAR                       19.933 LAYER ME4 ;
END DI36
PIN DO36
  DIRECTION OUTPUT ;
 PORT
  LAYER ME4 ;
  RECT 149.178 0.000 149.498 0.600 ;
  LAYER ME3 ;
  RECT 149.178 0.000 149.498 0.600 ;
  LAYER ME2 ;
  RECT 149.178 0.000 149.498 0.600 ;
  LAYER ME1 ;
  RECT 149.178 0.000 149.498 0.600 ;
 END
 ANTENNAPARTIALMETALAREA                  5.602 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME3 ;
 ANTENNADIFFAREA                          1.293 LAYER ME4 ;
END DO36
PIN WEB3
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 147.176 0.000 147.496 0.600 ;
  LAYER ME3 ;
  RECT 147.176 0.000 147.496 0.600 ;
  LAYER ME2 ;
  RECT 147.176 0.000 147.496 0.600 ;
  LAYER ME1 ;
  RECT 147.176 0.000 147.496 0.600 ;
 END
 ANTENNAPARTIALMETALAREA                  1.036 LAYER ME2 ;
 ANTENNAGATEAREA                          0.288 LAYER ME2 ;
 ANTENNAGATEAREA                          0.288 LAYER ME3 ;
 ANTENNAGATEAREA                          0.288 LAYER ME4 ;
 ANTENNADIFFAREA                          0.206 LAYER ME2 ;
 ANTENNADIFFAREA                          0.206 LAYER ME3 ;
 ANTENNADIFFAREA                          0.206 LAYER ME4 ;
 ANTENNAMAXAREACAR                        5.844 LAYER ME2 ;
 ANTENNAMAXAREACAR                        6.511 LAYER ME3 ;
 ANTENNAMAXAREACAR                        7.178 LAYER ME4 ;
END WEB3
PIN DI35
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 145.174 0.000 145.494 0.600 ;
  LAYER ME3 ;
  RECT 145.174 0.000 145.494 0.600 ;
  LAYER ME2 ;
  RECT 145.174 0.000 145.494 0.600 ;
  LAYER ME1 ;
  RECT 145.174 0.000 145.494 0.600 ;
 END
 ANTENNAPARTIALMETALAREA                  1.058 LAYER ME2 ;
 ANTENNAGATEAREA                          0.072 LAYER ME2 ;
 ANTENNAGATEAREA                          0.072 LAYER ME3 ;
 ANTENNAGATEAREA                          0.072 LAYER ME4 ;
 ANTENNADIFFAREA                          0.160 LAYER ME2 ;
 ANTENNADIFFAREA                          0.160 LAYER ME3 ;
 ANTENNADIFFAREA                          0.160 LAYER ME4 ;
 ANTENNAMAXAREACAR                       21.782 LAYER ME2 ;
 ANTENNAMAXAREACAR                       24.449 LAYER ME3 ;
 ANTENNAMAXAREACAR                       27.116 LAYER ME4 ;
END DI35
PIN DO35
  DIRECTION OUTPUT ;
 PORT
  LAYER ME4 ;
  RECT 144.612 0.000 144.932 0.600 ;
  LAYER ME3 ;
  RECT 144.612 0.000 144.932 0.600 ;
  LAYER ME2 ;
  RECT 144.612 0.000 144.932 0.600 ;
  LAYER ME1 ;
  RECT 144.612 0.000 144.932 0.600 ;
 END
 ANTENNAPARTIALMETALAREA                  5.273 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME3 ;
 ANTENNADIFFAREA                          1.293 LAYER ME4 ;
END DO35
PIN DI34
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 141.170 0.000 141.490 0.600 ;
  LAYER ME3 ;
  RECT 141.170 0.000 141.490 0.600 ;
  LAYER ME2 ;
  RECT 141.170 0.000 141.490 0.600 ;
  LAYER ME1 ;
  RECT 141.170 0.000 141.490 0.600 ;
 END
 ANTENNAPARTIALMETALAREA                  1.058 LAYER ME2 ;
 ANTENNAGATEAREA                          0.072 LAYER ME2 ;
 ANTENNAGATEAREA                          0.072 LAYER ME3 ;
 ANTENNAGATEAREA                          0.072 LAYER ME4 ;
 ANTENNADIFFAREA                          0.160 LAYER ME2 ;
 ANTENNADIFFAREA                          0.160 LAYER ME3 ;
 ANTENNADIFFAREA                          0.160 LAYER ME4 ;
 ANTENNAMAXAREACAR                       21.782 LAYER ME2 ;
 ANTENNAMAXAREACAR                       24.449 LAYER ME3 ;
 ANTENNAMAXAREACAR                       27.116 LAYER ME4 ;
END DI34
PIN DO34
  DIRECTION OUTPUT ;
 PORT
  LAYER ME4 ;
  RECT 140.608 0.000 140.928 0.600 ;
  LAYER ME3 ;
  RECT 140.608 0.000 140.928 0.600 ;
  LAYER ME2 ;
  RECT 140.608 0.000 140.928 0.600 ;
  LAYER ME1 ;
  RECT 140.608 0.000 140.928 0.600 ;
 END
 ANTENNAPARTIALMETALAREA                  5.273 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME3 ;
 ANTENNADIFFAREA                          1.293 LAYER ME4 ;
END DO34
PIN DI33
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 137.166 0.000 137.486 0.600 ;
  LAYER ME3 ;
  RECT 137.166 0.000 137.486 0.600 ;
  LAYER ME2 ;
  RECT 137.166 0.000 137.486 0.600 ;
  LAYER ME1 ;
  RECT 137.166 0.000 137.486 0.600 ;
 END
 ANTENNAPARTIALMETALAREA                  1.058 LAYER ME2 ;
 ANTENNAGATEAREA                          0.072 LAYER ME2 ;
 ANTENNAGATEAREA                          0.072 LAYER ME3 ;
 ANTENNAGATEAREA                          0.072 LAYER ME4 ;
 ANTENNADIFFAREA                          0.160 LAYER ME2 ;
 ANTENNADIFFAREA                          0.160 LAYER ME3 ;
 ANTENNADIFFAREA                          0.160 LAYER ME4 ;
 ANTENNAMAXAREACAR                       21.782 LAYER ME2 ;
 ANTENNAMAXAREACAR                       24.449 LAYER ME3 ;
 ANTENNAMAXAREACAR                       27.116 LAYER ME4 ;
END DI33
PIN DO33
  DIRECTION OUTPUT ;
 PORT
  LAYER ME4 ;
  RECT 136.604 0.000 136.924 0.600 ;
  LAYER ME3 ;
  RECT 136.604 0.000 136.924 0.600 ;
  LAYER ME2 ;
  RECT 136.604 0.000 136.924 0.600 ;
  LAYER ME1 ;
  RECT 136.604 0.000 136.924 0.600 ;
 END
 ANTENNAPARTIALMETALAREA                  5.273 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME3 ;
 ANTENNADIFFAREA                          1.293 LAYER ME4 ;
END DO33
PIN DI32
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 133.162 0.000 133.482 0.600 ;
  LAYER ME3 ;
  RECT 133.162 0.000 133.482 0.600 ;
  LAYER ME2 ;
  RECT 133.162 0.000 133.482 0.600 ;
  LAYER ME1 ;
  RECT 133.162 0.000 133.482 0.600 ;
 END
 ANTENNAPARTIALMETALAREA                  1.058 LAYER ME2 ;
 ANTENNAGATEAREA                          0.072 LAYER ME2 ;
 ANTENNAGATEAREA                          0.072 LAYER ME3 ;
 ANTENNAGATEAREA                          0.072 LAYER ME4 ;
 ANTENNADIFFAREA                          0.160 LAYER ME2 ;
 ANTENNADIFFAREA                          0.160 LAYER ME3 ;
 ANTENNADIFFAREA                          0.160 LAYER ME4 ;
 ANTENNAMAXAREACAR                       21.782 LAYER ME2 ;
 ANTENNAMAXAREACAR                       24.449 LAYER ME3 ;
 ANTENNAMAXAREACAR                       27.116 LAYER ME4 ;
END DI32
PIN DO32
  DIRECTION OUTPUT ;
 PORT
  LAYER ME4 ;
  RECT 132.600 0.000 132.920 0.600 ;
  LAYER ME3 ;
  RECT 132.600 0.000 132.920 0.600 ;
  LAYER ME2 ;
  RECT 132.600 0.000 132.920 0.600 ;
  LAYER ME1 ;
  RECT 132.600 0.000 132.920 0.600 ;
 END
 ANTENNAPARTIALMETALAREA                  5.273 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME3 ;
 ANTENNADIFFAREA                          1.293 LAYER ME4 ;
END DO32
PIN DI31
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 129.158 0.000 129.478 0.600 ;
  LAYER ME3 ;
  RECT 129.158 0.000 129.478 0.600 ;
  LAYER ME2 ;
  RECT 129.158 0.000 129.478 0.600 ;
  LAYER ME1 ;
  RECT 129.158 0.000 129.478 0.600 ;
 END
 ANTENNAPARTIALMETALAREA                  1.058 LAYER ME2 ;
 ANTENNAGATEAREA                          0.072 LAYER ME2 ;
 ANTENNAGATEAREA                          0.072 LAYER ME3 ;
 ANTENNAGATEAREA                          0.072 LAYER ME4 ;
 ANTENNADIFFAREA                          0.160 LAYER ME2 ;
 ANTENNADIFFAREA                          0.160 LAYER ME3 ;
 ANTENNADIFFAREA                          0.160 LAYER ME4 ;
 ANTENNAMAXAREACAR                       21.782 LAYER ME2 ;
 ANTENNAMAXAREACAR                       24.449 LAYER ME3 ;
 ANTENNAMAXAREACAR                       27.116 LAYER ME4 ;
END DI31
PIN DO31
  DIRECTION OUTPUT ;
 PORT
  LAYER ME4 ;
  RECT 128.596 0.000 128.916 0.600 ;
  LAYER ME3 ;
  RECT 128.596 0.000 128.916 0.600 ;
  LAYER ME2 ;
  RECT 128.596 0.000 128.916 0.600 ;
  LAYER ME1 ;
  RECT 128.596 0.000 128.916 0.600 ;
 END
 ANTENNAPARTIALMETALAREA                  5.273 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME3 ;
 ANTENNADIFFAREA                          1.293 LAYER ME4 ;
END DO31
PIN DI30
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 125.154 0.000 125.474 0.600 ;
  LAYER ME3 ;
  RECT 125.154 0.000 125.474 0.600 ;
  LAYER ME2 ;
  RECT 125.154 0.000 125.474 0.600 ;
  LAYER ME1 ;
  RECT 125.154 0.000 125.474 0.600 ;
 END
 ANTENNAPARTIALMETALAREA                  1.058 LAYER ME2 ;
 ANTENNAGATEAREA                          0.072 LAYER ME2 ;
 ANTENNAGATEAREA                          0.072 LAYER ME3 ;
 ANTENNAGATEAREA                          0.072 LAYER ME4 ;
 ANTENNADIFFAREA                          0.160 LAYER ME2 ;
 ANTENNADIFFAREA                          0.160 LAYER ME3 ;
 ANTENNADIFFAREA                          0.160 LAYER ME4 ;
 ANTENNAMAXAREACAR                       21.782 LAYER ME2 ;
 ANTENNAMAXAREACAR                       24.449 LAYER ME3 ;
 ANTENNAMAXAREACAR                       27.116 LAYER ME4 ;
END DI30
PIN DO30
  DIRECTION OUTPUT ;
 PORT
  LAYER ME4 ;
  RECT 124.592 0.000 124.912 0.600 ;
  LAYER ME3 ;
  RECT 124.592 0.000 124.912 0.600 ;
  LAYER ME2 ;
  RECT 124.592 0.000 124.912 0.600 ;
  LAYER ME1 ;
  RECT 124.592 0.000 124.912 0.600 ;
 END
 ANTENNAPARTIALMETALAREA                  5.273 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME3 ;
 ANTENNADIFFAREA                          1.293 LAYER ME4 ;
END DO30
PIN DI29
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 121.150 0.000 121.470 0.600 ;
  LAYER ME3 ;
  RECT 121.150 0.000 121.470 0.600 ;
  LAYER ME2 ;
  RECT 121.150 0.000 121.470 0.600 ;
  LAYER ME1 ;
  RECT 121.150 0.000 121.470 0.600 ;
 END
 ANTENNAPARTIALMETALAREA                  1.058 LAYER ME2 ;
 ANTENNAGATEAREA                          0.072 LAYER ME2 ;
 ANTENNAGATEAREA                          0.072 LAYER ME3 ;
 ANTENNAGATEAREA                          0.072 LAYER ME4 ;
 ANTENNADIFFAREA                          0.160 LAYER ME2 ;
 ANTENNADIFFAREA                          0.160 LAYER ME3 ;
 ANTENNADIFFAREA                          0.160 LAYER ME4 ;
 ANTENNAMAXAREACAR                       21.782 LAYER ME2 ;
 ANTENNAMAXAREACAR                       24.449 LAYER ME3 ;
 ANTENNAMAXAREACAR                       27.116 LAYER ME4 ;
END DI29
PIN DO29
  DIRECTION OUTPUT ;
 PORT
  LAYER ME4 ;
  RECT 120.588 0.000 120.908 0.600 ;
  LAYER ME3 ;
  RECT 120.588 0.000 120.908 0.600 ;
  LAYER ME2 ;
  RECT 120.588 0.000 120.908 0.600 ;
  LAYER ME1 ;
  RECT 120.588 0.000 120.908 0.600 ;
 END
 ANTENNAPARTIALMETALAREA                  5.273 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME3 ;
 ANTENNADIFFAREA                          1.293 LAYER ME4 ;
END DO29
PIN DI28
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 117.146 0.000 117.466 0.600 ;
  LAYER ME3 ;
  RECT 117.146 0.000 117.466 0.600 ;
  LAYER ME2 ;
  RECT 117.146 0.000 117.466 0.600 ;
  LAYER ME1 ;
  RECT 117.146 0.000 117.466 0.600 ;
 END
 ANTENNAPARTIALMETALAREA                  1.058 LAYER ME2 ;
 ANTENNAGATEAREA                          0.072 LAYER ME2 ;
 ANTENNAGATEAREA                          0.072 LAYER ME3 ;
 ANTENNAGATEAREA                          0.072 LAYER ME4 ;
 ANTENNADIFFAREA                          0.160 LAYER ME2 ;
 ANTENNADIFFAREA                          0.160 LAYER ME3 ;
 ANTENNADIFFAREA                          0.160 LAYER ME4 ;
 ANTENNAMAXAREACAR                       21.782 LAYER ME2 ;
 ANTENNAMAXAREACAR                       24.449 LAYER ME3 ;
 ANTENNAMAXAREACAR                       27.116 LAYER ME4 ;
END DI28
PIN DO28
  DIRECTION OUTPUT ;
 PORT
  LAYER ME4 ;
  RECT 116.584 0.000 116.904 0.600 ;
  LAYER ME3 ;
  RECT 116.584 0.000 116.904 0.600 ;
  LAYER ME2 ;
  RECT 116.584 0.000 116.904 0.600 ;
  LAYER ME1 ;
  RECT 116.584 0.000 116.904 0.600 ;
 END
 ANTENNAPARTIALMETALAREA                  5.273 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME3 ;
 ANTENNADIFFAREA                          1.293 LAYER ME4 ;
END DO28
PIN DI27
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 113.142 0.000 113.462 0.600 ;
  LAYER ME3 ;
  RECT 113.142 0.000 113.462 0.600 ;
  LAYER ME2 ;
  RECT 113.142 0.000 113.462 0.600 ;
  LAYER ME1 ;
  RECT 113.142 0.000 113.462 0.600 ;
 END
 ANTENNAPARTIALMETALAREA                  1.058 LAYER ME2 ;
 ANTENNAGATEAREA                          0.072 LAYER ME2 ;
 ANTENNAGATEAREA                          0.072 LAYER ME3 ;
 ANTENNAGATEAREA                          0.072 LAYER ME4 ;
 ANTENNADIFFAREA                          0.160 LAYER ME2 ;
 ANTENNADIFFAREA                          0.160 LAYER ME3 ;
 ANTENNADIFFAREA                          0.160 LAYER ME4 ;
 ANTENNAMAXAREACAR                       21.782 LAYER ME2 ;
 ANTENNAMAXAREACAR                       24.449 LAYER ME3 ;
 ANTENNAMAXAREACAR                       27.116 LAYER ME4 ;
END DI27
PIN DO27
  DIRECTION OUTPUT ;
 PORT
  LAYER ME4 ;
  RECT 112.580 0.000 112.900 0.600 ;
  LAYER ME3 ;
  RECT 112.580 0.000 112.900 0.600 ;
  LAYER ME2 ;
  RECT 112.580 0.000 112.900 0.600 ;
  LAYER ME1 ;
  RECT 112.580 0.000 112.900 0.600 ;
 END
 ANTENNAPARTIALMETALAREA                  5.273 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME3 ;
 ANTENNADIFFAREA                          1.293 LAYER ME4 ;
END DO27
PIN DI26
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 109.138 0.000 109.458 0.600 ;
  LAYER ME3 ;
  RECT 109.138 0.000 109.458 0.600 ;
  LAYER ME2 ;
  RECT 109.138 0.000 109.458 0.600 ;
  LAYER ME1 ;
  RECT 109.138 0.000 109.458 0.600 ;
 END
 ANTENNAPARTIALMETALAREA                  1.058 LAYER ME2 ;
 ANTENNAGATEAREA                          0.072 LAYER ME2 ;
 ANTENNAGATEAREA                          0.072 LAYER ME3 ;
 ANTENNAGATEAREA                          0.072 LAYER ME4 ;
 ANTENNADIFFAREA                          0.160 LAYER ME2 ;
 ANTENNADIFFAREA                          0.160 LAYER ME3 ;
 ANTENNADIFFAREA                          0.160 LAYER ME4 ;
 ANTENNAMAXAREACAR                       21.782 LAYER ME2 ;
 ANTENNAMAXAREACAR                       24.449 LAYER ME3 ;
 ANTENNAMAXAREACAR                       27.116 LAYER ME4 ;
END DI26
PIN DO26
  DIRECTION OUTPUT ;
 PORT
  LAYER ME4 ;
  RECT 108.576 0.000 108.896 0.600 ;
  LAYER ME3 ;
  RECT 108.576 0.000 108.896 0.600 ;
  LAYER ME2 ;
  RECT 108.576 0.000 108.896 0.600 ;
  LAYER ME1 ;
  RECT 108.576 0.000 108.896 0.600 ;
 END
 ANTENNAPARTIALMETALAREA                  5.273 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME3 ;
 ANTENNADIFFAREA                          1.293 LAYER ME4 ;
END DO26
PIN DI25
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 105.134 0.000 105.454 0.600 ;
  LAYER ME3 ;
  RECT 105.134 0.000 105.454 0.600 ;
  LAYER ME2 ;
  RECT 105.134 0.000 105.454 0.600 ;
  LAYER ME1 ;
  RECT 105.134 0.000 105.454 0.600 ;
 END
 ANTENNAPARTIALMETALAREA                  1.058 LAYER ME2 ;
 ANTENNAGATEAREA                          0.072 LAYER ME2 ;
 ANTENNAGATEAREA                          0.072 LAYER ME3 ;
 ANTENNAGATEAREA                          0.072 LAYER ME4 ;
 ANTENNADIFFAREA                          0.160 LAYER ME2 ;
 ANTENNADIFFAREA                          0.160 LAYER ME3 ;
 ANTENNADIFFAREA                          0.160 LAYER ME4 ;
 ANTENNAMAXAREACAR                       21.782 LAYER ME2 ;
 ANTENNAMAXAREACAR                       24.449 LAYER ME3 ;
 ANTENNAMAXAREACAR                       27.116 LAYER ME4 ;
END DI25
PIN DO25
  DIRECTION OUTPUT ;
 PORT
  LAYER ME4 ;
  RECT 104.572 0.000 104.892 0.600 ;
  LAYER ME3 ;
  RECT 104.572 0.000 104.892 0.600 ;
  LAYER ME2 ;
  RECT 104.572 0.000 104.892 0.600 ;
  LAYER ME1 ;
  RECT 104.572 0.000 104.892 0.600 ;
 END
 ANTENNAPARTIALMETALAREA                  5.273 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME3 ;
 ANTENNADIFFAREA                          1.293 LAYER ME4 ;
END DO25
PIN DI24
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 100.568 0.000 100.888 0.600 ;
  LAYER ME3 ;
  RECT 100.568 0.000 100.888 0.600 ;
  LAYER ME2 ;
  RECT 100.568 0.000 100.888 0.600 ;
  LAYER ME1 ;
  RECT 100.568 0.000 100.888 0.600 ;
 END
 ANTENNAPARTIALMETALAREA                  0.346 LAYER ME1 ;
 ANTENNAPARTIALMETALAREA                  1.466 LAYER ME2 ;
 ANTENNAPARTIALMETALAREA                  0.508 LAYER ME3 ;
 ANTENNAGATEAREA                          0.072 LAYER ME3 ;
 ANTENNAGATEAREA                          0.072 LAYER ME4 ;
 ANTENNADIFFAREA                          0.218 LAYER ME1 ;
 ANTENNADIFFAREA                          0.218 LAYER ME2 ;
 ANTENNADIFFAREA                          0.218 LAYER ME3 ;
 ANTENNADIFFAREA                          0.218 LAYER ME4 ;
 ANTENNAMAXAREACAR                       17.267 LAYER ME3 ;
 ANTENNAMAXAREACAR                       19.933 LAYER ME4 ;
END DI24
PIN DO24
  DIRECTION OUTPUT ;
 PORT
  LAYER ME4 ;
  RECT 101.130 0.000 101.450 0.600 ;
  LAYER ME3 ;
  RECT 101.130 0.000 101.450 0.600 ;
  LAYER ME2 ;
  RECT 101.130 0.000 101.450 0.600 ;
  LAYER ME1 ;
  RECT 101.130 0.000 101.450 0.600 ;
 END
 ANTENNAPARTIALMETALAREA                  5.602 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME3 ;
 ANTENNADIFFAREA                          1.293 LAYER ME4 ;
END DO24
PIN WEB2
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 99.128 0.000 99.448 0.600 ;
  LAYER ME3 ;
  RECT 99.128 0.000 99.448 0.600 ;
  LAYER ME2 ;
  RECT 99.128 0.000 99.448 0.600 ;
  LAYER ME1 ;
  RECT 99.128 0.000 99.448 0.600 ;
 END
 ANTENNAPARTIALMETALAREA                  1.036 LAYER ME2 ;
 ANTENNAGATEAREA                          0.288 LAYER ME2 ;
 ANTENNAGATEAREA                          0.288 LAYER ME3 ;
 ANTENNAGATEAREA                          0.288 LAYER ME4 ;
 ANTENNADIFFAREA                          0.206 LAYER ME2 ;
 ANTENNADIFFAREA                          0.206 LAYER ME3 ;
 ANTENNADIFFAREA                          0.206 LAYER ME4 ;
 ANTENNAMAXAREACAR                        5.844 LAYER ME2 ;
 ANTENNAMAXAREACAR                        6.511 LAYER ME3 ;
 ANTENNAMAXAREACAR                        7.178 LAYER ME4 ;
END WEB2
PIN DI23
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 97.126 0.000 97.446 0.600 ;
  LAYER ME3 ;
  RECT 97.126 0.000 97.446 0.600 ;
  LAYER ME2 ;
  RECT 97.126 0.000 97.446 0.600 ;
  LAYER ME1 ;
  RECT 97.126 0.000 97.446 0.600 ;
 END
 ANTENNAPARTIALMETALAREA                  1.058 LAYER ME2 ;
 ANTENNAGATEAREA                          0.072 LAYER ME2 ;
 ANTENNAGATEAREA                          0.072 LAYER ME3 ;
 ANTENNAGATEAREA                          0.072 LAYER ME4 ;
 ANTENNADIFFAREA                          0.160 LAYER ME2 ;
 ANTENNADIFFAREA                          0.160 LAYER ME3 ;
 ANTENNADIFFAREA                          0.160 LAYER ME4 ;
 ANTENNAMAXAREACAR                       21.782 LAYER ME2 ;
 ANTENNAMAXAREACAR                       24.449 LAYER ME3 ;
 ANTENNAMAXAREACAR                       27.116 LAYER ME4 ;
END DI23
PIN DO23
  DIRECTION OUTPUT ;
 PORT
  LAYER ME4 ;
  RECT 96.564 0.000 96.884 0.600 ;
  LAYER ME3 ;
  RECT 96.564 0.000 96.884 0.600 ;
  LAYER ME2 ;
  RECT 96.564 0.000 96.884 0.600 ;
  LAYER ME1 ;
  RECT 96.564 0.000 96.884 0.600 ;
 END
 ANTENNAPARTIALMETALAREA                  5.273 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME3 ;
 ANTENNADIFFAREA                          1.293 LAYER ME4 ;
END DO23
PIN DI22
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 93.122 0.000 93.442 0.600 ;
  LAYER ME3 ;
  RECT 93.122 0.000 93.442 0.600 ;
  LAYER ME2 ;
  RECT 93.122 0.000 93.442 0.600 ;
  LAYER ME1 ;
  RECT 93.122 0.000 93.442 0.600 ;
 END
 ANTENNAPARTIALMETALAREA                  1.058 LAYER ME2 ;
 ANTENNAGATEAREA                          0.072 LAYER ME2 ;
 ANTENNAGATEAREA                          0.072 LAYER ME3 ;
 ANTENNAGATEAREA                          0.072 LAYER ME4 ;
 ANTENNADIFFAREA                          0.160 LAYER ME2 ;
 ANTENNADIFFAREA                          0.160 LAYER ME3 ;
 ANTENNADIFFAREA                          0.160 LAYER ME4 ;
 ANTENNAMAXAREACAR                       21.782 LAYER ME2 ;
 ANTENNAMAXAREACAR                       24.449 LAYER ME3 ;
 ANTENNAMAXAREACAR                       27.116 LAYER ME4 ;
END DI22
PIN DO22
  DIRECTION OUTPUT ;
 PORT
  LAYER ME4 ;
  RECT 92.560 0.000 92.880 0.600 ;
  LAYER ME3 ;
  RECT 92.560 0.000 92.880 0.600 ;
  LAYER ME2 ;
  RECT 92.560 0.000 92.880 0.600 ;
  LAYER ME1 ;
  RECT 92.560 0.000 92.880 0.600 ;
 END
 ANTENNAPARTIALMETALAREA                  5.273 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME3 ;
 ANTENNADIFFAREA                          1.293 LAYER ME4 ;
END DO22
PIN DI21
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 89.118 0.000 89.438 0.600 ;
  LAYER ME3 ;
  RECT 89.118 0.000 89.438 0.600 ;
  LAYER ME2 ;
  RECT 89.118 0.000 89.438 0.600 ;
  LAYER ME1 ;
  RECT 89.118 0.000 89.438 0.600 ;
 END
 ANTENNAPARTIALMETALAREA                  1.058 LAYER ME2 ;
 ANTENNAGATEAREA                          0.072 LAYER ME2 ;
 ANTENNAGATEAREA                          0.072 LAYER ME3 ;
 ANTENNAGATEAREA                          0.072 LAYER ME4 ;
 ANTENNADIFFAREA                          0.160 LAYER ME2 ;
 ANTENNADIFFAREA                          0.160 LAYER ME3 ;
 ANTENNADIFFAREA                          0.160 LAYER ME4 ;
 ANTENNAMAXAREACAR                       21.782 LAYER ME2 ;
 ANTENNAMAXAREACAR                       24.449 LAYER ME3 ;
 ANTENNAMAXAREACAR                       27.116 LAYER ME4 ;
END DI21
PIN DO21
  DIRECTION OUTPUT ;
 PORT
  LAYER ME4 ;
  RECT 88.556 0.000 88.876 0.600 ;
  LAYER ME3 ;
  RECT 88.556 0.000 88.876 0.600 ;
  LAYER ME2 ;
  RECT 88.556 0.000 88.876 0.600 ;
  LAYER ME1 ;
  RECT 88.556 0.000 88.876 0.600 ;
 END
 ANTENNAPARTIALMETALAREA                  5.273 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME3 ;
 ANTENNADIFFAREA                          1.293 LAYER ME4 ;
END DO21
PIN DI20
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 85.114 0.000 85.434 0.600 ;
  LAYER ME3 ;
  RECT 85.114 0.000 85.434 0.600 ;
  LAYER ME2 ;
  RECT 85.114 0.000 85.434 0.600 ;
  LAYER ME1 ;
  RECT 85.114 0.000 85.434 0.600 ;
 END
 ANTENNAPARTIALMETALAREA                  1.058 LAYER ME2 ;
 ANTENNAGATEAREA                          0.072 LAYER ME2 ;
 ANTENNAGATEAREA                          0.072 LAYER ME3 ;
 ANTENNAGATEAREA                          0.072 LAYER ME4 ;
 ANTENNADIFFAREA                          0.160 LAYER ME2 ;
 ANTENNADIFFAREA                          0.160 LAYER ME3 ;
 ANTENNADIFFAREA                          0.160 LAYER ME4 ;
 ANTENNAMAXAREACAR                       21.782 LAYER ME2 ;
 ANTENNAMAXAREACAR                       24.449 LAYER ME3 ;
 ANTENNAMAXAREACAR                       27.116 LAYER ME4 ;
END DI20
PIN DO20
  DIRECTION OUTPUT ;
 PORT
  LAYER ME4 ;
  RECT 84.552 0.000 84.872 0.600 ;
  LAYER ME3 ;
  RECT 84.552 0.000 84.872 0.600 ;
  LAYER ME2 ;
  RECT 84.552 0.000 84.872 0.600 ;
  LAYER ME1 ;
  RECT 84.552 0.000 84.872 0.600 ;
 END
 ANTENNAPARTIALMETALAREA                  5.273 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME3 ;
 ANTENNADIFFAREA                          1.293 LAYER ME4 ;
END DO20
PIN DI19
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 81.110 0.000 81.430 0.600 ;
  LAYER ME3 ;
  RECT 81.110 0.000 81.430 0.600 ;
  LAYER ME2 ;
  RECT 81.110 0.000 81.430 0.600 ;
  LAYER ME1 ;
  RECT 81.110 0.000 81.430 0.600 ;
 END
 ANTENNAPARTIALMETALAREA                  1.058 LAYER ME2 ;
 ANTENNAGATEAREA                          0.072 LAYER ME2 ;
 ANTENNAGATEAREA                          0.072 LAYER ME3 ;
 ANTENNAGATEAREA                          0.072 LAYER ME4 ;
 ANTENNADIFFAREA                          0.160 LAYER ME2 ;
 ANTENNADIFFAREA                          0.160 LAYER ME3 ;
 ANTENNADIFFAREA                          0.160 LAYER ME4 ;
 ANTENNAMAXAREACAR                       21.782 LAYER ME2 ;
 ANTENNAMAXAREACAR                       24.449 LAYER ME3 ;
 ANTENNAMAXAREACAR                       27.116 LAYER ME4 ;
END DI19
PIN DO19
  DIRECTION OUTPUT ;
 PORT
  LAYER ME4 ;
  RECT 80.548 0.000 80.868 0.600 ;
  LAYER ME3 ;
  RECT 80.548 0.000 80.868 0.600 ;
  LAYER ME2 ;
  RECT 80.548 0.000 80.868 0.600 ;
  LAYER ME1 ;
  RECT 80.548 0.000 80.868 0.600 ;
 END
 ANTENNAPARTIALMETALAREA                  5.273 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME3 ;
 ANTENNADIFFAREA                          1.293 LAYER ME4 ;
END DO19
PIN DI18
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 77.106 0.000 77.426 0.600 ;
  LAYER ME3 ;
  RECT 77.106 0.000 77.426 0.600 ;
  LAYER ME2 ;
  RECT 77.106 0.000 77.426 0.600 ;
  LAYER ME1 ;
  RECT 77.106 0.000 77.426 0.600 ;
 END
 ANTENNAPARTIALMETALAREA                  1.058 LAYER ME2 ;
 ANTENNAGATEAREA                          0.072 LAYER ME2 ;
 ANTENNAGATEAREA                          0.072 LAYER ME3 ;
 ANTENNAGATEAREA                          0.072 LAYER ME4 ;
 ANTENNADIFFAREA                          0.160 LAYER ME2 ;
 ANTENNADIFFAREA                          0.160 LAYER ME3 ;
 ANTENNADIFFAREA                          0.160 LAYER ME4 ;
 ANTENNAMAXAREACAR                       21.782 LAYER ME2 ;
 ANTENNAMAXAREACAR                       24.449 LAYER ME3 ;
 ANTENNAMAXAREACAR                       27.116 LAYER ME4 ;
END DI18
PIN DO18
  DIRECTION OUTPUT ;
 PORT
  LAYER ME4 ;
  RECT 76.544 0.000 76.864 0.600 ;
  LAYER ME3 ;
  RECT 76.544 0.000 76.864 0.600 ;
  LAYER ME2 ;
  RECT 76.544 0.000 76.864 0.600 ;
  LAYER ME1 ;
  RECT 76.544 0.000 76.864 0.600 ;
 END
 ANTENNAPARTIALMETALAREA                  5.273 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME3 ;
 ANTENNADIFFAREA                          1.293 LAYER ME4 ;
END DO18
PIN DI17
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 73.102 0.000 73.422 0.600 ;
  LAYER ME3 ;
  RECT 73.102 0.000 73.422 0.600 ;
  LAYER ME2 ;
  RECT 73.102 0.000 73.422 0.600 ;
  LAYER ME1 ;
  RECT 73.102 0.000 73.422 0.600 ;
 END
 ANTENNAPARTIALMETALAREA                  1.058 LAYER ME2 ;
 ANTENNAGATEAREA                          0.072 LAYER ME2 ;
 ANTENNAGATEAREA                          0.072 LAYER ME3 ;
 ANTENNAGATEAREA                          0.072 LAYER ME4 ;
 ANTENNADIFFAREA                          0.160 LAYER ME2 ;
 ANTENNADIFFAREA                          0.160 LAYER ME3 ;
 ANTENNADIFFAREA                          0.160 LAYER ME4 ;
 ANTENNAMAXAREACAR                       21.782 LAYER ME2 ;
 ANTENNAMAXAREACAR                       24.449 LAYER ME3 ;
 ANTENNAMAXAREACAR                       27.116 LAYER ME4 ;
END DI17
PIN DO17
  DIRECTION OUTPUT ;
 PORT
  LAYER ME4 ;
  RECT 72.540 0.000 72.860 0.600 ;
  LAYER ME3 ;
  RECT 72.540 0.000 72.860 0.600 ;
  LAYER ME2 ;
  RECT 72.540 0.000 72.860 0.600 ;
  LAYER ME1 ;
  RECT 72.540 0.000 72.860 0.600 ;
 END
 ANTENNAPARTIALMETALAREA                  5.273 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME3 ;
 ANTENNADIFFAREA                          1.293 LAYER ME4 ;
END DO17
PIN DI16
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 69.098 0.000 69.418 0.600 ;
  LAYER ME3 ;
  RECT 69.098 0.000 69.418 0.600 ;
  LAYER ME2 ;
  RECT 69.098 0.000 69.418 0.600 ;
  LAYER ME1 ;
  RECT 69.098 0.000 69.418 0.600 ;
 END
 ANTENNAPARTIALMETALAREA                  1.058 LAYER ME2 ;
 ANTENNAGATEAREA                          0.072 LAYER ME2 ;
 ANTENNAGATEAREA                          0.072 LAYER ME3 ;
 ANTENNAGATEAREA                          0.072 LAYER ME4 ;
 ANTENNADIFFAREA                          0.160 LAYER ME2 ;
 ANTENNADIFFAREA                          0.160 LAYER ME3 ;
 ANTENNADIFFAREA                          0.160 LAYER ME4 ;
 ANTENNAMAXAREACAR                       21.782 LAYER ME2 ;
 ANTENNAMAXAREACAR                       24.449 LAYER ME3 ;
 ANTENNAMAXAREACAR                       27.116 LAYER ME4 ;
END DI16
PIN DO16
  DIRECTION OUTPUT ;
 PORT
  LAYER ME4 ;
  RECT 68.536 0.000 68.856 0.600 ;
  LAYER ME3 ;
  RECT 68.536 0.000 68.856 0.600 ;
  LAYER ME2 ;
  RECT 68.536 0.000 68.856 0.600 ;
  LAYER ME1 ;
  RECT 68.536 0.000 68.856 0.600 ;
 END
 ANTENNAPARTIALMETALAREA                  5.273 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME3 ;
 ANTENNADIFFAREA                          1.293 LAYER ME4 ;
END DO16
PIN DI15
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 65.094 0.000 65.414 0.600 ;
  LAYER ME3 ;
  RECT 65.094 0.000 65.414 0.600 ;
  LAYER ME2 ;
  RECT 65.094 0.000 65.414 0.600 ;
  LAYER ME1 ;
  RECT 65.094 0.000 65.414 0.600 ;
 END
 ANTENNAPARTIALMETALAREA                  1.058 LAYER ME2 ;
 ANTENNAGATEAREA                          0.072 LAYER ME2 ;
 ANTENNAGATEAREA                          0.072 LAYER ME3 ;
 ANTENNAGATEAREA                          0.072 LAYER ME4 ;
 ANTENNADIFFAREA                          0.160 LAYER ME2 ;
 ANTENNADIFFAREA                          0.160 LAYER ME3 ;
 ANTENNADIFFAREA                          0.160 LAYER ME4 ;
 ANTENNAMAXAREACAR                       21.782 LAYER ME2 ;
 ANTENNAMAXAREACAR                       24.449 LAYER ME3 ;
 ANTENNAMAXAREACAR                       27.116 LAYER ME4 ;
END DI15
PIN DO15
  DIRECTION OUTPUT ;
 PORT
  LAYER ME4 ;
  RECT 64.532 0.000 64.852 0.600 ;
  LAYER ME3 ;
  RECT 64.532 0.000 64.852 0.600 ;
  LAYER ME2 ;
  RECT 64.532 0.000 64.852 0.600 ;
  LAYER ME1 ;
  RECT 64.532 0.000 64.852 0.600 ;
 END
 ANTENNAPARTIALMETALAREA                  5.273 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME3 ;
 ANTENNADIFFAREA                          1.293 LAYER ME4 ;
END DO15
PIN DI14
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 61.090 0.000 61.410 0.600 ;
  LAYER ME3 ;
  RECT 61.090 0.000 61.410 0.600 ;
  LAYER ME2 ;
  RECT 61.090 0.000 61.410 0.600 ;
  LAYER ME1 ;
  RECT 61.090 0.000 61.410 0.600 ;
 END
 ANTENNAPARTIALMETALAREA                  1.058 LAYER ME2 ;
 ANTENNAGATEAREA                          0.072 LAYER ME2 ;
 ANTENNAGATEAREA                          0.072 LAYER ME3 ;
 ANTENNAGATEAREA                          0.072 LAYER ME4 ;
 ANTENNADIFFAREA                          0.160 LAYER ME2 ;
 ANTENNADIFFAREA                          0.160 LAYER ME3 ;
 ANTENNADIFFAREA                          0.160 LAYER ME4 ;
 ANTENNAMAXAREACAR                       21.782 LAYER ME2 ;
 ANTENNAMAXAREACAR                       24.449 LAYER ME3 ;
 ANTENNAMAXAREACAR                       27.116 LAYER ME4 ;
END DI14
PIN DO14
  DIRECTION OUTPUT ;
 PORT
  LAYER ME4 ;
  RECT 60.528 0.000 60.848 0.600 ;
  LAYER ME3 ;
  RECT 60.528 0.000 60.848 0.600 ;
  LAYER ME2 ;
  RECT 60.528 0.000 60.848 0.600 ;
  LAYER ME1 ;
  RECT 60.528 0.000 60.848 0.600 ;
 END
 ANTENNAPARTIALMETALAREA                  5.273 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME3 ;
 ANTENNADIFFAREA                          1.293 LAYER ME4 ;
END DO14
PIN DI13
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 57.086 0.000 57.406 0.600 ;
  LAYER ME3 ;
  RECT 57.086 0.000 57.406 0.600 ;
  LAYER ME2 ;
  RECT 57.086 0.000 57.406 0.600 ;
  LAYER ME1 ;
  RECT 57.086 0.000 57.406 0.600 ;
 END
 ANTENNAPARTIALMETALAREA                  1.058 LAYER ME2 ;
 ANTENNAGATEAREA                          0.072 LAYER ME2 ;
 ANTENNAGATEAREA                          0.072 LAYER ME3 ;
 ANTENNAGATEAREA                          0.072 LAYER ME4 ;
 ANTENNADIFFAREA                          0.160 LAYER ME2 ;
 ANTENNADIFFAREA                          0.160 LAYER ME3 ;
 ANTENNADIFFAREA                          0.160 LAYER ME4 ;
 ANTENNAMAXAREACAR                       21.782 LAYER ME2 ;
 ANTENNAMAXAREACAR                       24.449 LAYER ME3 ;
 ANTENNAMAXAREACAR                       27.116 LAYER ME4 ;
END DI13
PIN DO13
  DIRECTION OUTPUT ;
 PORT
  LAYER ME4 ;
  RECT 56.524 0.000 56.844 0.600 ;
  LAYER ME3 ;
  RECT 56.524 0.000 56.844 0.600 ;
  LAYER ME2 ;
  RECT 56.524 0.000 56.844 0.600 ;
  LAYER ME1 ;
  RECT 56.524 0.000 56.844 0.600 ;
 END
 ANTENNAPARTIALMETALAREA                  5.273 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME3 ;
 ANTENNADIFFAREA                          1.293 LAYER ME4 ;
END DO13
PIN DI12
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 52.520 0.000 52.840 0.600 ;
  LAYER ME3 ;
  RECT 52.520 0.000 52.840 0.600 ;
  LAYER ME2 ;
  RECT 52.520 0.000 52.840 0.600 ;
  LAYER ME1 ;
  RECT 52.520 0.000 52.840 0.600 ;
 END
 ANTENNAPARTIALMETALAREA                  0.346 LAYER ME1 ;
 ANTENNAPARTIALMETALAREA                  1.466 LAYER ME2 ;
 ANTENNAPARTIALMETALAREA                  0.508 LAYER ME3 ;
 ANTENNAGATEAREA                          0.072 LAYER ME3 ;
 ANTENNAGATEAREA                          0.072 LAYER ME4 ;
 ANTENNADIFFAREA                          0.218 LAYER ME1 ;
 ANTENNADIFFAREA                          0.218 LAYER ME2 ;
 ANTENNADIFFAREA                          0.218 LAYER ME3 ;
 ANTENNADIFFAREA                          0.218 LAYER ME4 ;
 ANTENNAMAXAREACAR                       17.267 LAYER ME3 ;
 ANTENNAMAXAREACAR                       19.933 LAYER ME4 ;
END DI12
PIN DO12
  DIRECTION OUTPUT ;
 PORT
  LAYER ME4 ;
  RECT 53.082 0.000 53.402 0.600 ;
  LAYER ME3 ;
  RECT 53.082 0.000 53.402 0.600 ;
  LAYER ME2 ;
  RECT 53.082 0.000 53.402 0.600 ;
  LAYER ME1 ;
  RECT 53.082 0.000 53.402 0.600 ;
 END
 ANTENNAPARTIALMETALAREA                  5.602 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME3 ;
 ANTENNADIFFAREA                          1.293 LAYER ME4 ;
END DO12
PIN WEB1
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 51.080 0.000 51.400 0.600 ;
  LAYER ME3 ;
  RECT 51.080 0.000 51.400 0.600 ;
  LAYER ME2 ;
  RECT 51.080 0.000 51.400 0.600 ;
  LAYER ME1 ;
  RECT 51.080 0.000 51.400 0.600 ;
 END
 ANTENNAPARTIALMETALAREA                  1.036 LAYER ME2 ;
 ANTENNAGATEAREA                          0.288 LAYER ME2 ;
 ANTENNAGATEAREA                          0.288 LAYER ME3 ;
 ANTENNAGATEAREA                          0.288 LAYER ME4 ;
 ANTENNADIFFAREA                          0.206 LAYER ME2 ;
 ANTENNADIFFAREA                          0.206 LAYER ME3 ;
 ANTENNADIFFAREA                          0.206 LAYER ME4 ;
 ANTENNAMAXAREACAR                        5.844 LAYER ME2 ;
 ANTENNAMAXAREACAR                        6.511 LAYER ME3 ;
 ANTENNAMAXAREACAR                        7.178 LAYER ME4 ;
END WEB1
PIN DI11
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 49.078 0.000 49.398 0.600 ;
  LAYER ME3 ;
  RECT 49.078 0.000 49.398 0.600 ;
  LAYER ME2 ;
  RECT 49.078 0.000 49.398 0.600 ;
  LAYER ME1 ;
  RECT 49.078 0.000 49.398 0.600 ;
 END
 ANTENNAPARTIALMETALAREA                  1.058 LAYER ME2 ;
 ANTENNAGATEAREA                          0.072 LAYER ME2 ;
 ANTENNAGATEAREA                          0.072 LAYER ME3 ;
 ANTENNAGATEAREA                          0.072 LAYER ME4 ;
 ANTENNADIFFAREA                          0.160 LAYER ME2 ;
 ANTENNADIFFAREA                          0.160 LAYER ME3 ;
 ANTENNADIFFAREA                          0.160 LAYER ME4 ;
 ANTENNAMAXAREACAR                       21.782 LAYER ME2 ;
 ANTENNAMAXAREACAR                       24.449 LAYER ME3 ;
 ANTENNAMAXAREACAR                       27.116 LAYER ME4 ;
END DI11
PIN DO11
  DIRECTION OUTPUT ;
 PORT
  LAYER ME4 ;
  RECT 48.516 0.000 48.836 0.600 ;
  LAYER ME3 ;
  RECT 48.516 0.000 48.836 0.600 ;
  LAYER ME2 ;
  RECT 48.516 0.000 48.836 0.600 ;
  LAYER ME1 ;
  RECT 48.516 0.000 48.836 0.600 ;
 END
 ANTENNAPARTIALMETALAREA                  5.273 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME3 ;
 ANTENNADIFFAREA                          1.293 LAYER ME4 ;
END DO11
PIN DI10
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 45.074 0.000 45.394 0.600 ;
  LAYER ME3 ;
  RECT 45.074 0.000 45.394 0.600 ;
  LAYER ME2 ;
  RECT 45.074 0.000 45.394 0.600 ;
  LAYER ME1 ;
  RECT 45.074 0.000 45.394 0.600 ;
 END
 ANTENNAPARTIALMETALAREA                  1.058 LAYER ME2 ;
 ANTENNAGATEAREA                          0.072 LAYER ME2 ;
 ANTENNAGATEAREA                          0.072 LAYER ME3 ;
 ANTENNAGATEAREA                          0.072 LAYER ME4 ;
 ANTENNADIFFAREA                          0.160 LAYER ME2 ;
 ANTENNADIFFAREA                          0.160 LAYER ME3 ;
 ANTENNADIFFAREA                          0.160 LAYER ME4 ;
 ANTENNAMAXAREACAR                       21.782 LAYER ME2 ;
 ANTENNAMAXAREACAR                       24.449 LAYER ME3 ;
 ANTENNAMAXAREACAR                       27.116 LAYER ME4 ;
END DI10
PIN DO10
  DIRECTION OUTPUT ;
 PORT
  LAYER ME4 ;
  RECT 44.512 0.000 44.832 0.600 ;
  LAYER ME3 ;
  RECT 44.512 0.000 44.832 0.600 ;
  LAYER ME2 ;
  RECT 44.512 0.000 44.832 0.600 ;
  LAYER ME1 ;
  RECT 44.512 0.000 44.832 0.600 ;
 END
 ANTENNAPARTIALMETALAREA                  5.273 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME3 ;
 ANTENNADIFFAREA                          1.293 LAYER ME4 ;
END DO10
PIN DI9
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 41.070 0.000 41.390 0.600 ;
  LAYER ME3 ;
  RECT 41.070 0.000 41.390 0.600 ;
  LAYER ME2 ;
  RECT 41.070 0.000 41.390 0.600 ;
  LAYER ME1 ;
  RECT 41.070 0.000 41.390 0.600 ;
 END
 ANTENNAPARTIALMETALAREA                  1.058 LAYER ME2 ;
 ANTENNAGATEAREA                          0.072 LAYER ME2 ;
 ANTENNAGATEAREA                          0.072 LAYER ME3 ;
 ANTENNAGATEAREA                          0.072 LAYER ME4 ;
 ANTENNADIFFAREA                          0.160 LAYER ME2 ;
 ANTENNADIFFAREA                          0.160 LAYER ME3 ;
 ANTENNADIFFAREA                          0.160 LAYER ME4 ;
 ANTENNAMAXAREACAR                       21.782 LAYER ME2 ;
 ANTENNAMAXAREACAR                       24.449 LAYER ME3 ;
 ANTENNAMAXAREACAR                       27.116 LAYER ME4 ;
END DI9
PIN DO9
  DIRECTION OUTPUT ;
 PORT
  LAYER ME4 ;
  RECT 40.508 0.000 40.828 0.600 ;
  LAYER ME3 ;
  RECT 40.508 0.000 40.828 0.600 ;
  LAYER ME2 ;
  RECT 40.508 0.000 40.828 0.600 ;
  LAYER ME1 ;
  RECT 40.508 0.000 40.828 0.600 ;
 END
 ANTENNAPARTIALMETALAREA                  5.273 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME3 ;
 ANTENNADIFFAREA                          1.293 LAYER ME4 ;
END DO9
PIN DI8
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 37.066 0.000 37.386 0.600 ;
  LAYER ME3 ;
  RECT 37.066 0.000 37.386 0.600 ;
  LAYER ME2 ;
  RECT 37.066 0.000 37.386 0.600 ;
  LAYER ME1 ;
  RECT 37.066 0.000 37.386 0.600 ;
 END
 ANTENNAPARTIALMETALAREA                  1.058 LAYER ME2 ;
 ANTENNAGATEAREA                          0.072 LAYER ME2 ;
 ANTENNAGATEAREA                          0.072 LAYER ME3 ;
 ANTENNAGATEAREA                          0.072 LAYER ME4 ;
 ANTENNADIFFAREA                          0.160 LAYER ME2 ;
 ANTENNADIFFAREA                          0.160 LAYER ME3 ;
 ANTENNADIFFAREA                          0.160 LAYER ME4 ;
 ANTENNAMAXAREACAR                       21.782 LAYER ME2 ;
 ANTENNAMAXAREACAR                       24.449 LAYER ME3 ;
 ANTENNAMAXAREACAR                       27.116 LAYER ME4 ;
END DI8
PIN DO8
  DIRECTION OUTPUT ;
 PORT
  LAYER ME4 ;
  RECT 36.504 0.000 36.824 0.600 ;
  LAYER ME3 ;
  RECT 36.504 0.000 36.824 0.600 ;
  LAYER ME2 ;
  RECT 36.504 0.000 36.824 0.600 ;
  LAYER ME1 ;
  RECT 36.504 0.000 36.824 0.600 ;
 END
 ANTENNAPARTIALMETALAREA                  5.273 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME3 ;
 ANTENNADIFFAREA                          1.293 LAYER ME4 ;
END DO8
PIN DI7
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 33.062 0.000 33.382 0.600 ;
  LAYER ME3 ;
  RECT 33.062 0.000 33.382 0.600 ;
  LAYER ME2 ;
  RECT 33.062 0.000 33.382 0.600 ;
  LAYER ME1 ;
  RECT 33.062 0.000 33.382 0.600 ;
 END
 ANTENNAPARTIALMETALAREA                  1.058 LAYER ME2 ;
 ANTENNAGATEAREA                          0.072 LAYER ME2 ;
 ANTENNAGATEAREA                          0.072 LAYER ME3 ;
 ANTENNAGATEAREA                          0.072 LAYER ME4 ;
 ANTENNADIFFAREA                          0.160 LAYER ME2 ;
 ANTENNADIFFAREA                          0.160 LAYER ME3 ;
 ANTENNADIFFAREA                          0.160 LAYER ME4 ;
 ANTENNAMAXAREACAR                       21.782 LAYER ME2 ;
 ANTENNAMAXAREACAR                       24.449 LAYER ME3 ;
 ANTENNAMAXAREACAR                       27.116 LAYER ME4 ;
END DI7
PIN DO7
  DIRECTION OUTPUT ;
 PORT
  LAYER ME4 ;
  RECT 32.500 0.000 32.820 0.600 ;
  LAYER ME3 ;
  RECT 32.500 0.000 32.820 0.600 ;
  LAYER ME2 ;
  RECT 32.500 0.000 32.820 0.600 ;
  LAYER ME1 ;
  RECT 32.500 0.000 32.820 0.600 ;
 END
 ANTENNAPARTIALMETALAREA                  5.273 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME3 ;
 ANTENNADIFFAREA                          1.293 LAYER ME4 ;
END DO7
PIN DI6
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 29.058 0.000 29.378 0.600 ;
  LAYER ME3 ;
  RECT 29.058 0.000 29.378 0.600 ;
  LAYER ME2 ;
  RECT 29.058 0.000 29.378 0.600 ;
  LAYER ME1 ;
  RECT 29.058 0.000 29.378 0.600 ;
 END
 ANTENNAPARTIALMETALAREA                  1.058 LAYER ME2 ;
 ANTENNAGATEAREA                          0.072 LAYER ME2 ;
 ANTENNAGATEAREA                          0.072 LAYER ME3 ;
 ANTENNAGATEAREA                          0.072 LAYER ME4 ;
 ANTENNADIFFAREA                          0.160 LAYER ME2 ;
 ANTENNADIFFAREA                          0.160 LAYER ME3 ;
 ANTENNADIFFAREA                          0.160 LAYER ME4 ;
 ANTENNAMAXAREACAR                       21.782 LAYER ME2 ;
 ANTENNAMAXAREACAR                       24.449 LAYER ME3 ;
 ANTENNAMAXAREACAR                       27.116 LAYER ME4 ;
END DI6
PIN DO6
  DIRECTION OUTPUT ;
 PORT
  LAYER ME4 ;
  RECT 28.496 0.000 28.816 0.600 ;
  LAYER ME3 ;
  RECT 28.496 0.000 28.816 0.600 ;
  LAYER ME2 ;
  RECT 28.496 0.000 28.816 0.600 ;
  LAYER ME1 ;
  RECT 28.496 0.000 28.816 0.600 ;
 END
 ANTENNAPARTIALMETALAREA                  5.273 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME3 ;
 ANTENNADIFFAREA                          1.293 LAYER ME4 ;
END DO6
PIN DI5
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 25.054 0.000 25.374 0.600 ;
  LAYER ME3 ;
  RECT 25.054 0.000 25.374 0.600 ;
  LAYER ME2 ;
  RECT 25.054 0.000 25.374 0.600 ;
  LAYER ME1 ;
  RECT 25.054 0.000 25.374 0.600 ;
 END
 ANTENNAPARTIALMETALAREA                  1.058 LAYER ME2 ;
 ANTENNAGATEAREA                          0.072 LAYER ME2 ;
 ANTENNAGATEAREA                          0.072 LAYER ME3 ;
 ANTENNAGATEAREA                          0.072 LAYER ME4 ;
 ANTENNADIFFAREA                          0.160 LAYER ME2 ;
 ANTENNADIFFAREA                          0.160 LAYER ME3 ;
 ANTENNADIFFAREA                          0.160 LAYER ME4 ;
 ANTENNAMAXAREACAR                       21.782 LAYER ME2 ;
 ANTENNAMAXAREACAR                       24.449 LAYER ME3 ;
 ANTENNAMAXAREACAR                       27.116 LAYER ME4 ;
END DI5
PIN DO5
  DIRECTION OUTPUT ;
 PORT
  LAYER ME4 ;
  RECT 24.492 0.000 24.812 0.600 ;
  LAYER ME3 ;
  RECT 24.492 0.000 24.812 0.600 ;
  LAYER ME2 ;
  RECT 24.492 0.000 24.812 0.600 ;
  LAYER ME1 ;
  RECT 24.492 0.000 24.812 0.600 ;
 END
 ANTENNAPARTIALMETALAREA                  5.273 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME3 ;
 ANTENNADIFFAREA                          1.293 LAYER ME4 ;
END DO5
PIN DI4
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 21.050 0.000 21.370 0.600 ;
  LAYER ME3 ;
  RECT 21.050 0.000 21.370 0.600 ;
  LAYER ME2 ;
  RECT 21.050 0.000 21.370 0.600 ;
  LAYER ME1 ;
  RECT 21.050 0.000 21.370 0.600 ;
 END
 ANTENNAPARTIALMETALAREA                  1.058 LAYER ME2 ;
 ANTENNAGATEAREA                          0.072 LAYER ME2 ;
 ANTENNAGATEAREA                          0.072 LAYER ME3 ;
 ANTENNAGATEAREA                          0.072 LAYER ME4 ;
 ANTENNADIFFAREA                          0.160 LAYER ME2 ;
 ANTENNADIFFAREA                          0.160 LAYER ME3 ;
 ANTENNADIFFAREA                          0.160 LAYER ME4 ;
 ANTENNAMAXAREACAR                       21.782 LAYER ME2 ;
 ANTENNAMAXAREACAR                       24.449 LAYER ME3 ;
 ANTENNAMAXAREACAR                       27.116 LAYER ME4 ;
END DI4
PIN DO4
  DIRECTION OUTPUT ;
 PORT
  LAYER ME4 ;
  RECT 20.488 0.000 20.808 0.600 ;
  LAYER ME3 ;
  RECT 20.488 0.000 20.808 0.600 ;
  LAYER ME2 ;
  RECT 20.488 0.000 20.808 0.600 ;
  LAYER ME1 ;
  RECT 20.488 0.000 20.808 0.600 ;
 END
 ANTENNAPARTIALMETALAREA                  5.273 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME3 ;
 ANTENNADIFFAREA                          1.293 LAYER ME4 ;
END DO4
PIN DI3
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 17.046 0.000 17.366 0.600 ;
  LAYER ME3 ;
  RECT 17.046 0.000 17.366 0.600 ;
  LAYER ME2 ;
  RECT 17.046 0.000 17.366 0.600 ;
  LAYER ME1 ;
  RECT 17.046 0.000 17.366 0.600 ;
 END
 ANTENNAPARTIALMETALAREA                  1.058 LAYER ME2 ;
 ANTENNAGATEAREA                          0.072 LAYER ME2 ;
 ANTENNAGATEAREA                          0.072 LAYER ME3 ;
 ANTENNAGATEAREA                          0.072 LAYER ME4 ;
 ANTENNADIFFAREA                          0.160 LAYER ME2 ;
 ANTENNADIFFAREA                          0.160 LAYER ME3 ;
 ANTENNADIFFAREA                          0.160 LAYER ME4 ;
 ANTENNAMAXAREACAR                       21.782 LAYER ME2 ;
 ANTENNAMAXAREACAR                       24.449 LAYER ME3 ;
 ANTENNAMAXAREACAR                       27.116 LAYER ME4 ;
END DI3
PIN DO3
  DIRECTION OUTPUT ;
 PORT
  LAYER ME4 ;
  RECT 16.484 0.000 16.804 0.600 ;
  LAYER ME3 ;
  RECT 16.484 0.000 16.804 0.600 ;
  LAYER ME2 ;
  RECT 16.484 0.000 16.804 0.600 ;
  LAYER ME1 ;
  RECT 16.484 0.000 16.804 0.600 ;
 END
 ANTENNAPARTIALMETALAREA                  5.273 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME3 ;
 ANTENNADIFFAREA                          1.293 LAYER ME4 ;
END DO3
PIN DI2
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 13.042 0.000 13.362 0.600 ;
  LAYER ME3 ;
  RECT 13.042 0.000 13.362 0.600 ;
  LAYER ME2 ;
  RECT 13.042 0.000 13.362 0.600 ;
  LAYER ME1 ;
  RECT 13.042 0.000 13.362 0.600 ;
 END
 ANTENNAPARTIALMETALAREA                  1.058 LAYER ME2 ;
 ANTENNAGATEAREA                          0.072 LAYER ME2 ;
 ANTENNAGATEAREA                          0.072 LAYER ME3 ;
 ANTENNAGATEAREA                          0.072 LAYER ME4 ;
 ANTENNADIFFAREA                          0.160 LAYER ME2 ;
 ANTENNADIFFAREA                          0.160 LAYER ME3 ;
 ANTENNADIFFAREA                          0.160 LAYER ME4 ;
 ANTENNAMAXAREACAR                       21.782 LAYER ME2 ;
 ANTENNAMAXAREACAR                       24.449 LAYER ME3 ;
 ANTENNAMAXAREACAR                       27.116 LAYER ME4 ;
END DI2
PIN DO2
  DIRECTION OUTPUT ;
 PORT
  LAYER ME4 ;
  RECT 12.480 0.000 12.800 0.600 ;
  LAYER ME3 ;
  RECT 12.480 0.000 12.800 0.600 ;
  LAYER ME2 ;
  RECT 12.480 0.000 12.800 0.600 ;
  LAYER ME1 ;
  RECT 12.480 0.000 12.800 0.600 ;
 END
 ANTENNAPARTIALMETALAREA                  5.273 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME3 ;
 ANTENNADIFFAREA                          1.293 LAYER ME4 ;
END DO2
PIN DI1
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 9.038 0.000 9.358 0.600 ;
  LAYER ME3 ;
  RECT 9.038 0.000 9.358 0.600 ;
  LAYER ME2 ;
  RECT 9.038 0.000 9.358 0.600 ;
  LAYER ME1 ;
  RECT 9.038 0.000 9.358 0.600 ;
 END
 ANTENNAPARTIALMETALAREA                  1.058 LAYER ME2 ;
 ANTENNAGATEAREA                          0.072 LAYER ME2 ;
 ANTENNAGATEAREA                          0.072 LAYER ME3 ;
 ANTENNAGATEAREA                          0.072 LAYER ME4 ;
 ANTENNADIFFAREA                          0.160 LAYER ME2 ;
 ANTENNADIFFAREA                          0.160 LAYER ME3 ;
 ANTENNADIFFAREA                          0.160 LAYER ME4 ;
 ANTENNAMAXAREACAR                       21.782 LAYER ME2 ;
 ANTENNAMAXAREACAR                       24.449 LAYER ME3 ;
 ANTENNAMAXAREACAR                       27.116 LAYER ME4 ;
END DI1
PIN DO1
  DIRECTION OUTPUT ;
 PORT
  LAYER ME4 ;
  RECT 8.476 0.000 8.796 0.600 ;
  LAYER ME3 ;
  RECT 8.476 0.000 8.796 0.600 ;
  LAYER ME2 ;
  RECT 8.476 0.000 8.796 0.600 ;
  LAYER ME1 ;
  RECT 8.476 0.000 8.796 0.600 ;
 END
 ANTENNAPARTIALMETALAREA                  5.273 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME3 ;
 ANTENNADIFFAREA                          1.293 LAYER ME4 ;
END DO1
PIN DI0
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 4.472 0.000 4.792 0.600 ;
  LAYER ME3 ;
  RECT 4.472 0.000 4.792 0.600 ;
  LAYER ME2 ;
  RECT 4.472 0.000 4.792 0.600 ;
  LAYER ME1 ;
  RECT 4.472 0.000 4.792 0.600 ;
 END
 ANTENNAPARTIALMETALAREA                  0.346 LAYER ME1 ;
 ANTENNAPARTIALMETALAREA                  1.466 LAYER ME2 ;
 ANTENNAPARTIALMETALAREA                  0.508 LAYER ME3 ;
 ANTENNAGATEAREA                          0.072 LAYER ME3 ;
 ANTENNAGATEAREA                          0.072 LAYER ME4 ;
 ANTENNADIFFAREA                          0.218 LAYER ME1 ;
 ANTENNADIFFAREA                          0.218 LAYER ME2 ;
 ANTENNADIFFAREA                          0.218 LAYER ME3 ;
 ANTENNADIFFAREA                          0.218 LAYER ME4 ;
 ANTENNAMAXAREACAR                       17.267 LAYER ME3 ;
 ANTENNAMAXAREACAR                       19.933 LAYER ME4 ;
END DI0
PIN DO0
  DIRECTION OUTPUT ;
 PORT
  LAYER ME4 ;
  RECT 5.034 0.000 5.354 0.600 ;
  LAYER ME3 ;
  RECT 5.034 0.000 5.354 0.600 ;
  LAYER ME2 ;
  RECT 5.034 0.000 5.354 0.600 ;
  LAYER ME1 ;
  RECT 5.034 0.000 5.354 0.600 ;
 END
 ANTENNAPARTIALMETALAREA                  5.602 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME3 ;
 ANTENNADIFFAREA                          1.293 LAYER ME4 ;
END DO0
PIN WEB0
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 3.032 0.000 3.352 0.600 ;
  LAYER ME3 ;
  RECT 3.032 0.000 3.352 0.600 ;
  LAYER ME2 ;
  RECT 3.032 0.000 3.352 0.600 ;
  LAYER ME1 ;
  RECT 3.032 0.000 3.352 0.600 ;
 END
 ANTENNAPARTIALMETALAREA                  1.036 LAYER ME2 ;
 ANTENNAGATEAREA                          0.288 LAYER ME2 ;
 ANTENNAGATEAREA                          0.288 LAYER ME3 ;
 ANTENNAGATEAREA                          0.288 LAYER ME4 ;
 ANTENNADIFFAREA                          0.206 LAYER ME2 ;
 ANTENNADIFFAREA                          0.206 LAYER ME3 ;
 ANTENNADIFFAREA                          0.206 LAYER ME4 ;
 ANTENNAMAXAREACAR                        5.844 LAYER ME2 ;
 ANTENNAMAXAREACAR                        6.511 LAYER ME3 ;
 ANTENNAMAXAREACAR                        7.178 LAYER ME4 ;
END WEB0
PIN A1
  DIRECTION INPUT ;
 PORT
  LAYER ME3 ;
  RECT 211.072 0.000 211.392 0.720 ;
  LAYER ME2 ;
  RECT 211.072 0.000 211.392 0.720 ;
  LAYER ME1 ;
  RECT 211.072 0.000 211.392 0.720 ;
 END
 ANTENNAPARTIALMETALAREA                  3.547 LAYER ME2 ;
 ANTENNAGATEAREA                          0.144 LAYER ME2 ;
 ANTENNAGATEAREA                          0.144 LAYER ME3 ;
 ANTENNADIFFAREA                          0.218 LAYER ME2 ;
 ANTENNADIFFAREA                          0.218 LAYER ME3 ;
 ANTENNAMAXAREACAR                       27.235 LAYER ME2 ;
 ANTENNAMAXAREACAR                       28.835 LAYER ME3 ;
END A1
PIN A2
  DIRECTION INPUT ;
 PORT
  LAYER ME3 ;
  RECT 211.642 0.000 211.962 0.720 ;
  LAYER ME2 ;
  RECT 211.642 0.000 211.962 0.720 ;
  LAYER ME1 ;
  RECT 211.642 0.000 211.962 0.720 ;
 END
 ANTENNAPARTIALMETALAREA                  3.688 LAYER ME2 ;
 ANTENNAGATEAREA                          0.144 LAYER ME2 ;
 ANTENNAGATEAREA                          0.144 LAYER ME3 ;
 ANTENNADIFFAREA                          0.218 LAYER ME2 ;
 ANTENNADIFFAREA                          0.218 LAYER ME3 ;
 ANTENNAMAXAREACAR                       28.214 LAYER ME2 ;
 ANTENNAMAXAREACAR                       29.814 LAYER ME3 ;
END A2
PIN A3
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 204.824 0.000 205.144 0.720 ;
  LAYER ME3 ;
  RECT 204.824 0.000 205.144 0.720 ;
  LAYER ME2 ;
  RECT 204.824 0.000 205.144 0.720 ;
  LAYER ME1 ;
  RECT 204.824 0.000 205.144 0.720 ;
 END
 ANTENNAPARTIALMETALAREA                  4.391 LAYER ME2 ;
 ANTENNAGATEAREA                          0.180 LAYER ME2 ;
 ANTENNAGATEAREA                          0.180 LAYER ME3 ;
 ANTENNAGATEAREA                          0.180 LAYER ME4 ;
 ANTENNADIFFAREA                          0.218 LAYER ME2 ;
 ANTENNADIFFAREA                          0.218 LAYER ME3 ;
 ANTENNADIFFAREA                          0.218 LAYER ME4 ;
 ANTENNAMAXAREACAR                       27.451 LAYER ME2 ;
 ANTENNAMAXAREACAR                       28.731 LAYER ME3 ;
 ANTENNAMAXAREACAR                       30.011 LAYER ME4 ;
END A3
PIN A4
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 204.144 0.000 204.464 0.720 ;
  LAYER ME3 ;
  RECT 204.144 0.000 204.464 0.720 ;
  LAYER ME2 ;
  RECT 204.144 0.000 204.464 0.720 ;
  LAYER ME1 ;
  RECT 204.144 0.000 204.464 0.720 ;
 END
 ANTENNAPARTIALMETALAREA                  3.928 LAYER ME2 ;
 ANTENNAGATEAREA                          0.180 LAYER ME2 ;
 ANTENNAGATEAREA                          0.180 LAYER ME3 ;
 ANTENNAGATEAREA                          0.180 LAYER ME4 ;
 ANTENNADIFFAREA                          0.218 LAYER ME2 ;
 ANTENNADIFFAREA                          0.218 LAYER ME3 ;
 ANTENNADIFFAREA                          0.218 LAYER ME4 ;
 ANTENNAMAXAREACAR                       26.813 LAYER ME2 ;
 ANTENNAMAXAREACAR                       28.093 LAYER ME3 ;
 ANTENNAMAXAREACAR                       29.373 LAYER ME4 ;
END A4
PIN A5
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 200.704 0.000 200.984 0.720 ;
  LAYER ME3 ;
  RECT 200.704 0.000 200.984 0.720 ;
  LAYER ME2 ;
  RECT 200.704 0.000 200.984 0.720 ;
  LAYER ME1 ;
  RECT 200.704 0.000 200.984 0.720 ;
 END
 ANTENNAPARTIALMETALAREA                  4.391 LAYER ME2 ;
 ANTENNAGATEAREA                          0.180 LAYER ME2 ;
 ANTENNAGATEAREA                          0.180 LAYER ME3 ;
 ANTENNAGATEAREA                          0.180 LAYER ME4 ;
 ANTENNADIFFAREA                          0.218 LAYER ME2 ;
 ANTENNADIFFAREA                          0.218 LAYER ME3 ;
 ANTENNADIFFAREA                          0.218 LAYER ME4 ;
 ANTENNAMAXAREACAR                       27.291 LAYER ME2 ;
 ANTENNAMAXAREACAR                       28.411 LAYER ME3 ;
 ANTENNAMAXAREACAR                       29.531 LAYER ME4 ;
END A5
PIN A0
  DIRECTION INPUT ;
 PORT
  LAYER ME3 ;
  RECT 221.658 0.000 221.978 0.662 ;
  LAYER ME2 ;
  RECT 221.658 0.000 221.978 0.662 ;
  LAYER ME1 ;
  RECT 221.658 0.000 221.978 0.662 ;
 END
 ANTENNAPARTIALMETALAREA                  5.907 LAYER ME2 ;
 ANTENNAGATEAREA                          0.108 LAYER ME2 ;
 ANTENNAGATEAREA                          0.108 LAYER ME3 ;
 ANTENNADIFFAREA                          0.218 LAYER ME2 ;
 ANTENNADIFFAREA                          0.218 LAYER ME3 ;
 ANTENNAMAXAREACAR                       58.521 LAYER ME2 ;
 ANTENNAMAXAREACAR                       60.482 LAYER ME3 ;
END A0
PIN DVSE
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 231.249 0.000 231.569 0.720 ;
  LAYER ME3 ;
  RECT 231.249 0.000 231.569 0.720 ;
  LAYER ME3 ;
  RECT 231.249 0.000 231.569 0.720 ;
  LAYER ME2 ;
  RECT 231.249 0.000 231.569 0.720 ;
  LAYER ME2 ;
  RECT 231.249 0.000 231.569 0.720 ;
  LAYER ME1 ;
  RECT 231.249 0.000 231.569 0.720 ;
  LAYER ME1 ;
  RECT 231.249 0.000 231.569 0.720 ;
 END
 ANTENNAPARTIALMETALAREA                  7.809 LAYER ME2 ;
 ANTENNAGATEAREA                          0.612 LAYER ME2 ;
 ANTENNAGATEAREA                          0.612 LAYER ME3 ;
 ANTENNAGATEAREA                          0.612 LAYER ME4 ;
 ANTENNADIFFAREA                          0.218 LAYER ME2 ;
 ANTENNADIFFAREA                          0.218 LAYER ME3 ;
 ANTENNADIFFAREA                          0.218 LAYER ME4 ;
 ANTENNAMAXAREACAR                       76.330 LAYER ME2 ;
 ANTENNAMAXAREACAR                       78.463 LAYER ME3 ;
 ANTENNAMAXAREACAR                       80.596 LAYER ME4 ;
END DVSE
PIN DVS3
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 230.729 0.000 231.049 0.720 ;
  LAYER ME3 ;
  RECT 230.729 0.000 231.049 0.720 ;
  LAYER ME3 ;
  RECT 230.729 0.000 231.049 0.720 ;
  LAYER ME2 ;
  RECT 230.729 0.000 231.049 0.720 ;
  LAYER ME2 ;
  RECT 230.729 0.000 231.049 0.720 ;
  LAYER ME1 ;
  RECT 230.729 0.000 231.049 0.720 ;
  LAYER ME1 ;
  RECT 230.729 0.000 231.049 0.720 ;
 END
 ANTENNAPARTIALMETALAREA                  6.179 LAYER ME2 ;
 ANTENNAGATEAREA                          0.108 LAYER ME2 ;
 ANTENNAGATEAREA                          0.108 LAYER ME3 ;
 ANTENNAGATEAREA                          0.108 LAYER ME4 ;
 ANTENNADIFFAREA                          0.218 LAYER ME2 ;
 ANTENNADIFFAREA                          0.218 LAYER ME3 ;
 ANTENNADIFFAREA                          0.218 LAYER ME4 ;
 ANTENNAMAXAREACAR                       68.823 LAYER ME2 ;
 ANTENNAMAXAREACAR                       70.956 LAYER ME3 ;
 ANTENNAMAXAREACAR                       73.089 LAYER ME4 ;
END DVS3
PIN DVS2
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 231.769 0.000 232.089 0.720 ;
  LAYER ME3 ;
  RECT 231.769 0.000 232.089 0.720 ;
  LAYER ME3 ;
  RECT 231.769 0.000 232.089 0.720 ;
  LAYER ME2 ;
  RECT 231.769 0.000 232.089 0.720 ;
  LAYER ME2 ;
  RECT 231.769 0.000 232.089 0.720 ;
  LAYER ME1 ;
  RECT 231.769 0.000 232.089 0.720 ;
  LAYER ME1 ;
  RECT 231.769 0.000 232.089 0.720 ;
 END
 ANTENNAPARTIALMETALAREA                  7.876 LAYER ME2 ;
 ANTENNAGATEAREA                          0.108 LAYER ME2 ;
 ANTENNAGATEAREA                          0.108 LAYER ME3 ;
 ANTENNAGATEAREA                          0.108 LAYER ME4 ;
 ANTENNADIFFAREA                          0.218 LAYER ME2 ;
 ANTENNADIFFAREA                          0.218 LAYER ME3 ;
 ANTENNADIFFAREA                          0.218 LAYER ME4 ;
 ANTENNAMAXAREACAR                       83.257 LAYER ME2 ;
 ANTENNAMAXAREACAR                       85.391 LAYER ME3 ;
 ANTENNAMAXAREACAR                       87.524 LAYER ME4 ;
END DVS2
PIN DVS1
  DIRECTION INPUT ;
 PORT
  LAYER ME3 ;
  RECT 228.113 0.000 228.433 0.720 ;
  LAYER ME2 ;
  RECT 228.113 0.000 228.433 0.720 ;
  LAYER ME1 ;
  RECT 228.113 0.000 228.433 0.720 ;
 END
 ANTENNAPARTIALMETALAREA                  6.247 LAYER ME2 ;
 ANTENNAGATEAREA                          0.108 LAYER ME2 ;
 ANTENNAGATEAREA                          0.108 LAYER ME3 ;
 ANTENNADIFFAREA                          0.218 LAYER ME2 ;
 ANTENNADIFFAREA                          0.218 LAYER ME3 ;
 ANTENNAMAXAREACAR                       69.294 LAYER ME2 ;
 ANTENNAMAXAREACAR                       71.427 LAYER ME3 ;
END DVS1
PIN DVS0
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 232.289 0.000 232.609 0.720 ;
  LAYER ME3 ;
  RECT 232.289 0.000 232.609 0.720 ;
  LAYER ME3 ;
  RECT 232.289 0.000 232.609 0.720 ;
  LAYER ME2 ;
  RECT 232.289 0.000 232.609 0.720 ;
  LAYER ME2 ;
  RECT 232.289 0.000 232.609 0.720 ;
  LAYER ME1 ;
  RECT 232.289 0.000 232.609 0.720 ;
  LAYER ME1 ;
  RECT 232.289 0.000 232.609 0.720 ;
 END
 ANTENNAPARTIALMETALAREA                  7.119 LAYER ME2 ;
 ANTENNAGATEAREA                          0.108 LAYER ME2 ;
 ANTENNAGATEAREA                          0.108 LAYER ME3 ;
 ANTENNAGATEAREA                          0.108 LAYER ME4 ;
 ANTENNADIFFAREA                          0.218 LAYER ME2 ;
 ANTENNADIFFAREA                          0.218 LAYER ME3 ;
 ANTENNADIFFAREA                          0.218 LAYER ME4 ;
 ANTENNAMAXAREACAR                       77.987 LAYER ME2 ;
 ANTENNAMAXAREACAR                       80.120 LAYER ME3 ;
 ANTENNAMAXAREACAR                       82.254 LAYER ME4 ;
END DVS0
PIN CK
  DIRECTION INPUT ;
 PORT
  LAYER ME3 ;
  RECT 224.197 0.000 224.517 0.720 ;
  LAYER ME2 ;
  RECT 224.197 0.000 224.517 0.720 ;
  LAYER ME1 ;
  RECT 224.197 0.000 224.517 0.720 ;
 END
 ANTENNAPARTIALMETALAREA                  5.257 LAYER ME2 ;
 ANTENNAPARTIALMETALAREA                  7.044 LAYER ME3 ;
 ANTENNAGATEAREA                          0.072 LAYER ME2 ;
 ANTENNAGATEAREA                          1.044 LAYER ME3 ;
 ANTENNADIFFAREA                          0.218 LAYER ME2 ;
 ANTENNADIFFAREA                          0.218 LAYER ME3 ;
 ANTENNAMAXAREACAR                       86.308 LAYER ME2 ;
 ANTENNAMAXAREACAR                      187.347 LAYER ME3 ;
END CK
PIN CSB
  DIRECTION INPUT ;
 PORT
  LAYER ME3 ;
  RECT 215.583 0.000 215.903 0.720 ;
  LAYER ME2 ;
  RECT 215.583 0.000 215.903 0.720 ;
  LAYER ME1 ;
  RECT 215.583 0.000 215.903 0.720 ;
 END
 ANTENNAPARTIALMETALAREA                  5.788 LAYER ME2 ;
 ANTENNAPARTIALMETALAREA                  7.100 LAYER ME3 ;
 ANTENNAGATEAREA                          2.508 LAYER ME2 ;
 ANTENNAGATEAREA                          3.480 LAYER ME3 ;
 ANTENNADIFFAREA                          0.218 LAYER ME2 ;
 ANTENNADIFFAREA                          0.218 LAYER ME3 ;
 ANTENNAMAXAREACAR                        3.046 LAYER ME2 ;
 ANTENNAMAXAREACAR                       36.487 LAYER ME3 ;
END CSB
PIN DI95
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 423.091 0.000 423.411 0.600 ;
  LAYER ME3 ;
  RECT 423.091 0.000 423.411 0.600 ;
  LAYER ME2 ;
  RECT 423.091 0.000 423.411 0.600 ;
  LAYER ME1 ;
  RECT 423.091 0.000 423.411 0.600 ;
 END
 ANTENNAPARTIALMETALAREA                  1.058 LAYER ME2 ;
 ANTENNAGATEAREA                          0.072 LAYER ME2 ;
 ANTENNAGATEAREA                          0.072 LAYER ME3 ;
 ANTENNAGATEAREA                          0.072 LAYER ME4 ;
 ANTENNADIFFAREA                          0.160 LAYER ME2 ;
 ANTENNADIFFAREA                          0.160 LAYER ME3 ;
 ANTENNADIFFAREA                          0.160 LAYER ME4 ;
 ANTENNAMAXAREACAR                       21.782 LAYER ME2 ;
 ANTENNAMAXAREACAR                       24.449 LAYER ME3 ;
 ANTENNAMAXAREACAR                       27.116 LAYER ME4 ;
END DI95
PIN DO95
  DIRECTION OUTPUT ;
 PORT
  LAYER ME4 ;
  RECT 422.529 0.000 422.849 0.600 ;
  LAYER ME3 ;
  RECT 422.529 0.000 422.849 0.600 ;
  LAYER ME2 ;
  RECT 422.529 0.000 422.849 0.600 ;
  LAYER ME1 ;
  RECT 422.529 0.000 422.849 0.600 ;
 END
 ANTENNAPARTIALMETALAREA                  5.273 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME3 ;
 ANTENNADIFFAREA                          1.293 LAYER ME4 ;
END DO95
PIN DI94
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 419.087 0.000 419.407 0.600 ;
  LAYER ME3 ;
  RECT 419.087 0.000 419.407 0.600 ;
  LAYER ME2 ;
  RECT 419.087 0.000 419.407 0.600 ;
  LAYER ME1 ;
  RECT 419.087 0.000 419.407 0.600 ;
 END
 ANTENNAPARTIALMETALAREA                  1.058 LAYER ME2 ;
 ANTENNAGATEAREA                          0.072 LAYER ME2 ;
 ANTENNAGATEAREA                          0.072 LAYER ME3 ;
 ANTENNAGATEAREA                          0.072 LAYER ME4 ;
 ANTENNADIFFAREA                          0.160 LAYER ME2 ;
 ANTENNADIFFAREA                          0.160 LAYER ME3 ;
 ANTENNADIFFAREA                          0.160 LAYER ME4 ;
 ANTENNAMAXAREACAR                       21.782 LAYER ME2 ;
 ANTENNAMAXAREACAR                       24.449 LAYER ME3 ;
 ANTENNAMAXAREACAR                       27.116 LAYER ME4 ;
END DI94
PIN DO94
  DIRECTION OUTPUT ;
 PORT
  LAYER ME4 ;
  RECT 418.525 0.000 418.845 0.600 ;
  LAYER ME3 ;
  RECT 418.525 0.000 418.845 0.600 ;
  LAYER ME2 ;
  RECT 418.525 0.000 418.845 0.600 ;
  LAYER ME1 ;
  RECT 418.525 0.000 418.845 0.600 ;
 END
 ANTENNAPARTIALMETALAREA                  5.273 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME3 ;
 ANTENNADIFFAREA                          1.293 LAYER ME4 ;
END DO94
PIN DI93
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 415.083 0.000 415.403 0.600 ;
  LAYER ME3 ;
  RECT 415.083 0.000 415.403 0.600 ;
  LAYER ME2 ;
  RECT 415.083 0.000 415.403 0.600 ;
  LAYER ME1 ;
  RECT 415.083 0.000 415.403 0.600 ;
 END
 ANTENNAPARTIALMETALAREA                  1.058 LAYER ME2 ;
 ANTENNAGATEAREA                          0.072 LAYER ME2 ;
 ANTENNAGATEAREA                          0.072 LAYER ME3 ;
 ANTENNAGATEAREA                          0.072 LAYER ME4 ;
 ANTENNADIFFAREA                          0.160 LAYER ME2 ;
 ANTENNADIFFAREA                          0.160 LAYER ME3 ;
 ANTENNADIFFAREA                          0.160 LAYER ME4 ;
 ANTENNAMAXAREACAR                       21.782 LAYER ME2 ;
 ANTENNAMAXAREACAR                       24.449 LAYER ME3 ;
 ANTENNAMAXAREACAR                       27.116 LAYER ME4 ;
END DI93
PIN DO93
  DIRECTION OUTPUT ;
 PORT
  LAYER ME4 ;
  RECT 414.521 0.000 414.841 0.600 ;
  LAYER ME3 ;
  RECT 414.521 0.000 414.841 0.600 ;
  LAYER ME2 ;
  RECT 414.521 0.000 414.841 0.600 ;
  LAYER ME1 ;
  RECT 414.521 0.000 414.841 0.600 ;
 END
 ANTENNAPARTIALMETALAREA                  5.273 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME3 ;
 ANTENNADIFFAREA                          1.293 LAYER ME4 ;
END DO93
PIN DI92
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 411.079 0.000 411.399 0.600 ;
  LAYER ME3 ;
  RECT 411.079 0.000 411.399 0.600 ;
  LAYER ME2 ;
  RECT 411.079 0.000 411.399 0.600 ;
  LAYER ME1 ;
  RECT 411.079 0.000 411.399 0.600 ;
 END
 ANTENNAPARTIALMETALAREA                  1.058 LAYER ME2 ;
 ANTENNAGATEAREA                          0.072 LAYER ME2 ;
 ANTENNAGATEAREA                          0.072 LAYER ME3 ;
 ANTENNAGATEAREA                          0.072 LAYER ME4 ;
 ANTENNADIFFAREA                          0.160 LAYER ME2 ;
 ANTENNADIFFAREA                          0.160 LAYER ME3 ;
 ANTENNADIFFAREA                          0.160 LAYER ME4 ;
 ANTENNAMAXAREACAR                       21.782 LAYER ME2 ;
 ANTENNAMAXAREACAR                       24.449 LAYER ME3 ;
 ANTENNAMAXAREACAR                       27.116 LAYER ME4 ;
END DI92
PIN DO92
  DIRECTION OUTPUT ;
 PORT
  LAYER ME4 ;
  RECT 410.517 0.000 410.837 0.600 ;
  LAYER ME3 ;
  RECT 410.517 0.000 410.837 0.600 ;
  LAYER ME2 ;
  RECT 410.517 0.000 410.837 0.600 ;
  LAYER ME1 ;
  RECT 410.517 0.000 410.837 0.600 ;
 END
 ANTENNAPARTIALMETALAREA                  5.273 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME3 ;
 ANTENNADIFFAREA                          1.293 LAYER ME4 ;
END DO92
PIN DI91
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 407.075 0.000 407.395 0.600 ;
  LAYER ME3 ;
  RECT 407.075 0.000 407.395 0.600 ;
  LAYER ME2 ;
  RECT 407.075 0.000 407.395 0.600 ;
  LAYER ME1 ;
  RECT 407.075 0.000 407.395 0.600 ;
 END
 ANTENNAPARTIALMETALAREA                  1.058 LAYER ME2 ;
 ANTENNAGATEAREA                          0.072 LAYER ME2 ;
 ANTENNAGATEAREA                          0.072 LAYER ME3 ;
 ANTENNAGATEAREA                          0.072 LAYER ME4 ;
 ANTENNADIFFAREA                          0.160 LAYER ME2 ;
 ANTENNADIFFAREA                          0.160 LAYER ME3 ;
 ANTENNADIFFAREA                          0.160 LAYER ME4 ;
 ANTENNAMAXAREACAR                       21.782 LAYER ME2 ;
 ANTENNAMAXAREACAR                       24.449 LAYER ME3 ;
 ANTENNAMAXAREACAR                       27.116 LAYER ME4 ;
END DI91
PIN DO91
  DIRECTION OUTPUT ;
 PORT
  LAYER ME4 ;
  RECT 406.513 0.000 406.833 0.600 ;
  LAYER ME3 ;
  RECT 406.513 0.000 406.833 0.600 ;
  LAYER ME2 ;
  RECT 406.513 0.000 406.833 0.600 ;
  LAYER ME1 ;
  RECT 406.513 0.000 406.833 0.600 ;
 END
 ANTENNAPARTIALMETALAREA                  5.273 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME3 ;
 ANTENNADIFFAREA                          1.293 LAYER ME4 ;
END DO91
PIN DI90
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 403.071 0.000 403.391 0.600 ;
  LAYER ME3 ;
  RECT 403.071 0.000 403.391 0.600 ;
  LAYER ME2 ;
  RECT 403.071 0.000 403.391 0.600 ;
  LAYER ME1 ;
  RECT 403.071 0.000 403.391 0.600 ;
 END
 ANTENNAPARTIALMETALAREA                  1.058 LAYER ME2 ;
 ANTENNAGATEAREA                          0.072 LAYER ME2 ;
 ANTENNAGATEAREA                          0.072 LAYER ME3 ;
 ANTENNAGATEAREA                          0.072 LAYER ME4 ;
 ANTENNADIFFAREA                          0.160 LAYER ME2 ;
 ANTENNADIFFAREA                          0.160 LAYER ME3 ;
 ANTENNADIFFAREA                          0.160 LAYER ME4 ;
 ANTENNAMAXAREACAR                       21.782 LAYER ME2 ;
 ANTENNAMAXAREACAR                       24.449 LAYER ME3 ;
 ANTENNAMAXAREACAR                       27.116 LAYER ME4 ;
END DI90
PIN DO90
  DIRECTION OUTPUT ;
 PORT
  LAYER ME4 ;
  RECT 402.509 0.000 402.829 0.600 ;
  LAYER ME3 ;
  RECT 402.509 0.000 402.829 0.600 ;
  LAYER ME2 ;
  RECT 402.509 0.000 402.829 0.600 ;
  LAYER ME1 ;
  RECT 402.509 0.000 402.829 0.600 ;
 END
 ANTENNAPARTIALMETALAREA                  5.273 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME3 ;
 ANTENNADIFFAREA                          1.293 LAYER ME4 ;
END DO90
PIN DI89
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 399.067 0.000 399.387 0.600 ;
  LAYER ME3 ;
  RECT 399.067 0.000 399.387 0.600 ;
  LAYER ME2 ;
  RECT 399.067 0.000 399.387 0.600 ;
  LAYER ME1 ;
  RECT 399.067 0.000 399.387 0.600 ;
 END
 ANTENNAPARTIALMETALAREA                  1.058 LAYER ME2 ;
 ANTENNAGATEAREA                          0.072 LAYER ME2 ;
 ANTENNAGATEAREA                          0.072 LAYER ME3 ;
 ANTENNAGATEAREA                          0.072 LAYER ME4 ;
 ANTENNADIFFAREA                          0.160 LAYER ME2 ;
 ANTENNADIFFAREA                          0.160 LAYER ME3 ;
 ANTENNADIFFAREA                          0.160 LAYER ME4 ;
 ANTENNAMAXAREACAR                       21.782 LAYER ME2 ;
 ANTENNAMAXAREACAR                       24.449 LAYER ME3 ;
 ANTENNAMAXAREACAR                       27.116 LAYER ME4 ;
END DI89
PIN DO89
  DIRECTION OUTPUT ;
 PORT
  LAYER ME4 ;
  RECT 398.505 0.000 398.825 0.600 ;
  LAYER ME3 ;
  RECT 398.505 0.000 398.825 0.600 ;
  LAYER ME2 ;
  RECT 398.505 0.000 398.825 0.600 ;
  LAYER ME1 ;
  RECT 398.505 0.000 398.825 0.600 ;
 END
 ANTENNAPARTIALMETALAREA                  5.273 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME3 ;
 ANTENNADIFFAREA                          1.293 LAYER ME4 ;
END DO89
PIN DI88
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 395.063 0.000 395.383 0.600 ;
  LAYER ME3 ;
  RECT 395.063 0.000 395.383 0.600 ;
  LAYER ME2 ;
  RECT 395.063 0.000 395.383 0.600 ;
  LAYER ME1 ;
  RECT 395.063 0.000 395.383 0.600 ;
 END
 ANTENNAPARTIALMETALAREA                  1.058 LAYER ME2 ;
 ANTENNAGATEAREA                          0.072 LAYER ME2 ;
 ANTENNAGATEAREA                          0.072 LAYER ME3 ;
 ANTENNAGATEAREA                          0.072 LAYER ME4 ;
 ANTENNADIFFAREA                          0.160 LAYER ME2 ;
 ANTENNADIFFAREA                          0.160 LAYER ME3 ;
 ANTENNADIFFAREA                          0.160 LAYER ME4 ;
 ANTENNAMAXAREACAR                       21.782 LAYER ME2 ;
 ANTENNAMAXAREACAR                       24.449 LAYER ME3 ;
 ANTENNAMAXAREACAR                       27.116 LAYER ME4 ;
END DI88
PIN DO88
  DIRECTION OUTPUT ;
 PORT
  LAYER ME4 ;
  RECT 394.501 0.000 394.821 0.600 ;
  LAYER ME3 ;
  RECT 394.501 0.000 394.821 0.600 ;
  LAYER ME2 ;
  RECT 394.501 0.000 394.821 0.600 ;
  LAYER ME1 ;
  RECT 394.501 0.000 394.821 0.600 ;
 END
 ANTENNAPARTIALMETALAREA                  5.273 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME3 ;
 ANTENNADIFFAREA                          1.293 LAYER ME4 ;
END DO88
PIN DI87
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 391.059 0.000 391.379 0.600 ;
  LAYER ME3 ;
  RECT 391.059 0.000 391.379 0.600 ;
  LAYER ME2 ;
  RECT 391.059 0.000 391.379 0.600 ;
  LAYER ME1 ;
  RECT 391.059 0.000 391.379 0.600 ;
 END
 ANTENNAPARTIALMETALAREA                  1.058 LAYER ME2 ;
 ANTENNAGATEAREA                          0.072 LAYER ME2 ;
 ANTENNAGATEAREA                          0.072 LAYER ME3 ;
 ANTENNAGATEAREA                          0.072 LAYER ME4 ;
 ANTENNADIFFAREA                          0.160 LAYER ME2 ;
 ANTENNADIFFAREA                          0.160 LAYER ME3 ;
 ANTENNADIFFAREA                          0.160 LAYER ME4 ;
 ANTENNAMAXAREACAR                       21.782 LAYER ME2 ;
 ANTENNAMAXAREACAR                       24.449 LAYER ME3 ;
 ANTENNAMAXAREACAR                       27.116 LAYER ME4 ;
END DI87
PIN DO87
  DIRECTION OUTPUT ;
 PORT
  LAYER ME4 ;
  RECT 390.497 0.000 390.817 0.600 ;
  LAYER ME3 ;
  RECT 390.497 0.000 390.817 0.600 ;
  LAYER ME2 ;
  RECT 390.497 0.000 390.817 0.600 ;
  LAYER ME1 ;
  RECT 390.497 0.000 390.817 0.600 ;
 END
 ANTENNAPARTIALMETALAREA                  5.273 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME3 ;
 ANTENNADIFFAREA                          1.293 LAYER ME4 ;
END DO87
PIN DI86
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 387.055 0.000 387.375 0.600 ;
  LAYER ME3 ;
  RECT 387.055 0.000 387.375 0.600 ;
  LAYER ME2 ;
  RECT 387.055 0.000 387.375 0.600 ;
  LAYER ME1 ;
  RECT 387.055 0.000 387.375 0.600 ;
 END
 ANTENNAPARTIALMETALAREA                  1.058 LAYER ME2 ;
 ANTENNAGATEAREA                          0.072 LAYER ME2 ;
 ANTENNAGATEAREA                          0.072 LAYER ME3 ;
 ANTENNAGATEAREA                          0.072 LAYER ME4 ;
 ANTENNADIFFAREA                          0.160 LAYER ME2 ;
 ANTENNADIFFAREA                          0.160 LAYER ME3 ;
 ANTENNADIFFAREA                          0.160 LAYER ME4 ;
 ANTENNAMAXAREACAR                       21.782 LAYER ME2 ;
 ANTENNAMAXAREACAR                       24.449 LAYER ME3 ;
 ANTENNAMAXAREACAR                       27.116 LAYER ME4 ;
END DI86
PIN DO86
  DIRECTION OUTPUT ;
 PORT
  LAYER ME4 ;
  RECT 386.493 0.000 386.813 0.600 ;
  LAYER ME3 ;
  RECT 386.493 0.000 386.813 0.600 ;
  LAYER ME2 ;
  RECT 386.493 0.000 386.813 0.600 ;
  LAYER ME1 ;
  RECT 386.493 0.000 386.813 0.600 ;
 END
 ANTENNAPARTIALMETALAREA                  5.273 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME3 ;
 ANTENNADIFFAREA                          1.293 LAYER ME4 ;
END DO86
PIN DI85
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 383.051 0.000 383.371 0.600 ;
  LAYER ME3 ;
  RECT 383.051 0.000 383.371 0.600 ;
  LAYER ME2 ;
  RECT 383.051 0.000 383.371 0.600 ;
  LAYER ME1 ;
  RECT 383.051 0.000 383.371 0.600 ;
 END
 ANTENNAPARTIALMETALAREA                  1.058 LAYER ME2 ;
 ANTENNAGATEAREA                          0.072 LAYER ME2 ;
 ANTENNAGATEAREA                          0.072 LAYER ME3 ;
 ANTENNAGATEAREA                          0.072 LAYER ME4 ;
 ANTENNADIFFAREA                          0.160 LAYER ME2 ;
 ANTENNADIFFAREA                          0.160 LAYER ME3 ;
 ANTENNADIFFAREA                          0.160 LAYER ME4 ;
 ANTENNAMAXAREACAR                       21.782 LAYER ME2 ;
 ANTENNAMAXAREACAR                       24.449 LAYER ME3 ;
 ANTENNAMAXAREACAR                       27.116 LAYER ME4 ;
END DI85
PIN DO85
  DIRECTION OUTPUT ;
 PORT
  LAYER ME4 ;
  RECT 382.489 0.000 382.809 0.600 ;
  LAYER ME3 ;
  RECT 382.489 0.000 382.809 0.600 ;
  LAYER ME2 ;
  RECT 382.489 0.000 382.809 0.600 ;
  LAYER ME1 ;
  RECT 382.489 0.000 382.809 0.600 ;
 END
 ANTENNAPARTIALMETALAREA                  5.273 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME3 ;
 ANTENNADIFFAREA                          1.293 LAYER ME4 ;
END DO85
PIN DI84
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 378.485 0.000 378.805 0.600 ;
  LAYER ME3 ;
  RECT 378.485 0.000 378.805 0.600 ;
  LAYER ME2 ;
  RECT 378.485 0.000 378.805 0.600 ;
  LAYER ME1 ;
  RECT 378.485 0.000 378.805 0.600 ;
 END
 ANTENNAPARTIALMETALAREA                  0.346 LAYER ME1 ;
 ANTENNAPARTIALMETALAREA                  1.466 LAYER ME2 ;
 ANTENNAPARTIALMETALAREA                  0.508 LAYER ME3 ;
 ANTENNAGATEAREA                          0.072 LAYER ME3 ;
 ANTENNAGATEAREA                          0.072 LAYER ME4 ;
 ANTENNADIFFAREA                          0.218 LAYER ME1 ;
 ANTENNADIFFAREA                          0.218 LAYER ME2 ;
 ANTENNADIFFAREA                          0.218 LAYER ME3 ;
 ANTENNADIFFAREA                          0.218 LAYER ME4 ;
 ANTENNAMAXAREACAR                       17.267 LAYER ME3 ;
 ANTENNAMAXAREACAR                       19.933 LAYER ME4 ;
END DI84
PIN DO84
  DIRECTION OUTPUT ;
 PORT
  LAYER ME4 ;
  RECT 379.047 0.000 379.367 0.600 ;
  LAYER ME3 ;
  RECT 379.047 0.000 379.367 0.600 ;
  LAYER ME2 ;
  RECT 379.047 0.000 379.367 0.600 ;
  LAYER ME1 ;
  RECT 379.047 0.000 379.367 0.600 ;
 END
 ANTENNAPARTIALMETALAREA                  5.602 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME3 ;
 ANTENNADIFFAREA                          1.293 LAYER ME4 ;
END DO84
PIN WEB7
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 377.045 0.000 377.365 0.600 ;
  LAYER ME3 ;
  RECT 377.045 0.000 377.365 0.600 ;
  LAYER ME2 ;
  RECT 377.045 0.000 377.365 0.600 ;
  LAYER ME1 ;
  RECT 377.045 0.000 377.365 0.600 ;
 END
 ANTENNAPARTIALMETALAREA                  1.036 LAYER ME2 ;
 ANTENNAGATEAREA                          0.288 LAYER ME2 ;
 ANTENNAGATEAREA                          0.288 LAYER ME3 ;
 ANTENNAGATEAREA                          0.288 LAYER ME4 ;
 ANTENNADIFFAREA                          0.206 LAYER ME2 ;
 ANTENNADIFFAREA                          0.206 LAYER ME3 ;
 ANTENNADIFFAREA                          0.206 LAYER ME4 ;
 ANTENNAMAXAREACAR                        5.844 LAYER ME2 ;
 ANTENNAMAXAREACAR                        6.511 LAYER ME3 ;
 ANTENNAMAXAREACAR                        7.178 LAYER ME4 ;
END WEB7
PIN DI83
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 375.043 0.000 375.363 0.600 ;
  LAYER ME3 ;
  RECT 375.043 0.000 375.363 0.600 ;
  LAYER ME2 ;
  RECT 375.043 0.000 375.363 0.600 ;
  LAYER ME1 ;
  RECT 375.043 0.000 375.363 0.600 ;
 END
 ANTENNAPARTIALMETALAREA                  1.058 LAYER ME2 ;
 ANTENNAGATEAREA                          0.072 LAYER ME2 ;
 ANTENNAGATEAREA                          0.072 LAYER ME3 ;
 ANTENNAGATEAREA                          0.072 LAYER ME4 ;
 ANTENNADIFFAREA                          0.160 LAYER ME2 ;
 ANTENNADIFFAREA                          0.160 LAYER ME3 ;
 ANTENNADIFFAREA                          0.160 LAYER ME4 ;
 ANTENNAMAXAREACAR                       21.782 LAYER ME2 ;
 ANTENNAMAXAREACAR                       24.449 LAYER ME3 ;
 ANTENNAMAXAREACAR                       27.116 LAYER ME4 ;
END DI83
PIN DO83
  DIRECTION OUTPUT ;
 PORT
  LAYER ME4 ;
  RECT 374.481 0.000 374.801 0.600 ;
  LAYER ME3 ;
  RECT 374.481 0.000 374.801 0.600 ;
  LAYER ME2 ;
  RECT 374.481 0.000 374.801 0.600 ;
  LAYER ME1 ;
  RECT 374.481 0.000 374.801 0.600 ;
 END
 ANTENNAPARTIALMETALAREA                  5.273 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME3 ;
 ANTENNADIFFAREA                          1.293 LAYER ME4 ;
END DO83
PIN DI82
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 371.039 0.000 371.359 0.600 ;
  LAYER ME3 ;
  RECT 371.039 0.000 371.359 0.600 ;
  LAYER ME2 ;
  RECT 371.039 0.000 371.359 0.600 ;
  LAYER ME1 ;
  RECT 371.039 0.000 371.359 0.600 ;
 END
 ANTENNAPARTIALMETALAREA                  1.058 LAYER ME2 ;
 ANTENNAGATEAREA                          0.072 LAYER ME2 ;
 ANTENNAGATEAREA                          0.072 LAYER ME3 ;
 ANTENNAGATEAREA                          0.072 LAYER ME4 ;
 ANTENNADIFFAREA                          0.160 LAYER ME2 ;
 ANTENNADIFFAREA                          0.160 LAYER ME3 ;
 ANTENNADIFFAREA                          0.160 LAYER ME4 ;
 ANTENNAMAXAREACAR                       21.782 LAYER ME2 ;
 ANTENNAMAXAREACAR                       24.449 LAYER ME3 ;
 ANTENNAMAXAREACAR                       27.116 LAYER ME4 ;
END DI82
PIN DO82
  DIRECTION OUTPUT ;
 PORT
  LAYER ME4 ;
  RECT 370.477 0.000 370.797 0.600 ;
  LAYER ME3 ;
  RECT 370.477 0.000 370.797 0.600 ;
  LAYER ME2 ;
  RECT 370.477 0.000 370.797 0.600 ;
  LAYER ME1 ;
  RECT 370.477 0.000 370.797 0.600 ;
 END
 ANTENNAPARTIALMETALAREA                  5.273 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME3 ;
 ANTENNADIFFAREA                          1.293 LAYER ME4 ;
END DO82
PIN DI81
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 367.035 0.000 367.355 0.600 ;
  LAYER ME3 ;
  RECT 367.035 0.000 367.355 0.600 ;
  LAYER ME2 ;
  RECT 367.035 0.000 367.355 0.600 ;
  LAYER ME1 ;
  RECT 367.035 0.000 367.355 0.600 ;
 END
 ANTENNAPARTIALMETALAREA                  1.058 LAYER ME2 ;
 ANTENNAGATEAREA                          0.072 LAYER ME2 ;
 ANTENNAGATEAREA                          0.072 LAYER ME3 ;
 ANTENNAGATEAREA                          0.072 LAYER ME4 ;
 ANTENNADIFFAREA                          0.160 LAYER ME2 ;
 ANTENNADIFFAREA                          0.160 LAYER ME3 ;
 ANTENNADIFFAREA                          0.160 LAYER ME4 ;
 ANTENNAMAXAREACAR                       21.782 LAYER ME2 ;
 ANTENNAMAXAREACAR                       24.449 LAYER ME3 ;
 ANTENNAMAXAREACAR                       27.116 LAYER ME4 ;
END DI81
PIN DO81
  DIRECTION OUTPUT ;
 PORT
  LAYER ME4 ;
  RECT 366.473 0.000 366.793 0.600 ;
  LAYER ME3 ;
  RECT 366.473 0.000 366.793 0.600 ;
  LAYER ME2 ;
  RECT 366.473 0.000 366.793 0.600 ;
  LAYER ME1 ;
  RECT 366.473 0.000 366.793 0.600 ;
 END
 ANTENNAPARTIALMETALAREA                  5.273 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME3 ;
 ANTENNADIFFAREA                          1.293 LAYER ME4 ;
END DO81
PIN DI80
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 363.031 0.000 363.351 0.600 ;
  LAYER ME3 ;
  RECT 363.031 0.000 363.351 0.600 ;
  LAYER ME2 ;
  RECT 363.031 0.000 363.351 0.600 ;
  LAYER ME1 ;
  RECT 363.031 0.000 363.351 0.600 ;
 END
 ANTENNAPARTIALMETALAREA                  1.058 LAYER ME2 ;
 ANTENNAGATEAREA                          0.072 LAYER ME2 ;
 ANTENNAGATEAREA                          0.072 LAYER ME3 ;
 ANTENNAGATEAREA                          0.072 LAYER ME4 ;
 ANTENNADIFFAREA                          0.160 LAYER ME2 ;
 ANTENNADIFFAREA                          0.160 LAYER ME3 ;
 ANTENNADIFFAREA                          0.160 LAYER ME4 ;
 ANTENNAMAXAREACAR                       21.782 LAYER ME2 ;
 ANTENNAMAXAREACAR                       24.449 LAYER ME3 ;
 ANTENNAMAXAREACAR                       27.116 LAYER ME4 ;
END DI80
PIN DO80
  DIRECTION OUTPUT ;
 PORT
  LAYER ME4 ;
  RECT 362.469 0.000 362.789 0.600 ;
  LAYER ME3 ;
  RECT 362.469 0.000 362.789 0.600 ;
  LAYER ME2 ;
  RECT 362.469 0.000 362.789 0.600 ;
  LAYER ME1 ;
  RECT 362.469 0.000 362.789 0.600 ;
 END
 ANTENNAPARTIALMETALAREA                  5.273 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME3 ;
 ANTENNADIFFAREA                          1.293 LAYER ME4 ;
END DO80
PIN DI79
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 359.027 0.000 359.347 0.600 ;
  LAYER ME3 ;
  RECT 359.027 0.000 359.347 0.600 ;
  LAYER ME2 ;
  RECT 359.027 0.000 359.347 0.600 ;
  LAYER ME1 ;
  RECT 359.027 0.000 359.347 0.600 ;
 END
 ANTENNAPARTIALMETALAREA                  1.058 LAYER ME2 ;
 ANTENNAGATEAREA                          0.072 LAYER ME2 ;
 ANTENNAGATEAREA                          0.072 LAYER ME3 ;
 ANTENNAGATEAREA                          0.072 LAYER ME4 ;
 ANTENNADIFFAREA                          0.160 LAYER ME2 ;
 ANTENNADIFFAREA                          0.160 LAYER ME3 ;
 ANTENNADIFFAREA                          0.160 LAYER ME4 ;
 ANTENNAMAXAREACAR                       21.782 LAYER ME2 ;
 ANTENNAMAXAREACAR                       24.449 LAYER ME3 ;
 ANTENNAMAXAREACAR                       27.116 LAYER ME4 ;
END DI79
PIN DO79
  DIRECTION OUTPUT ;
 PORT
  LAYER ME4 ;
  RECT 358.465 0.000 358.785 0.600 ;
  LAYER ME3 ;
  RECT 358.465 0.000 358.785 0.600 ;
  LAYER ME2 ;
  RECT 358.465 0.000 358.785 0.600 ;
  LAYER ME1 ;
  RECT 358.465 0.000 358.785 0.600 ;
 END
 ANTENNAPARTIALMETALAREA                  5.273 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME3 ;
 ANTENNADIFFAREA                          1.293 LAYER ME4 ;
END DO79
PIN DI78
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 355.023 0.000 355.343 0.600 ;
  LAYER ME3 ;
  RECT 355.023 0.000 355.343 0.600 ;
  LAYER ME2 ;
  RECT 355.023 0.000 355.343 0.600 ;
  LAYER ME1 ;
  RECT 355.023 0.000 355.343 0.600 ;
 END
 ANTENNAPARTIALMETALAREA                  1.058 LAYER ME2 ;
 ANTENNAGATEAREA                          0.072 LAYER ME2 ;
 ANTENNAGATEAREA                          0.072 LAYER ME3 ;
 ANTENNAGATEAREA                          0.072 LAYER ME4 ;
 ANTENNADIFFAREA                          0.160 LAYER ME2 ;
 ANTENNADIFFAREA                          0.160 LAYER ME3 ;
 ANTENNADIFFAREA                          0.160 LAYER ME4 ;
 ANTENNAMAXAREACAR                       21.782 LAYER ME2 ;
 ANTENNAMAXAREACAR                       24.449 LAYER ME3 ;
 ANTENNAMAXAREACAR                       27.116 LAYER ME4 ;
END DI78
PIN DO78
  DIRECTION OUTPUT ;
 PORT
  LAYER ME4 ;
  RECT 354.461 0.000 354.781 0.600 ;
  LAYER ME3 ;
  RECT 354.461 0.000 354.781 0.600 ;
  LAYER ME2 ;
  RECT 354.461 0.000 354.781 0.600 ;
  LAYER ME1 ;
  RECT 354.461 0.000 354.781 0.600 ;
 END
 ANTENNAPARTIALMETALAREA                  5.273 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME3 ;
 ANTENNADIFFAREA                          1.293 LAYER ME4 ;
END DO78
PIN DI77
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 351.019 0.000 351.339 0.600 ;
  LAYER ME3 ;
  RECT 351.019 0.000 351.339 0.600 ;
  LAYER ME2 ;
  RECT 351.019 0.000 351.339 0.600 ;
  LAYER ME1 ;
  RECT 351.019 0.000 351.339 0.600 ;
 END
 ANTENNAPARTIALMETALAREA                  1.058 LAYER ME2 ;
 ANTENNAGATEAREA                          0.072 LAYER ME2 ;
 ANTENNAGATEAREA                          0.072 LAYER ME3 ;
 ANTENNAGATEAREA                          0.072 LAYER ME4 ;
 ANTENNADIFFAREA                          0.160 LAYER ME2 ;
 ANTENNADIFFAREA                          0.160 LAYER ME3 ;
 ANTENNADIFFAREA                          0.160 LAYER ME4 ;
 ANTENNAMAXAREACAR                       21.782 LAYER ME2 ;
 ANTENNAMAXAREACAR                       24.449 LAYER ME3 ;
 ANTENNAMAXAREACAR                       27.116 LAYER ME4 ;
END DI77
PIN DO77
  DIRECTION OUTPUT ;
 PORT
  LAYER ME4 ;
  RECT 350.457 0.000 350.777 0.600 ;
  LAYER ME3 ;
  RECT 350.457 0.000 350.777 0.600 ;
  LAYER ME2 ;
  RECT 350.457 0.000 350.777 0.600 ;
  LAYER ME1 ;
  RECT 350.457 0.000 350.777 0.600 ;
 END
 ANTENNAPARTIALMETALAREA                  5.273 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME3 ;
 ANTENNADIFFAREA                          1.293 LAYER ME4 ;
END DO77
PIN DI76
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 347.015 0.000 347.335 0.600 ;
  LAYER ME3 ;
  RECT 347.015 0.000 347.335 0.600 ;
  LAYER ME2 ;
  RECT 347.015 0.000 347.335 0.600 ;
  LAYER ME1 ;
  RECT 347.015 0.000 347.335 0.600 ;
 END
 ANTENNAPARTIALMETALAREA                  1.058 LAYER ME2 ;
 ANTENNAGATEAREA                          0.072 LAYER ME2 ;
 ANTENNAGATEAREA                          0.072 LAYER ME3 ;
 ANTENNAGATEAREA                          0.072 LAYER ME4 ;
 ANTENNADIFFAREA                          0.160 LAYER ME2 ;
 ANTENNADIFFAREA                          0.160 LAYER ME3 ;
 ANTENNADIFFAREA                          0.160 LAYER ME4 ;
 ANTENNAMAXAREACAR                       21.782 LAYER ME2 ;
 ANTENNAMAXAREACAR                       24.449 LAYER ME3 ;
 ANTENNAMAXAREACAR                       27.116 LAYER ME4 ;
END DI76
PIN DO76
  DIRECTION OUTPUT ;
 PORT
  LAYER ME4 ;
  RECT 346.453 0.000 346.773 0.600 ;
  LAYER ME3 ;
  RECT 346.453 0.000 346.773 0.600 ;
  LAYER ME2 ;
  RECT 346.453 0.000 346.773 0.600 ;
  LAYER ME1 ;
  RECT 346.453 0.000 346.773 0.600 ;
 END
 ANTENNAPARTIALMETALAREA                  5.273 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME3 ;
 ANTENNADIFFAREA                          1.293 LAYER ME4 ;
END DO76
PIN DI75
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 343.011 0.000 343.331 0.600 ;
  LAYER ME3 ;
  RECT 343.011 0.000 343.331 0.600 ;
  LAYER ME2 ;
  RECT 343.011 0.000 343.331 0.600 ;
  LAYER ME1 ;
  RECT 343.011 0.000 343.331 0.600 ;
 END
 ANTENNAPARTIALMETALAREA                  1.058 LAYER ME2 ;
 ANTENNAGATEAREA                          0.072 LAYER ME2 ;
 ANTENNAGATEAREA                          0.072 LAYER ME3 ;
 ANTENNAGATEAREA                          0.072 LAYER ME4 ;
 ANTENNADIFFAREA                          0.160 LAYER ME2 ;
 ANTENNADIFFAREA                          0.160 LAYER ME3 ;
 ANTENNADIFFAREA                          0.160 LAYER ME4 ;
 ANTENNAMAXAREACAR                       21.782 LAYER ME2 ;
 ANTENNAMAXAREACAR                       24.449 LAYER ME3 ;
 ANTENNAMAXAREACAR                       27.116 LAYER ME4 ;
END DI75
PIN DO75
  DIRECTION OUTPUT ;
 PORT
  LAYER ME4 ;
  RECT 342.449 0.000 342.769 0.600 ;
  LAYER ME3 ;
  RECT 342.449 0.000 342.769 0.600 ;
  LAYER ME2 ;
  RECT 342.449 0.000 342.769 0.600 ;
  LAYER ME1 ;
  RECT 342.449 0.000 342.769 0.600 ;
 END
 ANTENNAPARTIALMETALAREA                  5.273 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME3 ;
 ANTENNADIFFAREA                          1.293 LAYER ME4 ;
END DO75
PIN DI74
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 339.007 0.000 339.327 0.600 ;
  LAYER ME3 ;
  RECT 339.007 0.000 339.327 0.600 ;
  LAYER ME2 ;
  RECT 339.007 0.000 339.327 0.600 ;
  LAYER ME1 ;
  RECT 339.007 0.000 339.327 0.600 ;
 END
 ANTENNAPARTIALMETALAREA                  1.058 LAYER ME2 ;
 ANTENNAGATEAREA                          0.072 LAYER ME2 ;
 ANTENNAGATEAREA                          0.072 LAYER ME3 ;
 ANTENNAGATEAREA                          0.072 LAYER ME4 ;
 ANTENNADIFFAREA                          0.160 LAYER ME2 ;
 ANTENNADIFFAREA                          0.160 LAYER ME3 ;
 ANTENNADIFFAREA                          0.160 LAYER ME4 ;
 ANTENNAMAXAREACAR                       21.782 LAYER ME2 ;
 ANTENNAMAXAREACAR                       24.449 LAYER ME3 ;
 ANTENNAMAXAREACAR                       27.116 LAYER ME4 ;
END DI74
PIN DO74
  DIRECTION OUTPUT ;
 PORT
  LAYER ME4 ;
  RECT 338.445 0.000 338.765 0.600 ;
  LAYER ME3 ;
  RECT 338.445 0.000 338.765 0.600 ;
  LAYER ME2 ;
  RECT 338.445 0.000 338.765 0.600 ;
  LAYER ME1 ;
  RECT 338.445 0.000 338.765 0.600 ;
 END
 ANTENNAPARTIALMETALAREA                  5.273 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME3 ;
 ANTENNADIFFAREA                          1.293 LAYER ME4 ;
END DO74
PIN DI73
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 335.003 0.000 335.323 0.600 ;
  LAYER ME3 ;
  RECT 335.003 0.000 335.323 0.600 ;
  LAYER ME2 ;
  RECT 335.003 0.000 335.323 0.600 ;
  LAYER ME1 ;
  RECT 335.003 0.000 335.323 0.600 ;
 END
 ANTENNAPARTIALMETALAREA                  1.058 LAYER ME2 ;
 ANTENNAGATEAREA                          0.072 LAYER ME2 ;
 ANTENNAGATEAREA                          0.072 LAYER ME3 ;
 ANTENNAGATEAREA                          0.072 LAYER ME4 ;
 ANTENNADIFFAREA                          0.160 LAYER ME2 ;
 ANTENNADIFFAREA                          0.160 LAYER ME3 ;
 ANTENNADIFFAREA                          0.160 LAYER ME4 ;
 ANTENNAMAXAREACAR                       21.782 LAYER ME2 ;
 ANTENNAMAXAREACAR                       24.449 LAYER ME3 ;
 ANTENNAMAXAREACAR                       27.116 LAYER ME4 ;
END DI73
PIN DO73
  DIRECTION OUTPUT ;
 PORT
  LAYER ME4 ;
  RECT 334.441 0.000 334.761 0.600 ;
  LAYER ME3 ;
  RECT 334.441 0.000 334.761 0.600 ;
  LAYER ME2 ;
  RECT 334.441 0.000 334.761 0.600 ;
  LAYER ME1 ;
  RECT 334.441 0.000 334.761 0.600 ;
 END
 ANTENNAPARTIALMETALAREA                  5.273 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME3 ;
 ANTENNADIFFAREA                          1.293 LAYER ME4 ;
END DO73
PIN DI72
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 330.437 0.000 330.757 0.600 ;
  LAYER ME3 ;
  RECT 330.437 0.000 330.757 0.600 ;
  LAYER ME2 ;
  RECT 330.437 0.000 330.757 0.600 ;
  LAYER ME1 ;
  RECT 330.437 0.000 330.757 0.600 ;
 END
 ANTENNAPARTIALMETALAREA                  0.346 LAYER ME1 ;
 ANTENNAPARTIALMETALAREA                  1.466 LAYER ME2 ;
 ANTENNAPARTIALMETALAREA                  0.508 LAYER ME3 ;
 ANTENNAGATEAREA                          0.072 LAYER ME3 ;
 ANTENNAGATEAREA                          0.072 LAYER ME4 ;
 ANTENNADIFFAREA                          0.218 LAYER ME1 ;
 ANTENNADIFFAREA                          0.218 LAYER ME2 ;
 ANTENNADIFFAREA                          0.218 LAYER ME3 ;
 ANTENNADIFFAREA                          0.218 LAYER ME4 ;
 ANTENNAMAXAREACAR                       17.267 LAYER ME3 ;
 ANTENNAMAXAREACAR                       19.933 LAYER ME4 ;
END DI72
PIN DO72
  DIRECTION OUTPUT ;
 PORT
  LAYER ME4 ;
  RECT 330.999 0.000 331.319 0.600 ;
  LAYER ME3 ;
  RECT 330.999 0.000 331.319 0.600 ;
  LAYER ME2 ;
  RECT 330.999 0.000 331.319 0.600 ;
  LAYER ME1 ;
  RECT 330.999 0.000 331.319 0.600 ;
 END
 ANTENNAPARTIALMETALAREA                  5.602 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME3 ;
 ANTENNADIFFAREA                          1.293 LAYER ME4 ;
END DO72
PIN WEB6
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 328.997 0.000 329.317 0.600 ;
  LAYER ME3 ;
  RECT 328.997 0.000 329.317 0.600 ;
  LAYER ME2 ;
  RECT 328.997 0.000 329.317 0.600 ;
  LAYER ME1 ;
  RECT 328.997 0.000 329.317 0.600 ;
 END
 ANTENNAPARTIALMETALAREA                  1.036 LAYER ME2 ;
 ANTENNAGATEAREA                          0.288 LAYER ME2 ;
 ANTENNAGATEAREA                          0.288 LAYER ME3 ;
 ANTENNAGATEAREA                          0.288 LAYER ME4 ;
 ANTENNADIFFAREA                          0.206 LAYER ME2 ;
 ANTENNADIFFAREA                          0.206 LAYER ME3 ;
 ANTENNADIFFAREA                          0.206 LAYER ME4 ;
 ANTENNAMAXAREACAR                        5.844 LAYER ME2 ;
 ANTENNAMAXAREACAR                        6.511 LAYER ME3 ;
 ANTENNAMAXAREACAR                        7.178 LAYER ME4 ;
END WEB6
PIN DI71
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 326.995 0.000 327.315 0.600 ;
  LAYER ME3 ;
  RECT 326.995 0.000 327.315 0.600 ;
  LAYER ME2 ;
  RECT 326.995 0.000 327.315 0.600 ;
  LAYER ME1 ;
  RECT 326.995 0.000 327.315 0.600 ;
 END
 ANTENNAPARTIALMETALAREA                  1.058 LAYER ME2 ;
 ANTENNAGATEAREA                          0.072 LAYER ME2 ;
 ANTENNAGATEAREA                          0.072 LAYER ME3 ;
 ANTENNAGATEAREA                          0.072 LAYER ME4 ;
 ANTENNADIFFAREA                          0.160 LAYER ME2 ;
 ANTENNADIFFAREA                          0.160 LAYER ME3 ;
 ANTENNADIFFAREA                          0.160 LAYER ME4 ;
 ANTENNAMAXAREACAR                       21.782 LAYER ME2 ;
 ANTENNAMAXAREACAR                       24.449 LAYER ME3 ;
 ANTENNAMAXAREACAR                       27.116 LAYER ME4 ;
END DI71
PIN DO71
  DIRECTION OUTPUT ;
 PORT
  LAYER ME4 ;
  RECT 326.433 0.000 326.753 0.600 ;
  LAYER ME3 ;
  RECT 326.433 0.000 326.753 0.600 ;
  LAYER ME2 ;
  RECT 326.433 0.000 326.753 0.600 ;
  LAYER ME1 ;
  RECT 326.433 0.000 326.753 0.600 ;
 END
 ANTENNAPARTIALMETALAREA                  5.273 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME3 ;
 ANTENNADIFFAREA                          1.293 LAYER ME4 ;
END DO71
PIN DI70
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 322.991 0.000 323.311 0.600 ;
  LAYER ME3 ;
  RECT 322.991 0.000 323.311 0.600 ;
  LAYER ME2 ;
  RECT 322.991 0.000 323.311 0.600 ;
  LAYER ME1 ;
  RECT 322.991 0.000 323.311 0.600 ;
 END
 ANTENNAPARTIALMETALAREA                  1.058 LAYER ME2 ;
 ANTENNAGATEAREA                          0.072 LAYER ME2 ;
 ANTENNAGATEAREA                          0.072 LAYER ME3 ;
 ANTENNAGATEAREA                          0.072 LAYER ME4 ;
 ANTENNADIFFAREA                          0.160 LAYER ME2 ;
 ANTENNADIFFAREA                          0.160 LAYER ME3 ;
 ANTENNADIFFAREA                          0.160 LAYER ME4 ;
 ANTENNAMAXAREACAR                       21.782 LAYER ME2 ;
 ANTENNAMAXAREACAR                       24.449 LAYER ME3 ;
 ANTENNAMAXAREACAR                       27.116 LAYER ME4 ;
END DI70
PIN DO70
  DIRECTION OUTPUT ;
 PORT
  LAYER ME4 ;
  RECT 322.429 0.000 322.749 0.600 ;
  LAYER ME3 ;
  RECT 322.429 0.000 322.749 0.600 ;
  LAYER ME2 ;
  RECT 322.429 0.000 322.749 0.600 ;
  LAYER ME1 ;
  RECT 322.429 0.000 322.749 0.600 ;
 END
 ANTENNAPARTIALMETALAREA                  5.273 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME3 ;
 ANTENNADIFFAREA                          1.293 LAYER ME4 ;
END DO70
PIN DI69
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 318.987 0.000 319.307 0.600 ;
  LAYER ME3 ;
  RECT 318.987 0.000 319.307 0.600 ;
  LAYER ME2 ;
  RECT 318.987 0.000 319.307 0.600 ;
  LAYER ME1 ;
  RECT 318.987 0.000 319.307 0.600 ;
 END
 ANTENNAPARTIALMETALAREA                  1.058 LAYER ME2 ;
 ANTENNAGATEAREA                          0.072 LAYER ME2 ;
 ANTENNAGATEAREA                          0.072 LAYER ME3 ;
 ANTENNAGATEAREA                          0.072 LAYER ME4 ;
 ANTENNADIFFAREA                          0.160 LAYER ME2 ;
 ANTENNADIFFAREA                          0.160 LAYER ME3 ;
 ANTENNADIFFAREA                          0.160 LAYER ME4 ;
 ANTENNAMAXAREACAR                       21.782 LAYER ME2 ;
 ANTENNAMAXAREACAR                       24.449 LAYER ME3 ;
 ANTENNAMAXAREACAR                       27.116 LAYER ME4 ;
END DI69
PIN DO69
  DIRECTION OUTPUT ;
 PORT
  LAYER ME4 ;
  RECT 318.425 0.000 318.745 0.600 ;
  LAYER ME3 ;
  RECT 318.425 0.000 318.745 0.600 ;
  LAYER ME2 ;
  RECT 318.425 0.000 318.745 0.600 ;
  LAYER ME1 ;
  RECT 318.425 0.000 318.745 0.600 ;
 END
 ANTENNAPARTIALMETALAREA                  5.273 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME3 ;
 ANTENNADIFFAREA                          1.293 LAYER ME4 ;
END DO69
PIN DI68
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 314.983 0.000 315.303 0.600 ;
  LAYER ME3 ;
  RECT 314.983 0.000 315.303 0.600 ;
  LAYER ME2 ;
  RECT 314.983 0.000 315.303 0.600 ;
  LAYER ME1 ;
  RECT 314.983 0.000 315.303 0.600 ;
 END
 ANTENNAPARTIALMETALAREA                  1.058 LAYER ME2 ;
 ANTENNAGATEAREA                          0.072 LAYER ME2 ;
 ANTENNAGATEAREA                          0.072 LAYER ME3 ;
 ANTENNAGATEAREA                          0.072 LAYER ME4 ;
 ANTENNADIFFAREA                          0.160 LAYER ME2 ;
 ANTENNADIFFAREA                          0.160 LAYER ME3 ;
 ANTENNADIFFAREA                          0.160 LAYER ME4 ;
 ANTENNAMAXAREACAR                       21.782 LAYER ME2 ;
 ANTENNAMAXAREACAR                       24.449 LAYER ME3 ;
 ANTENNAMAXAREACAR                       27.116 LAYER ME4 ;
END DI68
PIN DO68
  DIRECTION OUTPUT ;
 PORT
  LAYER ME4 ;
  RECT 314.421 0.000 314.741 0.600 ;
  LAYER ME3 ;
  RECT 314.421 0.000 314.741 0.600 ;
  LAYER ME2 ;
  RECT 314.421 0.000 314.741 0.600 ;
  LAYER ME1 ;
  RECT 314.421 0.000 314.741 0.600 ;
 END
 ANTENNAPARTIALMETALAREA                  5.273 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME3 ;
 ANTENNADIFFAREA                          1.293 LAYER ME4 ;
END DO68
PIN DI67
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 310.979 0.000 311.299 0.600 ;
  LAYER ME3 ;
  RECT 310.979 0.000 311.299 0.600 ;
  LAYER ME2 ;
  RECT 310.979 0.000 311.299 0.600 ;
  LAYER ME1 ;
  RECT 310.979 0.000 311.299 0.600 ;
 END
 ANTENNAPARTIALMETALAREA                  1.058 LAYER ME2 ;
 ANTENNAGATEAREA                          0.072 LAYER ME2 ;
 ANTENNAGATEAREA                          0.072 LAYER ME3 ;
 ANTENNAGATEAREA                          0.072 LAYER ME4 ;
 ANTENNADIFFAREA                          0.160 LAYER ME2 ;
 ANTENNADIFFAREA                          0.160 LAYER ME3 ;
 ANTENNADIFFAREA                          0.160 LAYER ME4 ;
 ANTENNAMAXAREACAR                       21.782 LAYER ME2 ;
 ANTENNAMAXAREACAR                       24.449 LAYER ME3 ;
 ANTENNAMAXAREACAR                       27.116 LAYER ME4 ;
END DI67
PIN DO67
  DIRECTION OUTPUT ;
 PORT
  LAYER ME4 ;
  RECT 310.417 0.000 310.737 0.600 ;
  LAYER ME3 ;
  RECT 310.417 0.000 310.737 0.600 ;
  LAYER ME2 ;
  RECT 310.417 0.000 310.737 0.600 ;
  LAYER ME1 ;
  RECT 310.417 0.000 310.737 0.600 ;
 END
 ANTENNAPARTIALMETALAREA                  5.273 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME3 ;
 ANTENNADIFFAREA                          1.293 LAYER ME4 ;
END DO67
PIN DI66
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 306.975 0.000 307.295 0.600 ;
  LAYER ME3 ;
  RECT 306.975 0.000 307.295 0.600 ;
  LAYER ME2 ;
  RECT 306.975 0.000 307.295 0.600 ;
  LAYER ME1 ;
  RECT 306.975 0.000 307.295 0.600 ;
 END
 ANTENNAPARTIALMETALAREA                  1.058 LAYER ME2 ;
 ANTENNAGATEAREA                          0.072 LAYER ME2 ;
 ANTENNAGATEAREA                          0.072 LAYER ME3 ;
 ANTENNAGATEAREA                          0.072 LAYER ME4 ;
 ANTENNADIFFAREA                          0.160 LAYER ME2 ;
 ANTENNADIFFAREA                          0.160 LAYER ME3 ;
 ANTENNADIFFAREA                          0.160 LAYER ME4 ;
 ANTENNAMAXAREACAR                       21.782 LAYER ME2 ;
 ANTENNAMAXAREACAR                       24.449 LAYER ME3 ;
 ANTENNAMAXAREACAR                       27.116 LAYER ME4 ;
END DI66
PIN DO66
  DIRECTION OUTPUT ;
 PORT
  LAYER ME4 ;
  RECT 306.413 0.000 306.733 0.600 ;
  LAYER ME3 ;
  RECT 306.413 0.000 306.733 0.600 ;
  LAYER ME2 ;
  RECT 306.413 0.000 306.733 0.600 ;
  LAYER ME1 ;
  RECT 306.413 0.000 306.733 0.600 ;
 END
 ANTENNAPARTIALMETALAREA                  5.273 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME3 ;
 ANTENNADIFFAREA                          1.293 LAYER ME4 ;
END DO66
PIN DI65
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 302.971 0.000 303.291 0.600 ;
  LAYER ME3 ;
  RECT 302.971 0.000 303.291 0.600 ;
  LAYER ME2 ;
  RECT 302.971 0.000 303.291 0.600 ;
  LAYER ME1 ;
  RECT 302.971 0.000 303.291 0.600 ;
 END
 ANTENNAPARTIALMETALAREA                  1.058 LAYER ME2 ;
 ANTENNAGATEAREA                          0.072 LAYER ME2 ;
 ANTENNAGATEAREA                          0.072 LAYER ME3 ;
 ANTENNAGATEAREA                          0.072 LAYER ME4 ;
 ANTENNADIFFAREA                          0.160 LAYER ME2 ;
 ANTENNADIFFAREA                          0.160 LAYER ME3 ;
 ANTENNADIFFAREA                          0.160 LAYER ME4 ;
 ANTENNAMAXAREACAR                       21.782 LAYER ME2 ;
 ANTENNAMAXAREACAR                       24.449 LAYER ME3 ;
 ANTENNAMAXAREACAR                       27.116 LAYER ME4 ;
END DI65
PIN DO65
  DIRECTION OUTPUT ;
 PORT
  LAYER ME4 ;
  RECT 302.409 0.000 302.729 0.600 ;
  LAYER ME3 ;
  RECT 302.409 0.000 302.729 0.600 ;
  LAYER ME2 ;
  RECT 302.409 0.000 302.729 0.600 ;
  LAYER ME1 ;
  RECT 302.409 0.000 302.729 0.600 ;
 END
 ANTENNAPARTIALMETALAREA                  5.273 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME3 ;
 ANTENNADIFFAREA                          1.293 LAYER ME4 ;
END DO65
PIN DI64
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 298.967 0.000 299.287 0.600 ;
  LAYER ME3 ;
  RECT 298.967 0.000 299.287 0.600 ;
  LAYER ME2 ;
  RECT 298.967 0.000 299.287 0.600 ;
  LAYER ME1 ;
  RECT 298.967 0.000 299.287 0.600 ;
 END
 ANTENNAPARTIALMETALAREA                  1.058 LAYER ME2 ;
 ANTENNAGATEAREA                          0.072 LAYER ME2 ;
 ANTENNAGATEAREA                          0.072 LAYER ME3 ;
 ANTENNAGATEAREA                          0.072 LAYER ME4 ;
 ANTENNADIFFAREA                          0.160 LAYER ME2 ;
 ANTENNADIFFAREA                          0.160 LAYER ME3 ;
 ANTENNADIFFAREA                          0.160 LAYER ME4 ;
 ANTENNAMAXAREACAR                       21.782 LAYER ME2 ;
 ANTENNAMAXAREACAR                       24.449 LAYER ME3 ;
 ANTENNAMAXAREACAR                       27.116 LAYER ME4 ;
END DI64
PIN DO64
  DIRECTION OUTPUT ;
 PORT
  LAYER ME4 ;
  RECT 298.405 0.000 298.725 0.600 ;
  LAYER ME3 ;
  RECT 298.405 0.000 298.725 0.600 ;
  LAYER ME2 ;
  RECT 298.405 0.000 298.725 0.600 ;
  LAYER ME1 ;
  RECT 298.405 0.000 298.725 0.600 ;
 END
 ANTENNAPARTIALMETALAREA                  5.273 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME3 ;
 ANTENNADIFFAREA                          1.293 LAYER ME4 ;
END DO64
PIN DI63
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 294.963 0.000 295.283 0.600 ;
  LAYER ME3 ;
  RECT 294.963 0.000 295.283 0.600 ;
  LAYER ME2 ;
  RECT 294.963 0.000 295.283 0.600 ;
  LAYER ME1 ;
  RECT 294.963 0.000 295.283 0.600 ;
 END
 ANTENNAPARTIALMETALAREA                  1.058 LAYER ME2 ;
 ANTENNAGATEAREA                          0.072 LAYER ME2 ;
 ANTENNAGATEAREA                          0.072 LAYER ME3 ;
 ANTENNAGATEAREA                          0.072 LAYER ME4 ;
 ANTENNADIFFAREA                          0.160 LAYER ME2 ;
 ANTENNADIFFAREA                          0.160 LAYER ME3 ;
 ANTENNADIFFAREA                          0.160 LAYER ME4 ;
 ANTENNAMAXAREACAR                       21.782 LAYER ME2 ;
 ANTENNAMAXAREACAR                       24.449 LAYER ME3 ;
 ANTENNAMAXAREACAR                       27.116 LAYER ME4 ;
END DI63
PIN DO63
  DIRECTION OUTPUT ;
 PORT
  LAYER ME4 ;
  RECT 294.401 0.000 294.721 0.600 ;
  LAYER ME3 ;
  RECT 294.401 0.000 294.721 0.600 ;
  LAYER ME2 ;
  RECT 294.401 0.000 294.721 0.600 ;
  LAYER ME1 ;
  RECT 294.401 0.000 294.721 0.600 ;
 END
 ANTENNAPARTIALMETALAREA                  5.273 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME3 ;
 ANTENNADIFFAREA                          1.293 LAYER ME4 ;
END DO63
PIN DI62
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 290.959 0.000 291.279 0.600 ;
  LAYER ME3 ;
  RECT 290.959 0.000 291.279 0.600 ;
  LAYER ME2 ;
  RECT 290.959 0.000 291.279 0.600 ;
  LAYER ME1 ;
  RECT 290.959 0.000 291.279 0.600 ;
 END
 ANTENNAPARTIALMETALAREA                  1.058 LAYER ME2 ;
 ANTENNAGATEAREA                          0.072 LAYER ME2 ;
 ANTENNAGATEAREA                          0.072 LAYER ME3 ;
 ANTENNAGATEAREA                          0.072 LAYER ME4 ;
 ANTENNADIFFAREA                          0.160 LAYER ME2 ;
 ANTENNADIFFAREA                          0.160 LAYER ME3 ;
 ANTENNADIFFAREA                          0.160 LAYER ME4 ;
 ANTENNAMAXAREACAR                       21.782 LAYER ME2 ;
 ANTENNAMAXAREACAR                       24.449 LAYER ME3 ;
 ANTENNAMAXAREACAR                       27.116 LAYER ME4 ;
END DI62
PIN DO62
  DIRECTION OUTPUT ;
 PORT
  LAYER ME4 ;
  RECT 290.397 0.000 290.717 0.600 ;
  LAYER ME3 ;
  RECT 290.397 0.000 290.717 0.600 ;
  LAYER ME2 ;
  RECT 290.397 0.000 290.717 0.600 ;
  LAYER ME1 ;
  RECT 290.397 0.000 290.717 0.600 ;
 END
 ANTENNAPARTIALMETALAREA                  5.273 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME3 ;
 ANTENNADIFFAREA                          1.293 LAYER ME4 ;
END DO62
PIN DI61
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 286.955 0.000 287.275 0.600 ;
  LAYER ME3 ;
  RECT 286.955 0.000 287.275 0.600 ;
  LAYER ME2 ;
  RECT 286.955 0.000 287.275 0.600 ;
  LAYER ME1 ;
  RECT 286.955 0.000 287.275 0.600 ;
 END
 ANTENNAPARTIALMETALAREA                  1.058 LAYER ME2 ;
 ANTENNAGATEAREA                          0.072 LAYER ME2 ;
 ANTENNAGATEAREA                          0.072 LAYER ME3 ;
 ANTENNAGATEAREA                          0.072 LAYER ME4 ;
 ANTENNADIFFAREA                          0.160 LAYER ME2 ;
 ANTENNADIFFAREA                          0.160 LAYER ME3 ;
 ANTENNADIFFAREA                          0.160 LAYER ME4 ;
 ANTENNAMAXAREACAR                       21.782 LAYER ME2 ;
 ANTENNAMAXAREACAR                       24.449 LAYER ME3 ;
 ANTENNAMAXAREACAR                       27.116 LAYER ME4 ;
END DI61
PIN DO61
  DIRECTION OUTPUT ;
 PORT
  LAYER ME4 ;
  RECT 286.393 0.000 286.713 0.600 ;
  LAYER ME3 ;
  RECT 286.393 0.000 286.713 0.600 ;
  LAYER ME2 ;
  RECT 286.393 0.000 286.713 0.600 ;
  LAYER ME1 ;
  RECT 286.393 0.000 286.713 0.600 ;
 END
 ANTENNAPARTIALMETALAREA                  5.273 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME3 ;
 ANTENNADIFFAREA                          1.293 LAYER ME4 ;
END DO61
PIN DI60
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 282.389 0.000 282.709 0.600 ;
  LAYER ME3 ;
  RECT 282.389 0.000 282.709 0.600 ;
  LAYER ME2 ;
  RECT 282.389 0.000 282.709 0.600 ;
  LAYER ME1 ;
  RECT 282.389 0.000 282.709 0.600 ;
 END
 ANTENNAPARTIALMETALAREA                  0.346 LAYER ME1 ;
 ANTENNAPARTIALMETALAREA                  1.466 LAYER ME2 ;
 ANTENNAPARTIALMETALAREA                  0.508 LAYER ME3 ;
 ANTENNAGATEAREA                          0.072 LAYER ME3 ;
 ANTENNAGATEAREA                          0.072 LAYER ME4 ;
 ANTENNADIFFAREA                          0.218 LAYER ME1 ;
 ANTENNADIFFAREA                          0.218 LAYER ME2 ;
 ANTENNADIFFAREA                          0.218 LAYER ME3 ;
 ANTENNADIFFAREA                          0.218 LAYER ME4 ;
 ANTENNAMAXAREACAR                       17.267 LAYER ME3 ;
 ANTENNAMAXAREACAR                       19.933 LAYER ME4 ;
END DI60
PIN DO60
  DIRECTION OUTPUT ;
 PORT
  LAYER ME4 ;
  RECT 282.951 0.000 283.271 0.600 ;
  LAYER ME3 ;
  RECT 282.951 0.000 283.271 0.600 ;
  LAYER ME2 ;
  RECT 282.951 0.000 283.271 0.600 ;
  LAYER ME1 ;
  RECT 282.951 0.000 283.271 0.600 ;
 END
 ANTENNAPARTIALMETALAREA                  5.602 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME3 ;
 ANTENNADIFFAREA                          1.293 LAYER ME4 ;
END DO60
PIN WEB5
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 280.949 0.000 281.269 0.600 ;
  LAYER ME3 ;
  RECT 280.949 0.000 281.269 0.600 ;
  LAYER ME2 ;
  RECT 280.949 0.000 281.269 0.600 ;
  LAYER ME1 ;
  RECT 280.949 0.000 281.269 0.600 ;
 END
 ANTENNAPARTIALMETALAREA                  1.036 LAYER ME2 ;
 ANTENNAGATEAREA                          0.288 LAYER ME2 ;
 ANTENNAGATEAREA                          0.288 LAYER ME3 ;
 ANTENNAGATEAREA                          0.288 LAYER ME4 ;
 ANTENNADIFFAREA                          0.206 LAYER ME2 ;
 ANTENNADIFFAREA                          0.206 LAYER ME3 ;
 ANTENNADIFFAREA                          0.206 LAYER ME4 ;
 ANTENNAMAXAREACAR                        5.844 LAYER ME2 ;
 ANTENNAMAXAREACAR                        6.511 LAYER ME3 ;
 ANTENNAMAXAREACAR                        7.178 LAYER ME4 ;
END WEB5
PIN DI59
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 278.947 0.000 279.267 0.600 ;
  LAYER ME3 ;
  RECT 278.947 0.000 279.267 0.600 ;
  LAYER ME2 ;
  RECT 278.947 0.000 279.267 0.600 ;
  LAYER ME1 ;
  RECT 278.947 0.000 279.267 0.600 ;
 END
 ANTENNAPARTIALMETALAREA                  1.058 LAYER ME2 ;
 ANTENNAGATEAREA                          0.072 LAYER ME2 ;
 ANTENNAGATEAREA                          0.072 LAYER ME3 ;
 ANTENNAGATEAREA                          0.072 LAYER ME4 ;
 ANTENNADIFFAREA                          0.160 LAYER ME2 ;
 ANTENNADIFFAREA                          0.160 LAYER ME3 ;
 ANTENNADIFFAREA                          0.160 LAYER ME4 ;
 ANTENNAMAXAREACAR                       21.782 LAYER ME2 ;
 ANTENNAMAXAREACAR                       24.449 LAYER ME3 ;
 ANTENNAMAXAREACAR                       27.116 LAYER ME4 ;
END DI59
PIN DO59
  DIRECTION OUTPUT ;
 PORT
  LAYER ME4 ;
  RECT 278.385 0.000 278.705 0.600 ;
  LAYER ME3 ;
  RECT 278.385 0.000 278.705 0.600 ;
  LAYER ME2 ;
  RECT 278.385 0.000 278.705 0.600 ;
  LAYER ME1 ;
  RECT 278.385 0.000 278.705 0.600 ;
 END
 ANTENNAPARTIALMETALAREA                  5.273 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME3 ;
 ANTENNADIFFAREA                          1.293 LAYER ME4 ;
END DO59
PIN DI58
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 274.943 0.000 275.263 0.600 ;
  LAYER ME3 ;
  RECT 274.943 0.000 275.263 0.600 ;
  LAYER ME2 ;
  RECT 274.943 0.000 275.263 0.600 ;
  LAYER ME1 ;
  RECT 274.943 0.000 275.263 0.600 ;
 END
 ANTENNAPARTIALMETALAREA                  1.058 LAYER ME2 ;
 ANTENNAGATEAREA                          0.072 LAYER ME2 ;
 ANTENNAGATEAREA                          0.072 LAYER ME3 ;
 ANTENNAGATEAREA                          0.072 LAYER ME4 ;
 ANTENNADIFFAREA                          0.160 LAYER ME2 ;
 ANTENNADIFFAREA                          0.160 LAYER ME3 ;
 ANTENNADIFFAREA                          0.160 LAYER ME4 ;
 ANTENNAMAXAREACAR                       21.782 LAYER ME2 ;
 ANTENNAMAXAREACAR                       24.449 LAYER ME3 ;
 ANTENNAMAXAREACAR                       27.116 LAYER ME4 ;
END DI58
PIN DO58
  DIRECTION OUTPUT ;
 PORT
  LAYER ME4 ;
  RECT 274.381 0.000 274.701 0.600 ;
  LAYER ME3 ;
  RECT 274.381 0.000 274.701 0.600 ;
  LAYER ME2 ;
  RECT 274.381 0.000 274.701 0.600 ;
  LAYER ME1 ;
  RECT 274.381 0.000 274.701 0.600 ;
 END
 ANTENNAPARTIALMETALAREA                  5.273 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME3 ;
 ANTENNADIFFAREA                          1.293 LAYER ME4 ;
END DO58
PIN DI57
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 270.939 0.000 271.259 0.600 ;
  LAYER ME3 ;
  RECT 270.939 0.000 271.259 0.600 ;
  LAYER ME2 ;
  RECT 270.939 0.000 271.259 0.600 ;
  LAYER ME1 ;
  RECT 270.939 0.000 271.259 0.600 ;
 END
 ANTENNAPARTIALMETALAREA                  1.058 LAYER ME2 ;
 ANTENNAGATEAREA                          0.072 LAYER ME2 ;
 ANTENNAGATEAREA                          0.072 LAYER ME3 ;
 ANTENNAGATEAREA                          0.072 LAYER ME4 ;
 ANTENNADIFFAREA                          0.160 LAYER ME2 ;
 ANTENNADIFFAREA                          0.160 LAYER ME3 ;
 ANTENNADIFFAREA                          0.160 LAYER ME4 ;
 ANTENNAMAXAREACAR                       21.782 LAYER ME2 ;
 ANTENNAMAXAREACAR                       24.449 LAYER ME3 ;
 ANTENNAMAXAREACAR                       27.116 LAYER ME4 ;
END DI57
PIN DO57
  DIRECTION OUTPUT ;
 PORT
  LAYER ME4 ;
  RECT 270.377 0.000 270.697 0.600 ;
  LAYER ME3 ;
  RECT 270.377 0.000 270.697 0.600 ;
  LAYER ME2 ;
  RECT 270.377 0.000 270.697 0.600 ;
  LAYER ME1 ;
  RECT 270.377 0.000 270.697 0.600 ;
 END
 ANTENNAPARTIALMETALAREA                  5.273 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME3 ;
 ANTENNADIFFAREA                          1.293 LAYER ME4 ;
END DO57
PIN DI56
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 266.935 0.000 267.255 0.600 ;
  LAYER ME3 ;
  RECT 266.935 0.000 267.255 0.600 ;
  LAYER ME2 ;
  RECT 266.935 0.000 267.255 0.600 ;
  LAYER ME1 ;
  RECT 266.935 0.000 267.255 0.600 ;
 END
 ANTENNAPARTIALMETALAREA                  1.058 LAYER ME2 ;
 ANTENNAGATEAREA                          0.072 LAYER ME2 ;
 ANTENNAGATEAREA                          0.072 LAYER ME3 ;
 ANTENNAGATEAREA                          0.072 LAYER ME4 ;
 ANTENNADIFFAREA                          0.160 LAYER ME2 ;
 ANTENNADIFFAREA                          0.160 LAYER ME3 ;
 ANTENNADIFFAREA                          0.160 LAYER ME4 ;
 ANTENNAMAXAREACAR                       21.782 LAYER ME2 ;
 ANTENNAMAXAREACAR                       24.449 LAYER ME3 ;
 ANTENNAMAXAREACAR                       27.116 LAYER ME4 ;
END DI56
PIN DO56
  DIRECTION OUTPUT ;
 PORT
  LAYER ME4 ;
  RECT 266.373 0.000 266.693 0.600 ;
  LAYER ME3 ;
  RECT 266.373 0.000 266.693 0.600 ;
  LAYER ME2 ;
  RECT 266.373 0.000 266.693 0.600 ;
  LAYER ME1 ;
  RECT 266.373 0.000 266.693 0.600 ;
 END
 ANTENNAPARTIALMETALAREA                  5.273 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME3 ;
 ANTENNADIFFAREA                          1.293 LAYER ME4 ;
END DO56
PIN DI55
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 262.931 0.000 263.251 0.600 ;
  LAYER ME3 ;
  RECT 262.931 0.000 263.251 0.600 ;
  LAYER ME2 ;
  RECT 262.931 0.000 263.251 0.600 ;
  LAYER ME1 ;
  RECT 262.931 0.000 263.251 0.600 ;
 END
 ANTENNAPARTIALMETALAREA                  1.058 LAYER ME2 ;
 ANTENNAGATEAREA                          0.072 LAYER ME2 ;
 ANTENNAGATEAREA                          0.072 LAYER ME3 ;
 ANTENNAGATEAREA                          0.072 LAYER ME4 ;
 ANTENNADIFFAREA                          0.160 LAYER ME2 ;
 ANTENNADIFFAREA                          0.160 LAYER ME3 ;
 ANTENNADIFFAREA                          0.160 LAYER ME4 ;
 ANTENNAMAXAREACAR                       21.782 LAYER ME2 ;
 ANTENNAMAXAREACAR                       24.449 LAYER ME3 ;
 ANTENNAMAXAREACAR                       27.116 LAYER ME4 ;
END DI55
PIN DO55
  DIRECTION OUTPUT ;
 PORT
  LAYER ME4 ;
  RECT 262.369 0.000 262.689 0.600 ;
  LAYER ME3 ;
  RECT 262.369 0.000 262.689 0.600 ;
  LAYER ME2 ;
  RECT 262.369 0.000 262.689 0.600 ;
  LAYER ME1 ;
  RECT 262.369 0.000 262.689 0.600 ;
 END
 ANTENNAPARTIALMETALAREA                  5.273 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME3 ;
 ANTENNADIFFAREA                          1.293 LAYER ME4 ;
END DO55
PIN DI54
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 258.927 0.000 259.247 0.600 ;
  LAYER ME3 ;
  RECT 258.927 0.000 259.247 0.600 ;
  LAYER ME2 ;
  RECT 258.927 0.000 259.247 0.600 ;
  LAYER ME1 ;
  RECT 258.927 0.000 259.247 0.600 ;
 END
 ANTENNAPARTIALMETALAREA                  1.058 LAYER ME2 ;
 ANTENNAGATEAREA                          0.072 LAYER ME2 ;
 ANTENNAGATEAREA                          0.072 LAYER ME3 ;
 ANTENNAGATEAREA                          0.072 LAYER ME4 ;
 ANTENNADIFFAREA                          0.160 LAYER ME2 ;
 ANTENNADIFFAREA                          0.160 LAYER ME3 ;
 ANTENNADIFFAREA                          0.160 LAYER ME4 ;
 ANTENNAMAXAREACAR                       21.782 LAYER ME2 ;
 ANTENNAMAXAREACAR                       24.449 LAYER ME3 ;
 ANTENNAMAXAREACAR                       27.116 LAYER ME4 ;
END DI54
PIN DO54
  DIRECTION OUTPUT ;
 PORT
  LAYER ME4 ;
  RECT 258.365 0.000 258.685 0.600 ;
  LAYER ME3 ;
  RECT 258.365 0.000 258.685 0.600 ;
  LAYER ME2 ;
  RECT 258.365 0.000 258.685 0.600 ;
  LAYER ME1 ;
  RECT 258.365 0.000 258.685 0.600 ;
 END
 ANTENNAPARTIALMETALAREA                  5.273 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME3 ;
 ANTENNADIFFAREA                          1.293 LAYER ME4 ;
END DO54
PIN DI53
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 254.923 0.000 255.243 0.600 ;
  LAYER ME3 ;
  RECT 254.923 0.000 255.243 0.600 ;
  LAYER ME2 ;
  RECT 254.923 0.000 255.243 0.600 ;
  LAYER ME1 ;
  RECT 254.923 0.000 255.243 0.600 ;
 END
 ANTENNAPARTIALMETALAREA                  1.058 LAYER ME2 ;
 ANTENNAGATEAREA                          0.072 LAYER ME2 ;
 ANTENNAGATEAREA                          0.072 LAYER ME3 ;
 ANTENNAGATEAREA                          0.072 LAYER ME4 ;
 ANTENNADIFFAREA                          0.160 LAYER ME2 ;
 ANTENNADIFFAREA                          0.160 LAYER ME3 ;
 ANTENNADIFFAREA                          0.160 LAYER ME4 ;
 ANTENNAMAXAREACAR                       21.782 LAYER ME2 ;
 ANTENNAMAXAREACAR                       24.449 LAYER ME3 ;
 ANTENNAMAXAREACAR                       27.116 LAYER ME4 ;
END DI53
PIN DO53
  DIRECTION OUTPUT ;
 PORT
  LAYER ME4 ;
  RECT 254.361 0.000 254.681 0.600 ;
  LAYER ME3 ;
  RECT 254.361 0.000 254.681 0.600 ;
  LAYER ME2 ;
  RECT 254.361 0.000 254.681 0.600 ;
  LAYER ME1 ;
  RECT 254.361 0.000 254.681 0.600 ;
 END
 ANTENNAPARTIALMETALAREA                  5.273 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME3 ;
 ANTENNADIFFAREA                          1.293 LAYER ME4 ;
END DO53
PIN DI52
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 250.919 0.000 251.239 0.600 ;
  LAYER ME3 ;
  RECT 250.919 0.000 251.239 0.600 ;
  LAYER ME2 ;
  RECT 250.919 0.000 251.239 0.600 ;
  LAYER ME1 ;
  RECT 250.919 0.000 251.239 0.600 ;
 END
 ANTENNAPARTIALMETALAREA                  1.058 LAYER ME2 ;
 ANTENNAGATEAREA                          0.072 LAYER ME2 ;
 ANTENNAGATEAREA                          0.072 LAYER ME3 ;
 ANTENNAGATEAREA                          0.072 LAYER ME4 ;
 ANTENNADIFFAREA                          0.160 LAYER ME2 ;
 ANTENNADIFFAREA                          0.160 LAYER ME3 ;
 ANTENNADIFFAREA                          0.160 LAYER ME4 ;
 ANTENNAMAXAREACAR                       21.782 LAYER ME2 ;
 ANTENNAMAXAREACAR                       24.449 LAYER ME3 ;
 ANTENNAMAXAREACAR                       27.116 LAYER ME4 ;
END DI52
PIN DO52
  DIRECTION OUTPUT ;
 PORT
  LAYER ME4 ;
  RECT 250.357 0.000 250.677 0.600 ;
  LAYER ME3 ;
  RECT 250.357 0.000 250.677 0.600 ;
  LAYER ME2 ;
  RECT 250.357 0.000 250.677 0.600 ;
  LAYER ME1 ;
  RECT 250.357 0.000 250.677 0.600 ;
 END
 ANTENNAPARTIALMETALAREA                  5.273 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME3 ;
 ANTENNADIFFAREA                          1.293 LAYER ME4 ;
END DO52
PIN DI51
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 246.915 0.000 247.235 0.600 ;
  LAYER ME3 ;
  RECT 246.915 0.000 247.235 0.600 ;
  LAYER ME2 ;
  RECT 246.915 0.000 247.235 0.600 ;
  LAYER ME1 ;
  RECT 246.915 0.000 247.235 0.600 ;
 END
 ANTENNAPARTIALMETALAREA                  1.058 LAYER ME2 ;
 ANTENNAGATEAREA                          0.072 LAYER ME2 ;
 ANTENNAGATEAREA                          0.072 LAYER ME3 ;
 ANTENNAGATEAREA                          0.072 LAYER ME4 ;
 ANTENNADIFFAREA                          0.160 LAYER ME2 ;
 ANTENNADIFFAREA                          0.160 LAYER ME3 ;
 ANTENNADIFFAREA                          0.160 LAYER ME4 ;
 ANTENNAMAXAREACAR                       21.782 LAYER ME2 ;
 ANTENNAMAXAREACAR                       24.449 LAYER ME3 ;
 ANTENNAMAXAREACAR                       27.116 LAYER ME4 ;
END DI51
PIN DO51
  DIRECTION OUTPUT ;
 PORT
  LAYER ME4 ;
  RECT 246.353 0.000 246.673 0.600 ;
  LAYER ME3 ;
  RECT 246.353 0.000 246.673 0.600 ;
  LAYER ME2 ;
  RECT 246.353 0.000 246.673 0.600 ;
  LAYER ME1 ;
  RECT 246.353 0.000 246.673 0.600 ;
 END
 ANTENNAPARTIALMETALAREA                  5.273 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME3 ;
 ANTENNADIFFAREA                          1.293 LAYER ME4 ;
END DO51
PIN DI50
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 242.911 0.000 243.231 0.600 ;
  LAYER ME3 ;
  RECT 242.911 0.000 243.231 0.600 ;
  LAYER ME2 ;
  RECT 242.911 0.000 243.231 0.600 ;
  LAYER ME1 ;
  RECT 242.911 0.000 243.231 0.600 ;
 END
 ANTENNAPARTIALMETALAREA                  1.058 LAYER ME2 ;
 ANTENNAGATEAREA                          0.072 LAYER ME2 ;
 ANTENNAGATEAREA                          0.072 LAYER ME3 ;
 ANTENNAGATEAREA                          0.072 LAYER ME4 ;
 ANTENNADIFFAREA                          0.160 LAYER ME2 ;
 ANTENNADIFFAREA                          0.160 LAYER ME3 ;
 ANTENNADIFFAREA                          0.160 LAYER ME4 ;
 ANTENNAMAXAREACAR                       21.782 LAYER ME2 ;
 ANTENNAMAXAREACAR                       24.449 LAYER ME3 ;
 ANTENNAMAXAREACAR                       27.116 LAYER ME4 ;
END DI50
PIN DO50
  DIRECTION OUTPUT ;
 PORT
  LAYER ME4 ;
  RECT 242.349 0.000 242.669 0.600 ;
  LAYER ME3 ;
  RECT 242.349 0.000 242.669 0.600 ;
  LAYER ME2 ;
  RECT 242.349 0.000 242.669 0.600 ;
  LAYER ME1 ;
  RECT 242.349 0.000 242.669 0.600 ;
 END
 ANTENNAPARTIALMETALAREA                  5.273 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME3 ;
 ANTENNADIFFAREA                          1.293 LAYER ME4 ;
END DO50
PIN DI49
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 238.907 0.000 239.227 0.600 ;
  LAYER ME3 ;
  RECT 238.907 0.000 239.227 0.600 ;
  LAYER ME2 ;
  RECT 238.907 0.000 239.227 0.600 ;
  LAYER ME1 ;
  RECT 238.907 0.000 239.227 0.600 ;
 END
 ANTENNAPARTIALMETALAREA                  1.058 LAYER ME2 ;
 ANTENNAGATEAREA                          0.072 LAYER ME2 ;
 ANTENNAGATEAREA                          0.072 LAYER ME3 ;
 ANTENNAGATEAREA                          0.072 LAYER ME4 ;
 ANTENNADIFFAREA                          0.160 LAYER ME2 ;
 ANTENNADIFFAREA                          0.160 LAYER ME3 ;
 ANTENNADIFFAREA                          0.160 LAYER ME4 ;
 ANTENNAMAXAREACAR                       21.782 LAYER ME2 ;
 ANTENNAMAXAREACAR                       24.449 LAYER ME3 ;
 ANTENNAMAXAREACAR                       27.116 LAYER ME4 ;
END DI49
PIN DO49
  DIRECTION OUTPUT ;
 PORT
  LAYER ME4 ;
  RECT 238.345 0.000 238.665 0.600 ;
  LAYER ME3 ;
  RECT 238.345 0.000 238.665 0.600 ;
  LAYER ME2 ;
  RECT 238.345 0.000 238.665 0.600 ;
  LAYER ME1 ;
  RECT 238.345 0.000 238.665 0.600 ;
 END
 ANTENNAPARTIALMETALAREA                  5.273 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME3 ;
 ANTENNADIFFAREA                          1.293 LAYER ME4 ;
END DO49
PIN DI48
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 234.341 0.000 234.661 0.600 ;
  LAYER ME3 ;
  RECT 234.341 0.000 234.661 0.600 ;
  LAYER ME2 ;
  RECT 234.341 0.000 234.661 0.600 ;
  LAYER ME1 ;
  RECT 234.341 0.000 234.661 0.600 ;
 END
 ANTENNAPARTIALMETALAREA                  0.346 LAYER ME1 ;
 ANTENNAPARTIALMETALAREA                  1.466 LAYER ME2 ;
 ANTENNAPARTIALMETALAREA                  0.508 LAYER ME3 ;
 ANTENNAGATEAREA                          0.072 LAYER ME3 ;
 ANTENNAGATEAREA                          0.072 LAYER ME4 ;
 ANTENNADIFFAREA                          0.218 LAYER ME1 ;
 ANTENNADIFFAREA                          0.218 LAYER ME2 ;
 ANTENNADIFFAREA                          0.218 LAYER ME3 ;
 ANTENNADIFFAREA                          0.218 LAYER ME4 ;
 ANTENNAMAXAREACAR                       17.267 LAYER ME3 ;
 ANTENNAMAXAREACAR                       19.933 LAYER ME4 ;
END DI48
PIN DO48
  DIRECTION OUTPUT ;
 PORT
  LAYER ME4 ;
  RECT 234.903 0.000 235.223 0.600 ;
  LAYER ME3 ;
  RECT 234.903 0.000 235.223 0.600 ;
  LAYER ME2 ;
  RECT 234.903 0.000 235.223 0.600 ;
  LAYER ME1 ;
  RECT 234.903 0.000 235.223 0.600 ;
 END
 ANTENNAPARTIALMETALAREA                  5.602 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME3 ;
 ANTENNADIFFAREA                          1.293 LAYER ME4 ;
END DO48
PIN WEB4
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 232.901 0.000 233.221 0.600 ;
  LAYER ME3 ;
  RECT 232.901 0.000 233.221 0.600 ;
  LAYER ME2 ;
  RECT 232.901 0.000 233.221 0.600 ;
  LAYER ME1 ;
  RECT 232.901 0.000 233.221 0.600 ;
 END
 ANTENNAPARTIALMETALAREA                  1.036 LAYER ME2 ;
 ANTENNAGATEAREA                          0.288 LAYER ME2 ;
 ANTENNAGATEAREA                          0.288 LAYER ME3 ;
 ANTENNAGATEAREA                          0.288 LAYER ME4 ;
 ANTENNADIFFAREA                          0.206 LAYER ME2 ;
 ANTENNADIFFAREA                          0.206 LAYER ME3 ;
 ANTENNADIFFAREA                          0.206 LAYER ME4 ;
 ANTENNAMAXAREACAR                        5.844 LAYER ME2 ;
 ANTENNAMAXAREACAR                        6.511 LAYER ME3 ;
 ANTENNAMAXAREACAR                        7.178 LAYER ME4 ;
END WEB4
OBS
  LAYER ME3 SPACING 0.260 ;
  RECT 0.000 0.000 427.883 80.703 ;
  LAYER ME2 SPACING 0.260 ;
  RECT 0.000 0.000 427.883 80.703 ;
  LAYER ME1 SPACING 0.260 ;
  RECT 0.000 0.000 427.883 80.703 ;
  LAYER ME4 SPACING 0.260 ;
  RECT 0.000 0.000 207.934 80.703 ;
  LAYER ME4 SPACING 0.260 ;
  RECT 209.588 0.000 210.708 80.703 ;
  LAYER ME4 SPACING 0.260 ;
  RECT 212.303 0.000 213.023 80.703 ;
  LAYER ME4 SPACING 0.260 ;
  RECT 213.753 0.000 214.473 80.703 ;
  LAYER ME4 SPACING 0.260 ;
  RECT 216.533 0.000 217.133 80.703 ;
  LAYER ME4 SPACING 0.260 ;
  RECT 219.747 0.000 221.433 80.703 ;
  LAYER ME4 SPACING 0.260 ;
  RECT 222.823 0.000 223.943 80.703 ;
  LAYER ME4 SPACING 0.260 ;
  RECT 225.218 0.000 225.938 80.703 ;
  LAYER ME4 SPACING 0.260 ;
  RECT 226.933 0.000 227.653 80.703 ;
  LAYER ME4 SPACING 0.260 ;
  RECT 228.853 0.000 427.883 80.703 ;
END
END SYKB110_64X12X8CM2
END LIBRARY





