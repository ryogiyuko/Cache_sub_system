# ________________________________________________________________________________________________
# 
# 
#             Synchronous High-Density Single-Port SRAM Compiler
# 
#                 UMC 0.11um LL AE Logic Process
# 
# ________________________________________________________________________________________________
# 
#               
#         Copyright (C) 2024 Faraday Technology Corporation. All Rights Reserved.       
#                
#         This source code is an unpublished work belongs to Faraday Technology Corporation       
#         It is considered a trade secret and is not to be divulged or       
#         used by parties who have not received written authorization from       
#         Faraday Technology Corporation       
#                
#         Faraday's home page can be found at: http://www.faraday-tech.com/       
#                
# ________________________________________________________________________________________________
# 
#        IP Name            :  FSR0K_D_SH                
#        IP Version         :  1.3.0                     
#        IP Release Status  :  Active                    
#        Word               :  4224                      
#        Bit                :  8                         
#        Byte               :  16                        
#        Mux                :  1                         
#        Output Loading     :  0.01                      
#        Clock Input Slew   :  0.016                     
#        Data Input Slew    :  0.016                     
#        Ring Type          :  Ring Shape Model          
#        Ring Width         :  2                         
#        Bus Format         :  0                         
#        Memaker Path       :  /home/mem/Desktop/memlib  
#        GUI Version        :  m20230904                 
#        Date               :  2024/12/23 09:47:17       
# ________________________________________________________________________________________________
# 

VERSION 5.5 ;
NAMESCASESENSITIVE ON ;
MACRO SHKD110_4224X8X16BM1
CLASS BLOCK ;
FOREIGN SHKD110_4224X8X16BM1 0.000 0.000 ;
ORIGIN 0.000 0.000 ;
SIZE 2692.940 BY 565.930 ;
SYMMETRY x y r90 ;
SITE core ;
PIN DO127
  DIRECTION OUTPUT ;
 PORT
  LAYER ME4 ;
  RECT 2680.800 0.000 2681.600 1.000 ;
  LAYER ME3 ;
  RECT 2680.800 0.000 2681.600 1.000 ;
  LAYER ME2 ;
  RECT 2680.800 0.000 2681.600 1.000 ;
  LAYER ME1 ;
  RECT 2680.800 0.000 2681.600 1.000 ;
 END
 ANTENNAPARTIALMETALAREA                  4.176 LAYER ME2 ;
 ANTENNADIFFAREA                          5.472 LAYER ME2 ;
 ANTENNADIFFAREA                          5.472 LAYER ME3 ;
 ANTENNADIFFAREA                          5.472 LAYER ME4 ;
END DO127
PIN DI127
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 2666.400 0.000 2667.200 1.000 ;
  LAYER ME3 ;
  RECT 2666.400 0.000 2667.200 1.000 ;
  LAYER ME2 ;
  RECT 2666.400 0.000 2667.200 1.000 ;
  LAYER ME1 ;
  RECT 2666.400 0.000 2667.200 1.000 ;
 END
 ANTENNAPARTIALMETALAREA                  3.126 LAYER ME2 ;
 ANTENNAGATEAREA                          0.086 LAYER ME2 ;
 ANTENNAGATEAREA                          0.086 LAYER ME3 ;
 ANTENNAGATEAREA                          0.086 LAYER ME4 ;
 ANTENNADIFFAREA                          0.160 LAYER ME2 ;
 ANTENNADIFFAREA                          0.160 LAYER ME3 ;
 ANTENNADIFFAREA                          0.160 LAYER ME4 ;
 ANTENNAMAXAREACAR                       48.523 LAYER ME2 ;
 ANTENNAMAXAREACAR                       57.782 LAYER ME3 ;
 ANTENNAMAXAREACAR                       67.042 LAYER ME4 ;
END DI127
PIN DO126
  DIRECTION OUTPUT ;
 PORT
  LAYER ME4 ;
  RECT 2661.200 0.000 2662.000 1.000 ;
  LAYER ME3 ;
  RECT 2661.200 0.000 2662.000 1.000 ;
  LAYER ME2 ;
  RECT 2661.200 0.000 2662.000 1.000 ;
  LAYER ME1 ;
  RECT 2661.200 0.000 2662.000 1.000 ;
 END
 ANTENNAPARTIALMETALAREA                  4.152 LAYER ME2 ;
 ANTENNADIFFAREA                          5.472 LAYER ME2 ;
 ANTENNADIFFAREA                          5.472 LAYER ME3 ;
 ANTENNADIFFAREA                          5.472 LAYER ME4 ;
END DO126
PIN DI126
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 2646.400 0.000 2647.200 1.000 ;
  LAYER ME3 ;
  RECT 2646.400 0.000 2647.200 1.000 ;
  LAYER ME2 ;
  RECT 2646.400 0.000 2647.200 1.000 ;
  LAYER ME1 ;
  RECT 2646.400 0.000 2647.200 1.000 ;
 END
 ANTENNAPARTIALMETALAREA                  3.138 LAYER ME2 ;
 ANTENNAGATEAREA                          0.086 LAYER ME2 ;
 ANTENNAGATEAREA                          0.086 LAYER ME3 ;
 ANTENNAGATEAREA                          0.086 LAYER ME4 ;
 ANTENNADIFFAREA                          0.160 LAYER ME2 ;
 ANTENNADIFFAREA                          0.160 LAYER ME3 ;
 ANTENNADIFFAREA                          0.160 LAYER ME4 ;
 ANTENNAMAXAREACAR                       48.662 LAYER ME2 ;
 ANTENNAMAXAREACAR                       57.921 LAYER ME3 ;
 ANTENNAMAXAREACAR                       67.181 LAYER ME4 ;
END DI126
PIN DO125
  DIRECTION OUTPUT ;
 PORT
  LAYER ME4 ;
  RECT 2640.000 0.000 2640.800 1.000 ;
  LAYER ME3 ;
  RECT 2640.000 0.000 2640.800 1.000 ;
  LAYER ME2 ;
  RECT 2640.000 0.000 2640.800 1.000 ;
  LAYER ME1 ;
  RECT 2640.000 0.000 2640.800 1.000 ;
 END
 ANTENNAPARTIALMETALAREA                  4.152 LAYER ME2 ;
 ANTENNADIFFAREA                          5.472 LAYER ME2 ;
 ANTENNADIFFAREA                          5.472 LAYER ME3 ;
 ANTENNADIFFAREA                          5.472 LAYER ME4 ;
END DO125
PIN DI125
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 2625.600 0.000 2626.400 1.000 ;
  LAYER ME3 ;
  RECT 2625.600 0.000 2626.400 1.000 ;
  LAYER ME2 ;
  RECT 2625.600 0.000 2626.400 1.000 ;
  LAYER ME1 ;
  RECT 2625.600 0.000 2626.400 1.000 ;
 END
 ANTENNAPARTIALMETALAREA                  3.150 LAYER ME2 ;
 ANTENNAGATEAREA                          0.086 LAYER ME2 ;
 ANTENNAGATEAREA                          0.086 LAYER ME3 ;
 ANTENNAGATEAREA                          0.086 LAYER ME4 ;
 ANTENNADIFFAREA                          0.160 LAYER ME2 ;
 ANTENNADIFFAREA                          0.160 LAYER ME3 ;
 ANTENNADIFFAREA                          0.160 LAYER ME4 ;
 ANTENNAMAXAREACAR                       48.801 LAYER ME2 ;
 ANTENNAMAXAREACAR                       58.060 LAYER ME3 ;
 ANTENNAMAXAREACAR                       67.319 LAYER ME4 ;
END DI125
PIN DO124
  DIRECTION OUTPUT ;
 PORT
  LAYER ME4 ;
  RECT 2620.400 0.000 2621.200 1.000 ;
  LAYER ME3 ;
  RECT 2620.400 0.000 2621.200 1.000 ;
  LAYER ME2 ;
  RECT 2620.400 0.000 2621.200 1.000 ;
  LAYER ME1 ;
  RECT 2620.400 0.000 2621.200 1.000 ;
 END
 ANTENNAPARTIALMETALAREA                  4.176 LAYER ME2 ;
 ANTENNADIFFAREA                          5.472 LAYER ME2 ;
 ANTENNADIFFAREA                          5.472 LAYER ME3 ;
 ANTENNADIFFAREA                          5.472 LAYER ME4 ;
END DO124
PIN DI124
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 2605.600 0.000 2606.400 1.000 ;
  LAYER ME3 ;
  RECT 2605.600 0.000 2606.400 1.000 ;
  LAYER ME2 ;
  RECT 2605.600 0.000 2606.400 1.000 ;
  LAYER ME1 ;
  RECT 2605.600 0.000 2606.400 1.000 ;
 END
 ANTENNAPARTIALMETALAREA                  3.118 LAYER ME2 ;
 ANTENNAGATEAREA                          0.086 LAYER ME2 ;
 ANTENNAGATEAREA                          0.086 LAYER ME3 ;
 ANTENNAGATEAREA                          0.086 LAYER ME4 ;
 ANTENNADIFFAREA                          0.160 LAYER ME2 ;
 ANTENNADIFFAREA                          0.160 LAYER ME3 ;
 ANTENNADIFFAREA                          0.160 LAYER ME4 ;
 ANTENNAMAXAREACAR                       48.431 LAYER ME2 ;
 ANTENNAMAXAREACAR                       57.690 LAYER ME3 ;
 ANTENNAMAXAREACAR                       66.949 LAYER ME4 ;
END DI124
PIN DO123
  DIRECTION OUTPUT ;
 PORT
  LAYER ME4 ;
  RECT 2599.200 0.000 2600.000 1.000 ;
  LAYER ME3 ;
  RECT 2599.200 0.000 2600.000 1.000 ;
  LAYER ME2 ;
  RECT 2599.200 0.000 2600.000 1.000 ;
  LAYER ME1 ;
  RECT 2599.200 0.000 2600.000 1.000 ;
 END
 ANTENNAPARTIALMETALAREA                  4.152 LAYER ME2 ;
 ANTENNADIFFAREA                          5.472 LAYER ME2 ;
 ANTENNADIFFAREA                          5.472 LAYER ME3 ;
 ANTENNADIFFAREA                          5.472 LAYER ME4 ;
END DO123
PIN DI123
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 2584.400 0.000 2585.200 1.000 ;
  LAYER ME3 ;
  RECT 2584.400 0.000 2585.200 1.000 ;
  LAYER ME2 ;
  RECT 2584.400 0.000 2585.200 1.000 ;
  LAYER ME1 ;
  RECT 2584.400 0.000 2585.200 1.000 ;
 END
 ANTENNAPARTIALMETALAREA                  3.138 LAYER ME2 ;
 ANTENNAGATEAREA                          0.086 LAYER ME2 ;
 ANTENNAGATEAREA                          0.086 LAYER ME3 ;
 ANTENNAGATEAREA                          0.086 LAYER ME4 ;
 ANTENNADIFFAREA                          0.160 LAYER ME2 ;
 ANTENNADIFFAREA                          0.160 LAYER ME3 ;
 ANTENNADIFFAREA                          0.160 LAYER ME4 ;
 ANTENNAMAXAREACAR                       48.662 LAYER ME2 ;
 ANTENNAMAXAREACAR                       57.921 LAYER ME3 ;
 ANTENNAMAXAREACAR                       67.181 LAYER ME4 ;
END DI123
PIN DO122
  DIRECTION OUTPUT ;
 PORT
  LAYER ME4 ;
  RECT 2579.200 0.000 2580.000 1.000 ;
  LAYER ME3 ;
  RECT 2579.200 0.000 2580.000 1.000 ;
  LAYER ME2 ;
  RECT 2579.200 0.000 2580.000 1.000 ;
  LAYER ME1 ;
  RECT 2579.200 0.000 2580.000 1.000 ;
 END
 ANTENNAPARTIALMETALAREA                  4.160 LAYER ME2 ;
 ANTENNADIFFAREA                          5.472 LAYER ME2 ;
 ANTENNADIFFAREA                          5.472 LAYER ME3 ;
 ANTENNADIFFAREA                          5.472 LAYER ME4 ;
END DO122
PIN DI122
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 2564.800 0.000 2565.600 1.000 ;
  LAYER ME3 ;
  RECT 2564.800 0.000 2565.600 1.000 ;
  LAYER ME2 ;
  RECT 2564.800 0.000 2565.600 1.000 ;
  LAYER ME1 ;
  RECT 2564.800 0.000 2565.600 1.000 ;
 END
 ANTENNAPARTIALMETALAREA                  3.142 LAYER ME2 ;
 ANTENNAGATEAREA                          0.086 LAYER ME2 ;
 ANTENNAGATEAREA                          0.086 LAYER ME3 ;
 ANTENNAGATEAREA                          0.086 LAYER ME4 ;
 ANTENNADIFFAREA                          0.160 LAYER ME2 ;
 ANTENNADIFFAREA                          0.160 LAYER ME3 ;
 ANTENNADIFFAREA                          0.160 LAYER ME4 ;
 ANTENNAMAXAREACAR                       48.708 LAYER ME2 ;
 ANTENNAMAXAREACAR                       57.968 LAYER ME3 ;
 ANTENNAMAXAREACAR                       67.227 LAYER ME4 ;
END DI122
PIN DO121
  DIRECTION OUTPUT ;
 PORT
  LAYER ME4 ;
  RECT 2558.400 0.000 2559.200 1.000 ;
  LAYER ME3 ;
  RECT 2558.400 0.000 2559.200 1.000 ;
  LAYER ME2 ;
  RECT 2558.400 0.000 2559.200 1.000 ;
  LAYER ME1 ;
  RECT 2558.400 0.000 2559.200 1.000 ;
 END
 ANTENNAPARTIALMETALAREA                  4.176 LAYER ME2 ;
 ANTENNADIFFAREA                          5.472 LAYER ME2 ;
 ANTENNADIFFAREA                          5.472 LAYER ME3 ;
 ANTENNADIFFAREA                          5.472 LAYER ME4 ;
END DO121
PIN DI121
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 2543.600 0.000 2544.400 1.000 ;
  LAYER ME3 ;
  RECT 2543.600 0.000 2544.400 1.000 ;
  LAYER ME2 ;
  RECT 2543.600 0.000 2544.400 1.000 ;
  LAYER ME1 ;
  RECT 2543.600 0.000 2544.400 1.000 ;
 END
 ANTENNAPARTIALMETALAREA                  3.118 LAYER ME2 ;
 ANTENNAGATEAREA                          0.086 LAYER ME2 ;
 ANTENNAGATEAREA                          0.086 LAYER ME3 ;
 ANTENNAGATEAREA                          0.086 LAYER ME4 ;
 ANTENNADIFFAREA                          0.160 LAYER ME2 ;
 ANTENNADIFFAREA                          0.160 LAYER ME3 ;
 ANTENNADIFFAREA                          0.160 LAYER ME4 ;
 ANTENNAMAXAREACAR                       48.431 LAYER ME2 ;
 ANTENNAMAXAREACAR                       57.690 LAYER ME3 ;
 ANTENNAMAXAREACAR                       66.949 LAYER ME4 ;
END DI121
PIN DO120
  DIRECTION OUTPUT ;
 PORT
  LAYER ME4 ;
  RECT 2538.400 0.000 2539.200 1.000 ;
  LAYER ME3 ;
  RECT 2538.400 0.000 2539.200 1.000 ;
  LAYER ME2 ;
  RECT 2538.400 0.000 2539.200 1.000 ;
  LAYER ME1 ;
  RECT 2538.400 0.000 2539.200 1.000 ;
 END
 ANTENNAPARTIALMETALAREA                  4.144 LAYER ME2 ;
 ANTENNADIFFAREA                          5.472 LAYER ME2 ;
 ANTENNADIFFAREA                          5.472 LAYER ME3 ;
 ANTENNADIFFAREA                          5.472 LAYER ME4 ;
END DO120
PIN WEB15
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 2525.600 0.000 2526.400 1.000 ;
  LAYER ME3 ;
  RECT 2525.600 0.000 2526.400 1.000 ;
  LAYER ME2 ;
  RECT 2525.600 0.000 2526.400 1.000 ;
  LAYER ME1 ;
  RECT 2525.600 0.000 2526.400 1.000 ;
 END
 ANTENNAPARTIALMETALAREA                  2.856 LAYER ME2 ;
 ANTENNAGATEAREA                          0.072 LAYER ME2 ;
 ANTENNAGATEAREA                          0.072 LAYER ME3 ;
 ANTENNAGATEAREA                          0.072 LAYER ME4 ;
 ANTENNADIFFAREA                          0.160 LAYER ME2 ;
 ANTENNADIFFAREA                          0.160 LAYER ME3 ;
 ANTENNADIFFAREA                          0.160 LAYER ME4 ;
 ANTENNAMAXAREACAR                       54.678 LAYER ME2 ;
 ANTENNAMAXAREACAR                       65.789 LAYER ME3 ;
 ANTENNAMAXAREACAR                       76.900 LAYER ME4 ;
END WEB15
PIN DI120
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 2523.600 0.000 2524.400 1.000 ;
  LAYER ME3 ;
  RECT 2523.600 0.000 2524.400 1.000 ;
  LAYER ME2 ;
  RECT 2523.600 0.000 2524.400 1.000 ;
  LAYER ME1 ;
  RECT 2523.600 0.000 2524.400 1.000 ;
 END
 ANTENNAPARTIALMETALAREA                  3.146 LAYER ME2 ;
 ANTENNAGATEAREA                          0.086 LAYER ME2 ;
 ANTENNAGATEAREA                          0.086 LAYER ME3 ;
 ANTENNAGATEAREA                          0.086 LAYER ME4 ;
 ANTENNADIFFAREA                          0.160 LAYER ME2 ;
 ANTENNADIFFAREA                          0.160 LAYER ME3 ;
 ANTENNADIFFAREA                          0.160 LAYER ME4 ;
 ANTENNAMAXAREACAR                       48.755 LAYER ME2 ;
 ANTENNAMAXAREACAR                       58.014 LAYER ME3 ;
 ANTENNAMAXAREACAR                       67.273 LAYER ME4 ;
END DI120
PIN DO119
  DIRECTION OUTPUT ;
 PORT
  LAYER ME4 ;
  RECT 2517.200 0.000 2518.000 1.000 ;
  LAYER ME3 ;
  RECT 2517.200 0.000 2518.000 1.000 ;
  LAYER ME2 ;
  RECT 2517.200 0.000 2518.000 1.000 ;
  LAYER ME1 ;
  RECT 2517.200 0.000 2518.000 1.000 ;
 END
 ANTENNAPARTIALMETALAREA                  4.160 LAYER ME2 ;
 ANTENNADIFFAREA                          5.472 LAYER ME2 ;
 ANTENNADIFFAREA                          5.472 LAYER ME3 ;
 ANTENNADIFFAREA                          5.472 LAYER ME4 ;
END DO119
PIN DI119
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 2502.800 0.000 2503.600 1.000 ;
  LAYER ME3 ;
  RECT 2502.800 0.000 2503.600 1.000 ;
  LAYER ME2 ;
  RECT 2502.800 0.000 2503.600 1.000 ;
  LAYER ME1 ;
  RECT 2502.800 0.000 2503.600 1.000 ;
 END
 ANTENNAPARTIALMETALAREA                  3.142 LAYER ME2 ;
 ANTENNAGATEAREA                          0.086 LAYER ME2 ;
 ANTENNAGATEAREA                          0.086 LAYER ME3 ;
 ANTENNAGATEAREA                          0.086 LAYER ME4 ;
 ANTENNADIFFAREA                          0.160 LAYER ME2 ;
 ANTENNADIFFAREA                          0.160 LAYER ME3 ;
 ANTENNADIFFAREA                          0.160 LAYER ME4 ;
 ANTENNAMAXAREACAR                       48.708 LAYER ME2 ;
 ANTENNAMAXAREACAR                       57.968 LAYER ME3 ;
 ANTENNAMAXAREACAR                       67.227 LAYER ME4 ;
END DI119
PIN DO118
  DIRECTION OUTPUT ;
 PORT
  LAYER ME4 ;
  RECT 2497.600 0.000 2498.400 1.000 ;
  LAYER ME3 ;
  RECT 2497.600 0.000 2498.400 1.000 ;
  LAYER ME2 ;
  RECT 2497.600 0.000 2498.400 1.000 ;
  LAYER ME1 ;
  RECT 2497.600 0.000 2498.400 1.000 ;
 END
 ANTENNAPARTIALMETALAREA                  4.168 LAYER ME2 ;
 ANTENNADIFFAREA                          5.472 LAYER ME2 ;
 ANTENNADIFFAREA                          5.472 LAYER ME3 ;
 ANTENNADIFFAREA                          5.472 LAYER ME4 ;
END DO118
PIN DI118
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 2482.800 0.000 2483.600 1.000 ;
  LAYER ME3 ;
  RECT 2482.800 0.000 2483.600 1.000 ;
  LAYER ME2 ;
  RECT 2482.800 0.000 2483.600 1.000 ;
  LAYER ME1 ;
  RECT 2482.800 0.000 2483.600 1.000 ;
 END
 ANTENNAPARTIALMETALAREA                  3.122 LAYER ME2 ;
 ANTENNAGATEAREA                          0.086 LAYER ME2 ;
 ANTENNAGATEAREA                          0.086 LAYER ME3 ;
 ANTENNAGATEAREA                          0.086 LAYER ME4 ;
 ANTENNADIFFAREA                          0.160 LAYER ME2 ;
 ANTENNADIFFAREA                          0.160 LAYER ME3 ;
 ANTENNADIFFAREA                          0.160 LAYER ME4 ;
 ANTENNAMAXAREACAR                       48.477 LAYER ME2 ;
 ANTENNAMAXAREACAR                       57.736 LAYER ME3 ;
 ANTENNAMAXAREACAR                       66.995 LAYER ME4 ;
END DI118
PIN DO117
  DIRECTION OUTPUT ;
 PORT
  LAYER ME4 ;
  RECT 2476.400 0.000 2477.200 1.000 ;
  LAYER ME3 ;
  RECT 2476.400 0.000 2477.200 1.000 ;
  LAYER ME2 ;
  RECT 2476.400 0.000 2477.200 1.000 ;
  LAYER ME1 ;
  RECT 2476.400 0.000 2477.200 1.000 ;
 END
 ANTENNAPARTIALMETALAREA                  4.144 LAYER ME2 ;
 ANTENNADIFFAREA                          5.472 LAYER ME2 ;
 ANTENNADIFFAREA                          5.472 LAYER ME3 ;
 ANTENNADIFFAREA                          5.472 LAYER ME4 ;
END DO117
PIN DI117
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 2461.600 0.000 2462.400 1.000 ;
  LAYER ME3 ;
  RECT 2461.600 0.000 2462.400 1.000 ;
  LAYER ME2 ;
  RECT 2461.600 0.000 2462.400 1.000 ;
  LAYER ME1 ;
  RECT 2461.600 0.000 2462.400 1.000 ;
 END
 ANTENNAPARTIALMETALAREA                  3.146 LAYER ME2 ;
 ANTENNAGATEAREA                          0.086 LAYER ME2 ;
 ANTENNAGATEAREA                          0.086 LAYER ME3 ;
 ANTENNAGATEAREA                          0.086 LAYER ME4 ;
 ANTENNADIFFAREA                          0.160 LAYER ME2 ;
 ANTENNADIFFAREA                          0.160 LAYER ME3 ;
 ANTENNADIFFAREA                          0.160 LAYER ME4 ;
 ANTENNAMAXAREACAR                       48.755 LAYER ME2 ;
 ANTENNAMAXAREACAR                       58.014 LAYER ME3 ;
 ANTENNAMAXAREACAR                       67.273 LAYER ME4 ;
END DI117
PIN DO116
  DIRECTION OUTPUT ;
 PORT
  LAYER ME4 ;
  RECT 2456.400 0.000 2457.200 1.000 ;
  LAYER ME3 ;
  RECT 2456.400 0.000 2457.200 1.000 ;
  LAYER ME2 ;
  RECT 2456.400 0.000 2457.200 1.000 ;
  LAYER ME1 ;
  RECT 2456.400 0.000 2457.200 1.000 ;
 END
 ANTENNAPARTIALMETALAREA                  4.168 LAYER ME2 ;
 ANTENNADIFFAREA                          5.472 LAYER ME2 ;
 ANTENNADIFFAREA                          5.472 LAYER ME3 ;
 ANTENNADIFFAREA                          5.472 LAYER ME4 ;
END DO116
PIN DI116
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 2442.000 0.000 2442.800 1.000 ;
  LAYER ME3 ;
  RECT 2442.000 0.000 2442.800 1.000 ;
  LAYER ME2 ;
  RECT 2442.000 0.000 2442.800 1.000 ;
  LAYER ME1 ;
  RECT 2442.000 0.000 2442.800 1.000 ;
 END
 ANTENNAPARTIALMETALAREA                  3.134 LAYER ME2 ;
 ANTENNAGATEAREA                          0.086 LAYER ME2 ;
 ANTENNAGATEAREA                          0.086 LAYER ME3 ;
 ANTENNAGATEAREA                          0.086 LAYER ME4 ;
 ANTENNADIFFAREA                          0.160 LAYER ME2 ;
 ANTENNADIFFAREA                          0.160 LAYER ME3 ;
 ANTENNADIFFAREA                          0.160 LAYER ME4 ;
 ANTENNAMAXAREACAR                       48.616 LAYER ME2 ;
 ANTENNAMAXAREACAR                       57.875 LAYER ME3 ;
 ANTENNAMAXAREACAR                       67.134 LAYER ME4 ;
END DI116
PIN DO115
  DIRECTION OUTPUT ;
 PORT
  LAYER ME4 ;
  RECT 2435.600 0.000 2436.400 1.000 ;
  LAYER ME3 ;
  RECT 2435.600 0.000 2436.400 1.000 ;
  LAYER ME2 ;
  RECT 2435.600 0.000 2436.400 1.000 ;
  LAYER ME1 ;
  RECT 2435.600 0.000 2436.400 1.000 ;
 END
 ANTENNAPARTIALMETALAREA                  4.168 LAYER ME2 ;
 ANTENNADIFFAREA                          5.472 LAYER ME2 ;
 ANTENNADIFFAREA                          5.472 LAYER ME3 ;
 ANTENNADIFFAREA                          5.472 LAYER ME4 ;
END DO115
PIN DI115
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 2420.800 0.000 2421.600 1.000 ;
  LAYER ME3 ;
  RECT 2420.800 0.000 2421.600 1.000 ;
  LAYER ME2 ;
  RECT 2420.800 0.000 2421.600 1.000 ;
  LAYER ME1 ;
  RECT 2420.800 0.000 2421.600 1.000 ;
 END
 ANTENNAPARTIALMETALAREA                  3.122 LAYER ME2 ;
 ANTENNAGATEAREA                          0.086 LAYER ME2 ;
 ANTENNAGATEAREA                          0.086 LAYER ME3 ;
 ANTENNAGATEAREA                          0.086 LAYER ME4 ;
 ANTENNADIFFAREA                          0.160 LAYER ME2 ;
 ANTENNADIFFAREA                          0.160 LAYER ME3 ;
 ANTENNADIFFAREA                          0.160 LAYER ME4 ;
 ANTENNAMAXAREACAR                       48.477 LAYER ME2 ;
 ANTENNAMAXAREACAR                       57.736 LAYER ME3 ;
 ANTENNAMAXAREACAR                       66.995 LAYER ME4 ;
END DI115
PIN DO114
  DIRECTION OUTPUT ;
 PORT
  LAYER ME4 ;
  RECT 2415.600 0.000 2416.400 1.000 ;
  LAYER ME3 ;
  RECT 2415.600 0.000 2416.400 1.000 ;
  LAYER ME2 ;
  RECT 2415.600 0.000 2416.400 1.000 ;
  LAYER ME1 ;
  RECT 2415.600 0.000 2416.400 1.000 ;
 END
 ANTENNAPARTIALMETALAREA                  4.144 LAYER ME2 ;
 ANTENNADIFFAREA                          5.472 LAYER ME2 ;
 ANTENNADIFFAREA                          5.472 LAYER ME3 ;
 ANTENNADIFFAREA                          5.472 LAYER ME4 ;
END DO114
PIN DI114
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 2400.800 0.000 2401.600 1.000 ;
  LAYER ME3 ;
  RECT 2400.800 0.000 2401.600 1.000 ;
  LAYER ME2 ;
  RECT 2400.800 0.000 2401.600 1.000 ;
  LAYER ME1 ;
  RECT 2400.800 0.000 2401.600 1.000 ;
 END
 ANTENNAPARTIALMETALAREA                  3.154 LAYER ME2 ;
 ANTENNAGATEAREA                          0.086 LAYER ME2 ;
 ANTENNAGATEAREA                          0.086 LAYER ME3 ;
 ANTENNAGATEAREA                          0.086 LAYER ME4 ;
 ANTENNADIFFAREA                          0.160 LAYER ME2 ;
 ANTENNADIFFAREA                          0.160 LAYER ME3 ;
 ANTENNADIFFAREA                          0.160 LAYER ME4 ;
 ANTENNAMAXAREACAR                       48.847 LAYER ME2 ;
 ANTENNAMAXAREACAR                       58.106 LAYER ME3 ;
 ANTENNAMAXAREACAR                       67.366 LAYER ME4 ;
END DI114
PIN DO113
  DIRECTION OUTPUT ;
 PORT
  LAYER ME4 ;
  RECT 2394.400 0.000 2395.200 1.000 ;
  LAYER ME3 ;
  RECT 2394.400 0.000 2395.200 1.000 ;
  LAYER ME2 ;
  RECT 2394.400 0.000 2395.200 1.000 ;
  LAYER ME1 ;
  RECT 2394.400 0.000 2395.200 1.000 ;
 END
 ANTENNAPARTIALMETALAREA                  4.168 LAYER ME2 ;
 ANTENNADIFFAREA                          5.472 LAYER ME2 ;
 ANTENNADIFFAREA                          5.472 LAYER ME3 ;
 ANTENNADIFFAREA                          5.472 LAYER ME4 ;
END DO113
PIN DI113
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 2380.000 0.000 2380.800 1.000 ;
  LAYER ME3 ;
  RECT 2380.000 0.000 2380.800 1.000 ;
  LAYER ME2 ;
  RECT 2380.000 0.000 2380.800 1.000 ;
  LAYER ME1 ;
  RECT 2380.000 0.000 2380.800 1.000 ;
 END
 ANTENNAPARTIALMETALAREA                  3.134 LAYER ME2 ;
 ANTENNAGATEAREA                          0.086 LAYER ME2 ;
 ANTENNAGATEAREA                          0.086 LAYER ME3 ;
 ANTENNAGATEAREA                          0.086 LAYER ME4 ;
 ANTENNADIFFAREA                          0.160 LAYER ME2 ;
 ANTENNADIFFAREA                          0.160 LAYER ME3 ;
 ANTENNADIFFAREA                          0.160 LAYER ME4 ;
 ANTENNAMAXAREACAR                       48.616 LAYER ME2 ;
 ANTENNAMAXAREACAR                       57.875 LAYER ME3 ;
 ANTENNAMAXAREACAR                       67.134 LAYER ME4 ;
END DI113
PIN DO112
  DIRECTION OUTPUT ;
 PORT
  LAYER ME4 ;
  RECT 2374.800 0.000 2375.600 1.000 ;
  LAYER ME3 ;
  RECT 2374.800 0.000 2375.600 1.000 ;
  LAYER ME2 ;
  RECT 2374.800 0.000 2375.600 1.000 ;
  LAYER ME1 ;
  RECT 2374.800 0.000 2375.600 1.000 ;
 END
 ANTENNAPARTIALMETALAREA                  4.160 LAYER ME2 ;
 ANTENNADIFFAREA                          5.472 LAYER ME2 ;
 ANTENNADIFFAREA                          5.472 LAYER ME3 ;
 ANTENNADIFFAREA                          5.472 LAYER ME4 ;
END DO112
PIN WEB14
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 2361.600 0.000 2362.400 1.000 ;
  LAYER ME3 ;
  RECT 2361.600 0.000 2362.400 1.000 ;
  LAYER ME2 ;
  RECT 2361.600 0.000 2362.400 1.000 ;
  LAYER ME1 ;
  RECT 2361.600 0.000 2362.400 1.000 ;
 END
 ANTENNAPARTIALMETALAREA                  2.868 LAYER ME2 ;
 ANTENNAGATEAREA                          0.072 LAYER ME2 ;
 ANTENNAGATEAREA                          0.072 LAYER ME3 ;
 ANTENNAGATEAREA                          0.072 LAYER ME4 ;
 ANTENNADIFFAREA                          0.160 LAYER ME2 ;
 ANTENNADIFFAREA                          0.160 LAYER ME3 ;
 ANTENNADIFFAREA                          0.160 LAYER ME4 ;
 ANTENNAMAXAREACAR                       54.844 LAYER ME2 ;
 ANTENNAMAXAREACAR                       65.956 LAYER ME3 ;
 ANTENNAMAXAREACAR                       77.067 LAYER ME4 ;
END WEB14
PIN DI112
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 2360.000 0.000 2360.800 1.000 ;
  LAYER ME3 ;
  RECT 2360.000 0.000 2360.800 1.000 ;
  LAYER ME2 ;
  RECT 2360.000 0.000 2360.800 1.000 ;
  LAYER ME1 ;
  RECT 2360.000 0.000 2360.800 1.000 ;
 END
 ANTENNAPARTIALMETALAREA                  3.130 LAYER ME2 ;
 ANTENNAGATEAREA                          0.086 LAYER ME2 ;
 ANTENNAGATEAREA                          0.086 LAYER ME3 ;
 ANTENNAGATEAREA                          0.086 LAYER ME4 ;
 ANTENNADIFFAREA                          0.160 LAYER ME2 ;
 ANTENNADIFFAREA                          0.160 LAYER ME3 ;
 ANTENNADIFFAREA                          0.160 LAYER ME4 ;
 ANTENNAMAXAREACAR                       48.569 LAYER ME2 ;
 ANTENNAMAXAREACAR                       57.829 LAYER ME3 ;
 ANTENNAMAXAREACAR                       67.088 LAYER ME4 ;
END DI112
PIN DO111
  DIRECTION OUTPUT ;
 PORT
  LAYER ME4 ;
  RECT 2353.600 0.000 2354.400 1.000 ;
  LAYER ME3 ;
  RECT 2353.600 0.000 2354.400 1.000 ;
  LAYER ME2 ;
  RECT 2353.600 0.000 2354.400 1.000 ;
  LAYER ME1 ;
  RECT 2353.600 0.000 2354.400 1.000 ;
 END
 ANTENNAPARTIALMETALAREA                  4.144 LAYER ME2 ;
 ANTENNADIFFAREA                          5.472 LAYER ME2 ;
 ANTENNADIFFAREA                          5.472 LAYER ME3 ;
 ANTENNADIFFAREA                          5.472 LAYER ME4 ;
END DO111
PIN DI111
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 2338.800 0.000 2339.600 1.000 ;
  LAYER ME3 ;
  RECT 2338.800 0.000 2339.600 1.000 ;
  LAYER ME2 ;
  RECT 2338.800 0.000 2339.600 1.000 ;
  LAYER ME1 ;
  RECT 2338.800 0.000 2339.600 1.000 ;
 END
 ANTENNAPARTIALMETALAREA                  3.154 LAYER ME2 ;
 ANTENNAGATEAREA                          0.086 LAYER ME2 ;
 ANTENNAGATEAREA                          0.086 LAYER ME3 ;
 ANTENNAGATEAREA                          0.086 LAYER ME4 ;
 ANTENNADIFFAREA                          0.160 LAYER ME2 ;
 ANTENNADIFFAREA                          0.160 LAYER ME3 ;
 ANTENNADIFFAREA                          0.160 LAYER ME4 ;
 ANTENNAMAXAREACAR                       48.847 LAYER ME2 ;
 ANTENNAMAXAREACAR                       58.106 LAYER ME3 ;
 ANTENNAMAXAREACAR                       67.366 LAYER ME4 ;
END DI111
PIN DO110
  DIRECTION OUTPUT ;
 PORT
  LAYER ME4 ;
  RECT 2333.600 0.000 2334.400 1.000 ;
  LAYER ME3 ;
  RECT 2333.600 0.000 2334.400 1.000 ;
  LAYER ME2 ;
  RECT 2333.600 0.000 2334.400 1.000 ;
  LAYER ME1 ;
  RECT 2333.600 0.000 2334.400 1.000 ;
 END
 ANTENNAPARTIALMETALAREA                  4.176 LAYER ME2 ;
 ANTENNADIFFAREA                          5.472 LAYER ME2 ;
 ANTENNADIFFAREA                          5.472 LAYER ME3 ;
 ANTENNADIFFAREA                          5.472 LAYER ME4 ;
END DO110
PIN DI110
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 2319.200 0.000 2320.000 1.000 ;
  LAYER ME3 ;
  RECT 2319.200 0.000 2320.000 1.000 ;
  LAYER ME2 ;
  RECT 2319.200 0.000 2320.000 1.000 ;
  LAYER ME1 ;
  RECT 2319.200 0.000 2320.000 1.000 ;
 END
 ANTENNAPARTIALMETALAREA                  3.126 LAYER ME2 ;
 ANTENNAGATEAREA                          0.086 LAYER ME2 ;
 ANTENNAGATEAREA                          0.086 LAYER ME3 ;
 ANTENNAGATEAREA                          0.086 LAYER ME4 ;
 ANTENNADIFFAREA                          0.160 LAYER ME2 ;
 ANTENNADIFFAREA                          0.160 LAYER ME3 ;
 ANTENNADIFFAREA                          0.160 LAYER ME4 ;
 ANTENNAMAXAREACAR                       48.523 LAYER ME2 ;
 ANTENNAMAXAREACAR                       57.782 LAYER ME3 ;
 ANTENNAMAXAREACAR                       67.042 LAYER ME4 ;
END DI110
PIN DO109
  DIRECTION OUTPUT ;
 PORT
  LAYER ME4 ;
  RECT 2312.800 0.000 2313.600 1.000 ;
  LAYER ME3 ;
  RECT 2312.800 0.000 2313.600 1.000 ;
  LAYER ME2 ;
  RECT 2312.800 0.000 2313.600 1.000 ;
  LAYER ME1 ;
  RECT 2312.800 0.000 2313.600 1.000 ;
 END
 ANTENNAPARTIALMETALAREA                  4.160 LAYER ME2 ;
 ANTENNADIFFAREA                          5.472 LAYER ME2 ;
 ANTENNADIFFAREA                          5.472 LAYER ME3 ;
 ANTENNADIFFAREA                          5.472 LAYER ME4 ;
END DO109
PIN DI109
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 2298.000 0.000 2298.800 1.000 ;
  LAYER ME3 ;
  RECT 2298.000 0.000 2298.800 1.000 ;
  LAYER ME2 ;
  RECT 2298.000 0.000 2298.800 1.000 ;
  LAYER ME1 ;
  RECT 2298.000 0.000 2298.800 1.000 ;
 END
 ANTENNAPARTIALMETALAREA                  3.130 LAYER ME2 ;
 ANTENNAGATEAREA                          0.086 LAYER ME2 ;
 ANTENNAGATEAREA                          0.086 LAYER ME3 ;
 ANTENNAGATEAREA                          0.086 LAYER ME4 ;
 ANTENNADIFFAREA                          0.160 LAYER ME2 ;
 ANTENNADIFFAREA                          0.160 LAYER ME3 ;
 ANTENNADIFFAREA                          0.160 LAYER ME4 ;
 ANTENNAMAXAREACAR                       48.569 LAYER ME2 ;
 ANTENNAMAXAREACAR                       57.829 LAYER ME3 ;
 ANTENNAMAXAREACAR                       67.088 LAYER ME4 ;
END DI109
PIN DO108
  DIRECTION OUTPUT ;
 PORT
  LAYER ME4 ;
  RECT 2292.800 0.000 2293.600 1.000 ;
  LAYER ME3 ;
  RECT 2292.800 0.000 2293.600 1.000 ;
  LAYER ME2 ;
  RECT 2292.800 0.000 2293.600 1.000 ;
  LAYER ME1 ;
  RECT 2292.800 0.000 2293.600 1.000 ;
 END
 ANTENNAPARTIALMETALAREA                  4.152 LAYER ME2 ;
 ANTENNADIFFAREA                          5.472 LAYER ME2 ;
 ANTENNADIFFAREA                          5.472 LAYER ME3 ;
 ANTENNADIFFAREA                          5.472 LAYER ME4 ;
END DO108
PIN DI108
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 2278.400 0.000 2279.200 1.000 ;
  LAYER ME3 ;
  RECT 2278.400 0.000 2279.200 1.000 ;
  LAYER ME2 ;
  RECT 2278.400 0.000 2279.200 1.000 ;
  LAYER ME1 ;
  RECT 2278.400 0.000 2279.200 1.000 ;
 END
 ANTENNAPARTIALMETALAREA                  3.150 LAYER ME2 ;
 ANTENNAGATEAREA                          0.086 LAYER ME2 ;
 ANTENNAGATEAREA                          0.086 LAYER ME3 ;
 ANTENNAGATEAREA                          0.086 LAYER ME4 ;
 ANTENNADIFFAREA                          0.160 LAYER ME2 ;
 ANTENNADIFFAREA                          0.160 LAYER ME3 ;
 ANTENNADIFFAREA                          0.160 LAYER ME4 ;
 ANTENNAMAXAREACAR                       48.801 LAYER ME2 ;
 ANTENNAMAXAREACAR                       58.060 LAYER ME3 ;
 ANTENNAMAXAREACAR                       67.319 LAYER ME4 ;
END DI108
PIN DO107
  DIRECTION OUTPUT ;
 PORT
  LAYER ME4 ;
  RECT 2271.600 0.000 2272.400 1.000 ;
  LAYER ME3 ;
  RECT 2271.600 0.000 2272.400 1.000 ;
  LAYER ME2 ;
  RECT 2271.600 0.000 2272.400 1.000 ;
  LAYER ME1 ;
  RECT 2271.600 0.000 2272.400 1.000 ;
 END
 ANTENNAPARTIALMETALAREA                  4.176 LAYER ME2 ;
 ANTENNADIFFAREA                          5.472 LAYER ME2 ;
 ANTENNADIFFAREA                          5.472 LAYER ME3 ;
 ANTENNADIFFAREA                          5.472 LAYER ME4 ;
END DO107
PIN DI107
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 2257.200 0.000 2258.000 1.000 ;
  LAYER ME3 ;
  RECT 2257.200 0.000 2258.000 1.000 ;
  LAYER ME2 ;
  RECT 2257.200 0.000 2258.000 1.000 ;
  LAYER ME1 ;
  RECT 2257.200 0.000 2258.000 1.000 ;
 END
 ANTENNAPARTIALMETALAREA                  3.126 LAYER ME2 ;
 ANTENNAGATEAREA                          0.086 LAYER ME2 ;
 ANTENNAGATEAREA                          0.086 LAYER ME3 ;
 ANTENNAGATEAREA                          0.086 LAYER ME4 ;
 ANTENNADIFFAREA                          0.160 LAYER ME2 ;
 ANTENNADIFFAREA                          0.160 LAYER ME3 ;
 ANTENNADIFFAREA                          0.160 LAYER ME4 ;
 ANTENNAMAXAREACAR                       48.523 LAYER ME2 ;
 ANTENNAMAXAREACAR                       57.782 LAYER ME3 ;
 ANTENNAMAXAREACAR                       67.042 LAYER ME4 ;
END DI107
PIN DO106
  DIRECTION OUTPUT ;
 PORT
  LAYER ME4 ;
  RECT 2252.000 0.000 2252.800 1.000 ;
  LAYER ME3 ;
  RECT 2252.000 0.000 2252.800 1.000 ;
  LAYER ME2 ;
  RECT 2252.000 0.000 2252.800 1.000 ;
  LAYER ME1 ;
  RECT 2252.000 0.000 2252.800 1.000 ;
 END
 ANTENNAPARTIALMETALAREA                  4.152 LAYER ME2 ;
 ANTENNADIFFAREA                          5.472 LAYER ME2 ;
 ANTENNADIFFAREA                          5.472 LAYER ME3 ;
 ANTENNADIFFAREA                          5.472 LAYER ME4 ;
END DO106
PIN DI106
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 2237.200 0.000 2238.000 1.000 ;
  LAYER ME3 ;
  RECT 2237.200 0.000 2238.000 1.000 ;
  LAYER ME2 ;
  RECT 2237.200 0.000 2238.000 1.000 ;
  LAYER ME1 ;
  RECT 2237.200 0.000 2238.000 1.000 ;
 END
 ANTENNAPARTIALMETALAREA                  3.138 LAYER ME2 ;
 ANTENNAGATEAREA                          0.086 LAYER ME2 ;
 ANTENNAGATEAREA                          0.086 LAYER ME3 ;
 ANTENNAGATEAREA                          0.086 LAYER ME4 ;
 ANTENNADIFFAREA                          0.160 LAYER ME2 ;
 ANTENNADIFFAREA                          0.160 LAYER ME3 ;
 ANTENNADIFFAREA                          0.160 LAYER ME4 ;
 ANTENNAMAXAREACAR                       48.662 LAYER ME2 ;
 ANTENNAMAXAREACAR                       57.921 LAYER ME3 ;
 ANTENNAMAXAREACAR                       67.181 LAYER ME4 ;
END DI106
PIN DO105
  DIRECTION OUTPUT ;
 PORT
  LAYER ME4 ;
  RECT 2230.800 0.000 2231.600 1.000 ;
  LAYER ME3 ;
  RECT 2230.800 0.000 2231.600 1.000 ;
  LAYER ME2 ;
  RECT 2230.800 0.000 2231.600 1.000 ;
  LAYER ME1 ;
  RECT 2230.800 0.000 2231.600 1.000 ;
 END
 ANTENNAPARTIALMETALAREA                  4.152 LAYER ME2 ;
 ANTENNADIFFAREA                          5.472 LAYER ME2 ;
 ANTENNADIFFAREA                          5.472 LAYER ME3 ;
 ANTENNADIFFAREA                          5.472 LAYER ME4 ;
END DO105
PIN DI105
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 2216.400 0.000 2217.200 1.000 ;
  LAYER ME3 ;
  RECT 2216.400 0.000 2217.200 1.000 ;
  LAYER ME2 ;
  RECT 2216.400 0.000 2217.200 1.000 ;
  LAYER ME1 ;
  RECT 2216.400 0.000 2217.200 1.000 ;
 END
 ANTENNAPARTIALMETALAREA                  3.150 LAYER ME2 ;
 ANTENNAGATEAREA                          0.086 LAYER ME2 ;
 ANTENNAGATEAREA                          0.086 LAYER ME3 ;
 ANTENNAGATEAREA                          0.086 LAYER ME4 ;
 ANTENNADIFFAREA                          0.160 LAYER ME2 ;
 ANTENNADIFFAREA                          0.160 LAYER ME3 ;
 ANTENNADIFFAREA                          0.160 LAYER ME4 ;
 ANTENNAMAXAREACAR                       48.801 LAYER ME2 ;
 ANTENNAMAXAREACAR                       58.060 LAYER ME3 ;
 ANTENNAMAXAREACAR                       67.319 LAYER ME4 ;
END DI105
PIN DO104
  DIRECTION OUTPUT ;
 PORT
  LAYER ME4 ;
  RECT 2211.200 0.000 2212.000 1.000 ;
  LAYER ME3 ;
  RECT 2211.200 0.000 2212.000 1.000 ;
  LAYER ME2 ;
  RECT 2211.200 0.000 2212.000 1.000 ;
  LAYER ME1 ;
  RECT 2211.200 0.000 2212.000 1.000 ;
 END
 ANTENNAPARTIALMETALAREA                  4.176 LAYER ME2 ;
 ANTENNADIFFAREA                          5.472 LAYER ME2 ;
 ANTENNADIFFAREA                          5.472 LAYER ME3 ;
 ANTENNADIFFAREA                          5.472 LAYER ME4 ;
END DO104
PIN WEB13
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 2198.000 0.000 2198.800 1.000 ;
  LAYER ME3 ;
  RECT 2198.000 0.000 2198.800 1.000 ;
  LAYER ME2 ;
  RECT 2198.000 0.000 2198.800 1.000 ;
  LAYER ME1 ;
  RECT 2198.000 0.000 2198.800 1.000 ;
 END
 ANTENNAPARTIALMETALAREA                  2.852 LAYER ME2 ;
 ANTENNAGATEAREA                          0.072 LAYER ME2 ;
 ANTENNAGATEAREA                          0.072 LAYER ME3 ;
 ANTENNAGATEAREA                          0.072 LAYER ME4 ;
 ANTENNADIFFAREA                          0.160 LAYER ME2 ;
 ANTENNADIFFAREA                          0.160 LAYER ME3 ;
 ANTENNADIFFAREA                          0.160 LAYER ME4 ;
 ANTENNAMAXAREACAR                       54.622 LAYER ME2 ;
 ANTENNAMAXAREACAR                       65.733 LAYER ME3 ;
 ANTENNAMAXAREACAR                       76.844 LAYER ME4 ;
END WEB13
PIN DI104
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 2196.400 0.000 2197.200 1.000 ;
  LAYER ME3 ;
  RECT 2196.400 0.000 2197.200 1.000 ;
  LAYER ME2 ;
  RECT 2196.400 0.000 2197.200 1.000 ;
  LAYER ME1 ;
  RECT 2196.400 0.000 2197.200 1.000 ;
 END
 ANTENNAPARTIALMETALAREA                  3.118 LAYER ME2 ;
 ANTENNAGATEAREA                          0.086 LAYER ME2 ;
 ANTENNAGATEAREA                          0.086 LAYER ME3 ;
 ANTENNAGATEAREA                          0.086 LAYER ME4 ;
 ANTENNADIFFAREA                          0.160 LAYER ME2 ;
 ANTENNADIFFAREA                          0.160 LAYER ME3 ;
 ANTENNADIFFAREA                          0.160 LAYER ME4 ;
 ANTENNAMAXAREACAR                       48.431 LAYER ME2 ;
 ANTENNAMAXAREACAR                       57.690 LAYER ME3 ;
 ANTENNAMAXAREACAR                       66.949 LAYER ME4 ;
END DI104
PIN DO103
  DIRECTION OUTPUT ;
 PORT
  LAYER ME4 ;
  RECT 2190.000 0.000 2190.800 1.000 ;
  LAYER ME3 ;
  RECT 2190.000 0.000 2190.800 1.000 ;
  LAYER ME2 ;
  RECT 2190.000 0.000 2190.800 1.000 ;
  LAYER ME1 ;
  RECT 2190.000 0.000 2190.800 1.000 ;
 END
 ANTENNAPARTIALMETALAREA                  4.152 LAYER ME2 ;
 ANTENNADIFFAREA                          5.472 LAYER ME2 ;
 ANTENNADIFFAREA                          5.472 LAYER ME3 ;
 ANTENNADIFFAREA                          5.472 LAYER ME4 ;
END DO103
PIN DI103
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 2175.200 0.000 2176.000 1.000 ;
  LAYER ME3 ;
  RECT 2175.200 0.000 2176.000 1.000 ;
  LAYER ME2 ;
  RECT 2175.200 0.000 2176.000 1.000 ;
  LAYER ME1 ;
  RECT 2175.200 0.000 2176.000 1.000 ;
 END
 ANTENNAPARTIALMETALAREA                  3.138 LAYER ME2 ;
 ANTENNAGATEAREA                          0.086 LAYER ME2 ;
 ANTENNAGATEAREA                          0.086 LAYER ME3 ;
 ANTENNAGATEAREA                          0.086 LAYER ME4 ;
 ANTENNADIFFAREA                          0.160 LAYER ME2 ;
 ANTENNADIFFAREA                          0.160 LAYER ME3 ;
 ANTENNADIFFAREA                          0.160 LAYER ME4 ;
 ANTENNAMAXAREACAR                       48.662 LAYER ME2 ;
 ANTENNAMAXAREACAR                       57.921 LAYER ME3 ;
 ANTENNAMAXAREACAR                       67.181 LAYER ME4 ;
END DI103
PIN DO102
  DIRECTION OUTPUT ;
 PORT
  LAYER ME4 ;
  RECT 2170.000 0.000 2170.800 1.000 ;
  LAYER ME3 ;
  RECT 2170.000 0.000 2170.800 1.000 ;
  LAYER ME2 ;
  RECT 2170.000 0.000 2170.800 1.000 ;
  LAYER ME1 ;
  RECT 2170.000 0.000 2170.800 1.000 ;
 END
 ANTENNAPARTIALMETALAREA                  4.160 LAYER ME2 ;
 ANTENNADIFFAREA                          5.472 LAYER ME2 ;
 ANTENNADIFFAREA                          5.472 LAYER ME3 ;
 ANTENNADIFFAREA                          5.472 LAYER ME4 ;
END DO102
PIN DI102
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 2155.600 0.000 2156.400 1.000 ;
  LAYER ME3 ;
  RECT 2155.600 0.000 2156.400 1.000 ;
  LAYER ME2 ;
  RECT 2155.600 0.000 2156.400 1.000 ;
  LAYER ME1 ;
  RECT 2155.600 0.000 2156.400 1.000 ;
 END
 ANTENNAPARTIALMETALAREA                  3.142 LAYER ME2 ;
 ANTENNAGATEAREA                          0.086 LAYER ME2 ;
 ANTENNAGATEAREA                          0.086 LAYER ME3 ;
 ANTENNAGATEAREA                          0.086 LAYER ME4 ;
 ANTENNADIFFAREA                          0.160 LAYER ME2 ;
 ANTENNADIFFAREA                          0.160 LAYER ME3 ;
 ANTENNADIFFAREA                          0.160 LAYER ME4 ;
 ANTENNAMAXAREACAR                       48.708 LAYER ME2 ;
 ANTENNAMAXAREACAR                       57.968 LAYER ME3 ;
 ANTENNAMAXAREACAR                       67.227 LAYER ME4 ;
END DI102
PIN DO101
  DIRECTION OUTPUT ;
 PORT
  LAYER ME4 ;
  RECT 2149.200 0.000 2150.000 1.000 ;
  LAYER ME3 ;
  RECT 2149.200 0.000 2150.000 1.000 ;
  LAYER ME2 ;
  RECT 2149.200 0.000 2150.000 1.000 ;
  LAYER ME1 ;
  RECT 2149.200 0.000 2150.000 1.000 ;
 END
 ANTENNAPARTIALMETALAREA                  4.176 LAYER ME2 ;
 ANTENNADIFFAREA                          5.472 LAYER ME2 ;
 ANTENNADIFFAREA                          5.472 LAYER ME3 ;
 ANTENNADIFFAREA                          5.472 LAYER ME4 ;
END DO101
PIN DI101
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 2134.400 0.000 2135.200 1.000 ;
  LAYER ME3 ;
  RECT 2134.400 0.000 2135.200 1.000 ;
  LAYER ME2 ;
  RECT 2134.400 0.000 2135.200 1.000 ;
  LAYER ME1 ;
  RECT 2134.400 0.000 2135.200 1.000 ;
 END
 ANTENNAPARTIALMETALAREA                  3.118 LAYER ME2 ;
 ANTENNAGATEAREA                          0.086 LAYER ME2 ;
 ANTENNAGATEAREA                          0.086 LAYER ME3 ;
 ANTENNAGATEAREA                          0.086 LAYER ME4 ;
 ANTENNADIFFAREA                          0.160 LAYER ME2 ;
 ANTENNADIFFAREA                          0.160 LAYER ME3 ;
 ANTENNADIFFAREA                          0.160 LAYER ME4 ;
 ANTENNAMAXAREACAR                       48.431 LAYER ME2 ;
 ANTENNAMAXAREACAR                       57.690 LAYER ME3 ;
 ANTENNAMAXAREACAR                       66.949 LAYER ME4 ;
END DI101
PIN DO100
  DIRECTION OUTPUT ;
 PORT
  LAYER ME4 ;
  RECT 2129.200 0.000 2130.000 1.000 ;
  LAYER ME3 ;
  RECT 2129.200 0.000 2130.000 1.000 ;
  LAYER ME2 ;
  RECT 2129.200 0.000 2130.000 1.000 ;
  LAYER ME1 ;
  RECT 2129.200 0.000 2130.000 1.000 ;
 END
 ANTENNAPARTIALMETALAREA                  4.144 LAYER ME2 ;
 ANTENNADIFFAREA                          5.472 LAYER ME2 ;
 ANTENNADIFFAREA                          5.472 LAYER ME3 ;
 ANTENNADIFFAREA                          5.472 LAYER ME4 ;
END DO100
PIN DI100
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 2114.400 0.000 2115.200 1.000 ;
  LAYER ME3 ;
  RECT 2114.400 0.000 2115.200 1.000 ;
  LAYER ME2 ;
  RECT 2114.400 0.000 2115.200 1.000 ;
  LAYER ME1 ;
  RECT 2114.400 0.000 2115.200 1.000 ;
 END
 ANTENNAPARTIALMETALAREA                  3.146 LAYER ME2 ;
 ANTENNAGATEAREA                          0.086 LAYER ME2 ;
 ANTENNAGATEAREA                          0.086 LAYER ME3 ;
 ANTENNAGATEAREA                          0.086 LAYER ME4 ;
 ANTENNADIFFAREA                          0.160 LAYER ME2 ;
 ANTENNADIFFAREA                          0.160 LAYER ME3 ;
 ANTENNADIFFAREA                          0.160 LAYER ME4 ;
 ANTENNAMAXAREACAR                       48.755 LAYER ME2 ;
 ANTENNAMAXAREACAR                       58.014 LAYER ME3 ;
 ANTENNAMAXAREACAR                       67.273 LAYER ME4 ;
END DI100
PIN DO99
  DIRECTION OUTPUT ;
 PORT
  LAYER ME4 ;
  RECT 2108.000 0.000 2108.800 1.000 ;
  LAYER ME3 ;
  RECT 2108.000 0.000 2108.800 1.000 ;
  LAYER ME2 ;
  RECT 2108.000 0.000 2108.800 1.000 ;
  LAYER ME1 ;
  RECT 2108.000 0.000 2108.800 1.000 ;
 END
 ANTENNAPARTIALMETALAREA                  4.160 LAYER ME2 ;
 ANTENNADIFFAREA                          5.472 LAYER ME2 ;
 ANTENNADIFFAREA                          5.472 LAYER ME3 ;
 ANTENNADIFFAREA                          5.472 LAYER ME4 ;
END DO99
PIN DI99
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 2093.600 0.000 2094.400 1.000 ;
  LAYER ME3 ;
  RECT 2093.600 0.000 2094.400 1.000 ;
  LAYER ME2 ;
  RECT 2093.600 0.000 2094.400 1.000 ;
  LAYER ME1 ;
  RECT 2093.600 0.000 2094.400 1.000 ;
 END
 ANTENNAPARTIALMETALAREA                  3.142 LAYER ME2 ;
 ANTENNAGATEAREA                          0.086 LAYER ME2 ;
 ANTENNAGATEAREA                          0.086 LAYER ME3 ;
 ANTENNAGATEAREA                          0.086 LAYER ME4 ;
 ANTENNADIFFAREA                          0.160 LAYER ME2 ;
 ANTENNADIFFAREA                          0.160 LAYER ME3 ;
 ANTENNADIFFAREA                          0.160 LAYER ME4 ;
 ANTENNAMAXAREACAR                       48.708 LAYER ME2 ;
 ANTENNAMAXAREACAR                       57.968 LAYER ME3 ;
 ANTENNAMAXAREACAR                       67.227 LAYER ME4 ;
END DI99
PIN DO98
  DIRECTION OUTPUT ;
 PORT
  LAYER ME4 ;
  RECT 2088.400 0.000 2089.200 1.000 ;
  LAYER ME3 ;
  RECT 2088.400 0.000 2089.200 1.000 ;
  LAYER ME2 ;
  RECT 2088.400 0.000 2089.200 1.000 ;
  LAYER ME1 ;
  RECT 2088.400 0.000 2089.200 1.000 ;
 END
 ANTENNAPARTIALMETALAREA                  4.168 LAYER ME2 ;
 ANTENNADIFFAREA                          5.472 LAYER ME2 ;
 ANTENNADIFFAREA                          5.472 LAYER ME3 ;
 ANTENNADIFFAREA                          5.472 LAYER ME4 ;
END DO98
PIN DI98
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 2073.600 0.000 2074.400 1.000 ;
  LAYER ME3 ;
  RECT 2073.600 0.000 2074.400 1.000 ;
  LAYER ME2 ;
  RECT 2073.600 0.000 2074.400 1.000 ;
  LAYER ME1 ;
  RECT 2073.600 0.000 2074.400 1.000 ;
 END
 ANTENNAPARTIALMETALAREA                  3.122 LAYER ME2 ;
 ANTENNAGATEAREA                          0.086 LAYER ME2 ;
 ANTENNAGATEAREA                          0.086 LAYER ME3 ;
 ANTENNAGATEAREA                          0.086 LAYER ME4 ;
 ANTENNADIFFAREA                          0.160 LAYER ME2 ;
 ANTENNADIFFAREA                          0.160 LAYER ME3 ;
 ANTENNADIFFAREA                          0.160 LAYER ME4 ;
 ANTENNAMAXAREACAR                       48.477 LAYER ME2 ;
 ANTENNAMAXAREACAR                       57.736 LAYER ME3 ;
 ANTENNAMAXAREACAR                       66.995 LAYER ME4 ;
END DI98
PIN DO97
  DIRECTION OUTPUT ;
 PORT
  LAYER ME4 ;
  RECT 2067.200 0.000 2068.000 1.000 ;
  LAYER ME3 ;
  RECT 2067.200 0.000 2068.000 1.000 ;
  LAYER ME2 ;
  RECT 2067.200 0.000 2068.000 1.000 ;
  LAYER ME1 ;
  RECT 2067.200 0.000 2068.000 1.000 ;
 END
 ANTENNAPARTIALMETALAREA                  4.144 LAYER ME2 ;
 ANTENNADIFFAREA                          5.472 LAYER ME2 ;
 ANTENNADIFFAREA                          5.472 LAYER ME3 ;
 ANTENNADIFFAREA                          5.472 LAYER ME4 ;
END DO97
PIN DI97
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 2052.400 0.000 2053.200 1.000 ;
  LAYER ME3 ;
  RECT 2052.400 0.000 2053.200 1.000 ;
  LAYER ME2 ;
  RECT 2052.400 0.000 2053.200 1.000 ;
  LAYER ME1 ;
  RECT 2052.400 0.000 2053.200 1.000 ;
 END
 ANTENNAPARTIALMETALAREA                  3.146 LAYER ME2 ;
 ANTENNAGATEAREA                          0.086 LAYER ME2 ;
 ANTENNAGATEAREA                          0.086 LAYER ME3 ;
 ANTENNAGATEAREA                          0.086 LAYER ME4 ;
 ANTENNADIFFAREA                          0.160 LAYER ME2 ;
 ANTENNADIFFAREA                          0.160 LAYER ME3 ;
 ANTENNADIFFAREA                          0.160 LAYER ME4 ;
 ANTENNAMAXAREACAR                       48.755 LAYER ME2 ;
 ANTENNAMAXAREACAR                       58.014 LAYER ME3 ;
 ANTENNAMAXAREACAR                       67.273 LAYER ME4 ;
END DI97
PIN DO96
  DIRECTION OUTPUT ;
 PORT
  LAYER ME4 ;
  RECT 2047.200 0.000 2048.000 1.000 ;
  LAYER ME3 ;
  RECT 2047.200 0.000 2048.000 1.000 ;
  LAYER ME2 ;
  RECT 2047.200 0.000 2048.000 1.000 ;
  LAYER ME1 ;
  RECT 2047.200 0.000 2048.000 1.000 ;
 END
 ANTENNAPARTIALMETALAREA                  4.168 LAYER ME2 ;
 ANTENNADIFFAREA                          5.472 LAYER ME2 ;
 ANTENNADIFFAREA                          5.472 LAYER ME3 ;
 ANTENNADIFFAREA                          5.472 LAYER ME4 ;
END DO96
PIN WEB12
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 2034.400 0.000 2035.200 1.000 ;
  LAYER ME3 ;
  RECT 2034.400 0.000 2035.200 1.000 ;
  LAYER ME2 ;
  RECT 2034.400 0.000 2035.200 1.000 ;
  LAYER ME1 ;
  RECT 2034.400 0.000 2035.200 1.000 ;
 END
 ANTENNAPARTIALMETALAREA                  2.836 LAYER ME2 ;
 ANTENNAGATEAREA                          0.072 LAYER ME2 ;
 ANTENNAGATEAREA                          0.072 LAYER ME3 ;
 ANTENNAGATEAREA                          0.072 LAYER ME4 ;
 ANTENNADIFFAREA                          0.160 LAYER ME2 ;
 ANTENNADIFFAREA                          0.160 LAYER ME3 ;
 ANTENNADIFFAREA                          0.160 LAYER ME4 ;
 ANTENNAMAXAREACAR                       54.400 LAYER ME2 ;
 ANTENNAMAXAREACAR                       65.511 LAYER ME3 ;
 ANTENNAMAXAREACAR                       76.622 LAYER ME4 ;
END WEB12
PIN DI96
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 2032.800 0.000 2033.600 1.000 ;
  LAYER ME3 ;
  RECT 2032.800 0.000 2033.600 1.000 ;
  LAYER ME2 ;
  RECT 2032.800 0.000 2033.600 1.000 ;
  LAYER ME1 ;
  RECT 2032.800 0.000 2033.600 1.000 ;
 END
 ANTENNAPARTIALMETALAREA                  3.134 LAYER ME2 ;
 ANTENNAGATEAREA                          0.086 LAYER ME2 ;
 ANTENNAGATEAREA                          0.086 LAYER ME3 ;
 ANTENNAGATEAREA                          0.086 LAYER ME4 ;
 ANTENNADIFFAREA                          0.160 LAYER ME2 ;
 ANTENNADIFFAREA                          0.160 LAYER ME3 ;
 ANTENNADIFFAREA                          0.160 LAYER ME4 ;
 ANTENNAMAXAREACAR                       48.616 LAYER ME2 ;
 ANTENNAMAXAREACAR                       57.875 LAYER ME3 ;
 ANTENNAMAXAREACAR                       67.134 LAYER ME4 ;
END DI96
PIN DO95
  DIRECTION OUTPUT ;
 PORT
  LAYER ME4 ;
  RECT 2026.400 0.000 2027.200 1.000 ;
  LAYER ME3 ;
  RECT 2026.400 0.000 2027.200 1.000 ;
  LAYER ME2 ;
  RECT 2026.400 0.000 2027.200 1.000 ;
  LAYER ME1 ;
  RECT 2026.400 0.000 2027.200 1.000 ;
 END
 ANTENNAPARTIALMETALAREA                  4.168 LAYER ME2 ;
 ANTENNADIFFAREA                          5.472 LAYER ME2 ;
 ANTENNADIFFAREA                          5.472 LAYER ME3 ;
 ANTENNADIFFAREA                          5.472 LAYER ME4 ;
END DO95
PIN DI95
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 2011.600 0.000 2012.400 1.000 ;
  LAYER ME3 ;
  RECT 2011.600 0.000 2012.400 1.000 ;
  LAYER ME2 ;
  RECT 2011.600 0.000 2012.400 1.000 ;
  LAYER ME1 ;
  RECT 2011.600 0.000 2012.400 1.000 ;
 END
 ANTENNAPARTIALMETALAREA                  3.122 LAYER ME2 ;
 ANTENNAGATEAREA                          0.086 LAYER ME2 ;
 ANTENNAGATEAREA                          0.086 LAYER ME3 ;
 ANTENNAGATEAREA                          0.086 LAYER ME4 ;
 ANTENNADIFFAREA                          0.160 LAYER ME2 ;
 ANTENNADIFFAREA                          0.160 LAYER ME3 ;
 ANTENNADIFFAREA                          0.160 LAYER ME4 ;
 ANTENNAMAXAREACAR                       48.477 LAYER ME2 ;
 ANTENNAMAXAREACAR                       57.736 LAYER ME3 ;
 ANTENNAMAXAREACAR                       66.995 LAYER ME4 ;
END DI95
PIN DO94
  DIRECTION OUTPUT ;
 PORT
  LAYER ME4 ;
  RECT 2006.400 0.000 2007.200 1.000 ;
  LAYER ME3 ;
  RECT 2006.400 0.000 2007.200 1.000 ;
  LAYER ME2 ;
  RECT 2006.400 0.000 2007.200 1.000 ;
  LAYER ME1 ;
  RECT 2006.400 0.000 2007.200 1.000 ;
 END
 ANTENNAPARTIALMETALAREA                  4.144 LAYER ME2 ;
 ANTENNADIFFAREA                          5.472 LAYER ME2 ;
 ANTENNADIFFAREA                          5.472 LAYER ME3 ;
 ANTENNADIFFAREA                          5.472 LAYER ME4 ;
END DO94
PIN DI94
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 1991.600 0.000 1992.400 1.000 ;
  LAYER ME3 ;
  RECT 1991.600 0.000 1992.400 1.000 ;
  LAYER ME2 ;
  RECT 1991.600 0.000 1992.400 1.000 ;
  LAYER ME1 ;
  RECT 1991.600 0.000 1992.400 1.000 ;
 END
 ANTENNAPARTIALMETALAREA                  3.154 LAYER ME2 ;
 ANTENNAGATEAREA                          0.086 LAYER ME2 ;
 ANTENNAGATEAREA                          0.086 LAYER ME3 ;
 ANTENNAGATEAREA                          0.086 LAYER ME4 ;
 ANTENNADIFFAREA                          0.160 LAYER ME2 ;
 ANTENNADIFFAREA                          0.160 LAYER ME3 ;
 ANTENNADIFFAREA                          0.160 LAYER ME4 ;
 ANTENNAMAXAREACAR                       48.847 LAYER ME2 ;
 ANTENNAMAXAREACAR                       58.106 LAYER ME3 ;
 ANTENNAMAXAREACAR                       67.366 LAYER ME4 ;
END DI94
PIN DO93
  DIRECTION OUTPUT ;
 PORT
  LAYER ME4 ;
  RECT 1985.200 0.000 1986.000 1.000 ;
  LAYER ME3 ;
  RECT 1985.200 0.000 1986.000 1.000 ;
  LAYER ME2 ;
  RECT 1985.200 0.000 1986.000 1.000 ;
  LAYER ME1 ;
  RECT 1985.200 0.000 1986.000 1.000 ;
 END
 ANTENNAPARTIALMETALAREA                  4.168 LAYER ME2 ;
 ANTENNADIFFAREA                          5.472 LAYER ME2 ;
 ANTENNADIFFAREA                          5.472 LAYER ME3 ;
 ANTENNADIFFAREA                          5.472 LAYER ME4 ;
END DO93
PIN DI93
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 1970.800 0.000 1971.600 1.000 ;
  LAYER ME3 ;
  RECT 1970.800 0.000 1971.600 1.000 ;
  LAYER ME2 ;
  RECT 1970.800 0.000 1971.600 1.000 ;
  LAYER ME1 ;
  RECT 1970.800 0.000 1971.600 1.000 ;
 END
 ANTENNAPARTIALMETALAREA                  3.134 LAYER ME2 ;
 ANTENNAGATEAREA                          0.086 LAYER ME2 ;
 ANTENNAGATEAREA                          0.086 LAYER ME3 ;
 ANTENNAGATEAREA                          0.086 LAYER ME4 ;
 ANTENNADIFFAREA                          0.160 LAYER ME2 ;
 ANTENNADIFFAREA                          0.160 LAYER ME3 ;
 ANTENNADIFFAREA                          0.160 LAYER ME4 ;
 ANTENNAMAXAREACAR                       48.616 LAYER ME2 ;
 ANTENNAMAXAREACAR                       57.875 LAYER ME3 ;
 ANTENNAMAXAREACAR                       67.134 LAYER ME4 ;
END DI93
PIN DO92
  DIRECTION OUTPUT ;
 PORT
  LAYER ME4 ;
  RECT 1965.600 0.000 1966.400 1.000 ;
  LAYER ME3 ;
  RECT 1965.600 0.000 1966.400 1.000 ;
  LAYER ME2 ;
  RECT 1965.600 0.000 1966.400 1.000 ;
  LAYER ME1 ;
  RECT 1965.600 0.000 1966.400 1.000 ;
 END
 ANTENNAPARTIALMETALAREA                  4.160 LAYER ME2 ;
 ANTENNADIFFAREA                          5.472 LAYER ME2 ;
 ANTENNADIFFAREA                          5.472 LAYER ME3 ;
 ANTENNADIFFAREA                          5.472 LAYER ME4 ;
END DO92
PIN DI92
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 1950.800 0.000 1951.600 1.000 ;
  LAYER ME3 ;
  RECT 1950.800 0.000 1951.600 1.000 ;
  LAYER ME2 ;
  RECT 1950.800 0.000 1951.600 1.000 ;
  LAYER ME1 ;
  RECT 1950.800 0.000 1951.600 1.000 ;
 END
 ANTENNAPARTIALMETALAREA                  3.130 LAYER ME2 ;
 ANTENNAGATEAREA                          0.086 LAYER ME2 ;
 ANTENNAGATEAREA                          0.086 LAYER ME3 ;
 ANTENNAGATEAREA                          0.086 LAYER ME4 ;
 ANTENNADIFFAREA                          0.160 LAYER ME2 ;
 ANTENNADIFFAREA                          0.160 LAYER ME3 ;
 ANTENNADIFFAREA                          0.160 LAYER ME4 ;
 ANTENNAMAXAREACAR                       48.569 LAYER ME2 ;
 ANTENNAMAXAREACAR                       57.829 LAYER ME3 ;
 ANTENNAMAXAREACAR                       67.088 LAYER ME4 ;
END DI92
PIN DO91
  DIRECTION OUTPUT ;
 PORT
  LAYER ME4 ;
  RECT 1944.400 0.000 1945.200 1.000 ;
  LAYER ME3 ;
  RECT 1944.400 0.000 1945.200 1.000 ;
  LAYER ME2 ;
  RECT 1944.400 0.000 1945.200 1.000 ;
  LAYER ME1 ;
  RECT 1944.400 0.000 1945.200 1.000 ;
 END
 ANTENNAPARTIALMETALAREA                  4.144 LAYER ME2 ;
 ANTENNADIFFAREA                          5.472 LAYER ME2 ;
 ANTENNADIFFAREA                          5.472 LAYER ME3 ;
 ANTENNADIFFAREA                          5.472 LAYER ME4 ;
END DO91
PIN DI91
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 1929.600 0.000 1930.400 1.000 ;
  LAYER ME3 ;
  RECT 1929.600 0.000 1930.400 1.000 ;
  LAYER ME2 ;
  RECT 1929.600 0.000 1930.400 1.000 ;
  LAYER ME1 ;
  RECT 1929.600 0.000 1930.400 1.000 ;
 END
 ANTENNAPARTIALMETALAREA                  3.154 LAYER ME2 ;
 ANTENNAGATEAREA                          0.086 LAYER ME2 ;
 ANTENNAGATEAREA                          0.086 LAYER ME3 ;
 ANTENNAGATEAREA                          0.086 LAYER ME4 ;
 ANTENNADIFFAREA                          0.160 LAYER ME2 ;
 ANTENNADIFFAREA                          0.160 LAYER ME3 ;
 ANTENNADIFFAREA                          0.160 LAYER ME4 ;
 ANTENNAMAXAREACAR                       48.847 LAYER ME2 ;
 ANTENNAMAXAREACAR                       58.106 LAYER ME3 ;
 ANTENNAMAXAREACAR                       67.366 LAYER ME4 ;
END DI91
PIN DO90
  DIRECTION OUTPUT ;
 PORT
  LAYER ME4 ;
  RECT 1924.400 0.000 1925.200 1.000 ;
  LAYER ME3 ;
  RECT 1924.400 0.000 1925.200 1.000 ;
  LAYER ME2 ;
  RECT 1924.400 0.000 1925.200 1.000 ;
  LAYER ME1 ;
  RECT 1924.400 0.000 1925.200 1.000 ;
 END
 ANTENNAPARTIALMETALAREA                  4.176 LAYER ME2 ;
 ANTENNADIFFAREA                          5.472 LAYER ME2 ;
 ANTENNADIFFAREA                          5.472 LAYER ME3 ;
 ANTENNADIFFAREA                          5.472 LAYER ME4 ;
END DO90
PIN DI90
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 1910.000 0.000 1910.800 1.000 ;
  LAYER ME3 ;
  RECT 1910.000 0.000 1910.800 1.000 ;
  LAYER ME2 ;
  RECT 1910.000 0.000 1910.800 1.000 ;
  LAYER ME1 ;
  RECT 1910.000 0.000 1910.800 1.000 ;
 END
 ANTENNAPARTIALMETALAREA                  3.126 LAYER ME2 ;
 ANTENNAGATEAREA                          0.086 LAYER ME2 ;
 ANTENNAGATEAREA                          0.086 LAYER ME3 ;
 ANTENNAGATEAREA                          0.086 LAYER ME4 ;
 ANTENNADIFFAREA                          0.160 LAYER ME2 ;
 ANTENNADIFFAREA                          0.160 LAYER ME3 ;
 ANTENNADIFFAREA                          0.160 LAYER ME4 ;
 ANTENNAMAXAREACAR                       48.523 LAYER ME2 ;
 ANTENNAMAXAREACAR                       57.782 LAYER ME3 ;
 ANTENNAMAXAREACAR                       67.042 LAYER ME4 ;
END DI90
PIN DO89
  DIRECTION OUTPUT ;
 PORT
  LAYER ME4 ;
  RECT 1903.600 0.000 1904.400 1.000 ;
  LAYER ME3 ;
  RECT 1903.600 0.000 1904.400 1.000 ;
  LAYER ME2 ;
  RECT 1903.600 0.000 1904.400 1.000 ;
  LAYER ME1 ;
  RECT 1903.600 0.000 1904.400 1.000 ;
 END
 ANTENNAPARTIALMETALAREA                  4.160 LAYER ME2 ;
 ANTENNADIFFAREA                          5.472 LAYER ME2 ;
 ANTENNADIFFAREA                          5.472 LAYER ME3 ;
 ANTENNADIFFAREA                          5.472 LAYER ME4 ;
END DO89
PIN DI89
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 1888.800 0.000 1889.600 1.000 ;
  LAYER ME3 ;
  RECT 1888.800 0.000 1889.600 1.000 ;
  LAYER ME2 ;
  RECT 1888.800 0.000 1889.600 1.000 ;
  LAYER ME1 ;
  RECT 1888.800 0.000 1889.600 1.000 ;
 END
 ANTENNAPARTIALMETALAREA                  3.130 LAYER ME2 ;
 ANTENNAGATEAREA                          0.086 LAYER ME2 ;
 ANTENNAGATEAREA                          0.086 LAYER ME3 ;
 ANTENNAGATEAREA                          0.086 LAYER ME4 ;
 ANTENNADIFFAREA                          0.160 LAYER ME2 ;
 ANTENNADIFFAREA                          0.160 LAYER ME3 ;
 ANTENNADIFFAREA                          0.160 LAYER ME4 ;
 ANTENNAMAXAREACAR                       48.569 LAYER ME2 ;
 ANTENNAMAXAREACAR                       57.829 LAYER ME3 ;
 ANTENNAMAXAREACAR                       67.088 LAYER ME4 ;
END DI89
PIN DO88
  DIRECTION OUTPUT ;
 PORT
  LAYER ME4 ;
  RECT 1883.600 0.000 1884.400 1.000 ;
  LAYER ME3 ;
  RECT 1883.600 0.000 1884.400 1.000 ;
  LAYER ME2 ;
  RECT 1883.600 0.000 1884.400 1.000 ;
  LAYER ME1 ;
  RECT 1883.600 0.000 1884.400 1.000 ;
 END
 ANTENNAPARTIALMETALAREA                  4.152 LAYER ME2 ;
 ANTENNADIFFAREA                          5.472 LAYER ME2 ;
 ANTENNADIFFAREA                          5.472 LAYER ME3 ;
 ANTENNADIFFAREA                          5.472 LAYER ME4 ;
END DO88
PIN WEB11
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 1870.800 0.000 1871.600 1.000 ;
  LAYER ME3 ;
  RECT 1870.800 0.000 1871.600 1.000 ;
  LAYER ME2 ;
  RECT 1870.800 0.000 1871.600 1.000 ;
  LAYER ME1 ;
  RECT 1870.800 0.000 1871.600 1.000 ;
 END
 ANTENNAPARTIALMETALAREA                  2.840 LAYER ME2 ;
 ANTENNAGATEAREA                          0.072 LAYER ME2 ;
 ANTENNAGATEAREA                          0.072 LAYER ME3 ;
 ANTENNAGATEAREA                          0.072 LAYER ME4 ;
 ANTENNADIFFAREA                          0.160 LAYER ME2 ;
 ANTENNADIFFAREA                          0.160 LAYER ME3 ;
 ANTENNADIFFAREA                          0.160 LAYER ME4 ;
 ANTENNAMAXAREACAR                       54.456 LAYER ME2 ;
 ANTENNAMAXAREACAR                       65.567 LAYER ME3 ;
 ANTENNAMAXAREACAR                       76.678 LAYER ME4 ;
END WEB11
PIN DI88
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 1869.200 0.000 1870.000 1.000 ;
  LAYER ME3 ;
  RECT 1869.200 0.000 1870.000 1.000 ;
  LAYER ME2 ;
  RECT 1869.200 0.000 1870.000 1.000 ;
  LAYER ME1 ;
  RECT 1869.200 0.000 1870.000 1.000 ;
 END
 ANTENNAPARTIALMETALAREA                  3.150 LAYER ME2 ;
 ANTENNAGATEAREA                          0.086 LAYER ME2 ;
 ANTENNAGATEAREA                          0.086 LAYER ME3 ;
 ANTENNAGATEAREA                          0.086 LAYER ME4 ;
 ANTENNADIFFAREA                          0.160 LAYER ME2 ;
 ANTENNADIFFAREA                          0.160 LAYER ME3 ;
 ANTENNADIFFAREA                          0.160 LAYER ME4 ;
 ANTENNAMAXAREACAR                       48.801 LAYER ME2 ;
 ANTENNAMAXAREACAR                       58.060 LAYER ME3 ;
 ANTENNAMAXAREACAR                       67.319 LAYER ME4 ;
END DI88
PIN DO87
  DIRECTION OUTPUT ;
 PORT
  LAYER ME4 ;
  RECT 1862.400 0.000 1863.200 1.000 ;
  LAYER ME3 ;
  RECT 1862.400 0.000 1863.200 1.000 ;
  LAYER ME2 ;
  RECT 1862.400 0.000 1863.200 1.000 ;
  LAYER ME1 ;
  RECT 1862.400 0.000 1863.200 1.000 ;
 END
 ANTENNAPARTIALMETALAREA                  4.176 LAYER ME2 ;
 ANTENNADIFFAREA                          5.472 LAYER ME2 ;
 ANTENNADIFFAREA                          5.472 LAYER ME3 ;
 ANTENNADIFFAREA                          5.472 LAYER ME4 ;
END DO87
PIN DI87
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 1848.000 0.000 1848.800 1.000 ;
  LAYER ME3 ;
  RECT 1848.000 0.000 1848.800 1.000 ;
  LAYER ME2 ;
  RECT 1848.000 0.000 1848.800 1.000 ;
  LAYER ME1 ;
  RECT 1848.000 0.000 1848.800 1.000 ;
 END
 ANTENNAPARTIALMETALAREA                  3.126 LAYER ME2 ;
 ANTENNAGATEAREA                          0.086 LAYER ME2 ;
 ANTENNAGATEAREA                          0.086 LAYER ME3 ;
 ANTENNAGATEAREA                          0.086 LAYER ME4 ;
 ANTENNADIFFAREA                          0.160 LAYER ME2 ;
 ANTENNADIFFAREA                          0.160 LAYER ME3 ;
 ANTENNADIFFAREA                          0.160 LAYER ME4 ;
 ANTENNAMAXAREACAR                       48.523 LAYER ME2 ;
 ANTENNAMAXAREACAR                       57.782 LAYER ME3 ;
 ANTENNAMAXAREACAR                       67.042 LAYER ME4 ;
END DI87
PIN DO86
  DIRECTION OUTPUT ;
 PORT
  LAYER ME4 ;
  RECT 1842.800 0.000 1843.600 1.000 ;
  LAYER ME3 ;
  RECT 1842.800 0.000 1843.600 1.000 ;
  LAYER ME2 ;
  RECT 1842.800 0.000 1843.600 1.000 ;
  LAYER ME1 ;
  RECT 1842.800 0.000 1843.600 1.000 ;
 END
 ANTENNAPARTIALMETALAREA                  4.152 LAYER ME2 ;
 ANTENNADIFFAREA                          5.472 LAYER ME2 ;
 ANTENNADIFFAREA                          5.472 LAYER ME3 ;
 ANTENNADIFFAREA                          5.472 LAYER ME4 ;
END DO86
PIN DI86
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 1828.000 0.000 1828.800 1.000 ;
  LAYER ME3 ;
  RECT 1828.000 0.000 1828.800 1.000 ;
  LAYER ME2 ;
  RECT 1828.000 0.000 1828.800 1.000 ;
  LAYER ME1 ;
  RECT 1828.000 0.000 1828.800 1.000 ;
 END
 ANTENNAPARTIALMETALAREA                  3.138 LAYER ME2 ;
 ANTENNAGATEAREA                          0.086 LAYER ME2 ;
 ANTENNAGATEAREA                          0.086 LAYER ME3 ;
 ANTENNAGATEAREA                          0.086 LAYER ME4 ;
 ANTENNADIFFAREA                          0.160 LAYER ME2 ;
 ANTENNADIFFAREA                          0.160 LAYER ME3 ;
 ANTENNADIFFAREA                          0.160 LAYER ME4 ;
 ANTENNAMAXAREACAR                       48.662 LAYER ME2 ;
 ANTENNAMAXAREACAR                       57.921 LAYER ME3 ;
 ANTENNAMAXAREACAR                       67.181 LAYER ME4 ;
END DI86
PIN DO85
  DIRECTION OUTPUT ;
 PORT
  LAYER ME4 ;
  RECT 1821.600 0.000 1822.400 1.000 ;
  LAYER ME3 ;
  RECT 1821.600 0.000 1822.400 1.000 ;
  LAYER ME2 ;
  RECT 1821.600 0.000 1822.400 1.000 ;
  LAYER ME1 ;
  RECT 1821.600 0.000 1822.400 1.000 ;
 END
 ANTENNAPARTIALMETALAREA                  4.152 LAYER ME2 ;
 ANTENNADIFFAREA                          5.472 LAYER ME2 ;
 ANTENNADIFFAREA                          5.472 LAYER ME3 ;
 ANTENNADIFFAREA                          5.472 LAYER ME4 ;
END DO85
PIN DI85
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 1807.200 0.000 1808.000 1.000 ;
  LAYER ME3 ;
  RECT 1807.200 0.000 1808.000 1.000 ;
  LAYER ME2 ;
  RECT 1807.200 0.000 1808.000 1.000 ;
  LAYER ME1 ;
  RECT 1807.200 0.000 1808.000 1.000 ;
 END
 ANTENNAPARTIALMETALAREA                  3.150 LAYER ME2 ;
 ANTENNAGATEAREA                          0.086 LAYER ME2 ;
 ANTENNAGATEAREA                          0.086 LAYER ME3 ;
 ANTENNAGATEAREA                          0.086 LAYER ME4 ;
 ANTENNADIFFAREA                          0.160 LAYER ME2 ;
 ANTENNADIFFAREA                          0.160 LAYER ME3 ;
 ANTENNADIFFAREA                          0.160 LAYER ME4 ;
 ANTENNAMAXAREACAR                       48.801 LAYER ME2 ;
 ANTENNAMAXAREACAR                       58.060 LAYER ME3 ;
 ANTENNAMAXAREACAR                       67.319 LAYER ME4 ;
END DI85
PIN DO84
  DIRECTION OUTPUT ;
 PORT
  LAYER ME4 ;
  RECT 1802.000 0.000 1802.800 1.000 ;
  LAYER ME3 ;
  RECT 1802.000 0.000 1802.800 1.000 ;
  LAYER ME2 ;
  RECT 1802.000 0.000 1802.800 1.000 ;
  LAYER ME1 ;
  RECT 1802.000 0.000 1802.800 1.000 ;
 END
 ANTENNAPARTIALMETALAREA                  4.176 LAYER ME2 ;
 ANTENNADIFFAREA                          5.472 LAYER ME2 ;
 ANTENNADIFFAREA                          5.472 LAYER ME3 ;
 ANTENNADIFFAREA                          5.472 LAYER ME4 ;
END DO84
PIN DI84
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 1787.200 0.000 1788.000 1.000 ;
  LAYER ME3 ;
  RECT 1787.200 0.000 1788.000 1.000 ;
  LAYER ME2 ;
  RECT 1787.200 0.000 1788.000 1.000 ;
  LAYER ME1 ;
  RECT 1787.200 0.000 1788.000 1.000 ;
 END
 ANTENNAPARTIALMETALAREA                  3.118 LAYER ME2 ;
 ANTENNAGATEAREA                          0.086 LAYER ME2 ;
 ANTENNAGATEAREA                          0.086 LAYER ME3 ;
 ANTENNAGATEAREA                          0.086 LAYER ME4 ;
 ANTENNADIFFAREA                          0.160 LAYER ME2 ;
 ANTENNADIFFAREA                          0.160 LAYER ME3 ;
 ANTENNADIFFAREA                          0.160 LAYER ME4 ;
 ANTENNAMAXAREACAR                       48.431 LAYER ME2 ;
 ANTENNAMAXAREACAR                       57.690 LAYER ME3 ;
 ANTENNAMAXAREACAR                       66.949 LAYER ME4 ;
END DI84
PIN DO83
  DIRECTION OUTPUT ;
 PORT
  LAYER ME4 ;
  RECT 1780.800 0.000 1781.600 1.000 ;
  LAYER ME3 ;
  RECT 1780.800 0.000 1781.600 1.000 ;
  LAYER ME2 ;
  RECT 1780.800 0.000 1781.600 1.000 ;
  LAYER ME1 ;
  RECT 1780.800 0.000 1781.600 1.000 ;
 END
 ANTENNAPARTIALMETALAREA                  4.152 LAYER ME2 ;
 ANTENNADIFFAREA                          5.472 LAYER ME2 ;
 ANTENNADIFFAREA                          5.472 LAYER ME3 ;
 ANTENNADIFFAREA                          5.472 LAYER ME4 ;
END DO83
PIN DI83
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 1766.000 0.000 1766.800 1.000 ;
  LAYER ME3 ;
  RECT 1766.000 0.000 1766.800 1.000 ;
  LAYER ME2 ;
  RECT 1766.000 0.000 1766.800 1.000 ;
  LAYER ME1 ;
  RECT 1766.000 0.000 1766.800 1.000 ;
 END
 ANTENNAPARTIALMETALAREA                  3.138 LAYER ME2 ;
 ANTENNAGATEAREA                          0.086 LAYER ME2 ;
 ANTENNAGATEAREA                          0.086 LAYER ME3 ;
 ANTENNAGATEAREA                          0.086 LAYER ME4 ;
 ANTENNADIFFAREA                          0.160 LAYER ME2 ;
 ANTENNADIFFAREA                          0.160 LAYER ME3 ;
 ANTENNADIFFAREA                          0.160 LAYER ME4 ;
 ANTENNAMAXAREACAR                       48.662 LAYER ME2 ;
 ANTENNAMAXAREACAR                       57.921 LAYER ME3 ;
 ANTENNAMAXAREACAR                       67.181 LAYER ME4 ;
END DI83
PIN DO82
  DIRECTION OUTPUT ;
 PORT
  LAYER ME4 ;
  RECT 1760.800 0.000 1761.600 1.000 ;
  LAYER ME3 ;
  RECT 1760.800 0.000 1761.600 1.000 ;
  LAYER ME2 ;
  RECT 1760.800 0.000 1761.600 1.000 ;
  LAYER ME1 ;
  RECT 1760.800 0.000 1761.600 1.000 ;
 END
 ANTENNAPARTIALMETALAREA                  4.160 LAYER ME2 ;
 ANTENNADIFFAREA                          5.472 LAYER ME2 ;
 ANTENNADIFFAREA                          5.472 LAYER ME3 ;
 ANTENNADIFFAREA                          5.472 LAYER ME4 ;
END DO82
PIN DI82
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 1746.400 0.000 1747.200 1.000 ;
  LAYER ME3 ;
  RECT 1746.400 0.000 1747.200 1.000 ;
  LAYER ME2 ;
  RECT 1746.400 0.000 1747.200 1.000 ;
  LAYER ME1 ;
  RECT 1746.400 0.000 1747.200 1.000 ;
 END
 ANTENNAPARTIALMETALAREA                  3.142 LAYER ME2 ;
 ANTENNAGATEAREA                          0.086 LAYER ME2 ;
 ANTENNAGATEAREA                          0.086 LAYER ME3 ;
 ANTENNAGATEAREA                          0.086 LAYER ME4 ;
 ANTENNADIFFAREA                          0.160 LAYER ME2 ;
 ANTENNADIFFAREA                          0.160 LAYER ME3 ;
 ANTENNADIFFAREA                          0.160 LAYER ME4 ;
 ANTENNAMAXAREACAR                       48.708 LAYER ME2 ;
 ANTENNAMAXAREACAR                       57.968 LAYER ME3 ;
 ANTENNAMAXAREACAR                       67.227 LAYER ME4 ;
END DI82
PIN DO81
  DIRECTION OUTPUT ;
 PORT
  LAYER ME4 ;
  RECT 1740.000 0.000 1740.800 1.000 ;
  LAYER ME3 ;
  RECT 1740.000 0.000 1740.800 1.000 ;
  LAYER ME2 ;
  RECT 1740.000 0.000 1740.800 1.000 ;
  LAYER ME1 ;
  RECT 1740.000 0.000 1740.800 1.000 ;
 END
 ANTENNAPARTIALMETALAREA                  4.176 LAYER ME2 ;
 ANTENNADIFFAREA                          5.472 LAYER ME2 ;
 ANTENNADIFFAREA                          5.472 LAYER ME3 ;
 ANTENNADIFFAREA                          5.472 LAYER ME4 ;
END DO81
PIN DI81
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 1725.200 0.000 1726.000 1.000 ;
  LAYER ME3 ;
  RECT 1725.200 0.000 1726.000 1.000 ;
  LAYER ME2 ;
  RECT 1725.200 0.000 1726.000 1.000 ;
  LAYER ME1 ;
  RECT 1725.200 0.000 1726.000 1.000 ;
 END
 ANTENNAPARTIALMETALAREA                  3.118 LAYER ME2 ;
 ANTENNAGATEAREA                          0.086 LAYER ME2 ;
 ANTENNAGATEAREA                          0.086 LAYER ME3 ;
 ANTENNAGATEAREA                          0.086 LAYER ME4 ;
 ANTENNADIFFAREA                          0.160 LAYER ME2 ;
 ANTENNADIFFAREA                          0.160 LAYER ME3 ;
 ANTENNADIFFAREA                          0.160 LAYER ME4 ;
 ANTENNAMAXAREACAR                       48.431 LAYER ME2 ;
 ANTENNAMAXAREACAR                       57.690 LAYER ME3 ;
 ANTENNAMAXAREACAR                       66.949 LAYER ME4 ;
END DI81
PIN DO80
  DIRECTION OUTPUT ;
 PORT
  LAYER ME4 ;
  RECT 1720.000 0.000 1720.800 1.000 ;
  LAYER ME3 ;
  RECT 1720.000 0.000 1720.800 1.000 ;
  LAYER ME2 ;
  RECT 1720.000 0.000 1720.800 1.000 ;
  LAYER ME1 ;
  RECT 1720.000 0.000 1720.800 1.000 ;
 END
 ANTENNAPARTIALMETALAREA                  4.144 LAYER ME2 ;
 ANTENNADIFFAREA                          5.472 LAYER ME2 ;
 ANTENNADIFFAREA                          5.472 LAYER ME3 ;
 ANTENNADIFFAREA                          5.472 LAYER ME4 ;
END DO80
PIN WEB10
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 1707.200 0.000 1708.000 1.000 ;
  LAYER ME3 ;
  RECT 1707.200 0.000 1708.000 1.000 ;
  LAYER ME2 ;
  RECT 1707.200 0.000 1708.000 1.000 ;
  LAYER ME1 ;
  RECT 1707.200 0.000 1708.000 1.000 ;
 END
 ANTENNAPARTIALMETALAREA                  2.856 LAYER ME2 ;
 ANTENNAGATEAREA                          0.072 LAYER ME2 ;
 ANTENNAGATEAREA                          0.072 LAYER ME3 ;
 ANTENNAGATEAREA                          0.072 LAYER ME4 ;
 ANTENNADIFFAREA                          0.160 LAYER ME2 ;
 ANTENNADIFFAREA                          0.160 LAYER ME3 ;
 ANTENNADIFFAREA                          0.160 LAYER ME4 ;
 ANTENNAMAXAREACAR                       54.678 LAYER ME2 ;
 ANTENNAMAXAREACAR                       65.789 LAYER ME3 ;
 ANTENNAMAXAREACAR                       76.900 LAYER ME4 ;
END WEB10
PIN DI80
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 1705.200 0.000 1706.000 1.000 ;
  LAYER ME3 ;
  RECT 1705.200 0.000 1706.000 1.000 ;
  LAYER ME2 ;
  RECT 1705.200 0.000 1706.000 1.000 ;
  LAYER ME1 ;
  RECT 1705.200 0.000 1706.000 1.000 ;
 END
 ANTENNAPARTIALMETALAREA                  3.146 LAYER ME2 ;
 ANTENNAGATEAREA                          0.086 LAYER ME2 ;
 ANTENNAGATEAREA                          0.086 LAYER ME3 ;
 ANTENNAGATEAREA                          0.086 LAYER ME4 ;
 ANTENNADIFFAREA                          0.160 LAYER ME2 ;
 ANTENNADIFFAREA                          0.160 LAYER ME3 ;
 ANTENNADIFFAREA                          0.160 LAYER ME4 ;
 ANTENNAMAXAREACAR                       48.755 LAYER ME2 ;
 ANTENNAMAXAREACAR                       58.014 LAYER ME3 ;
 ANTENNAMAXAREACAR                       67.273 LAYER ME4 ;
END DI80
PIN DO79
  DIRECTION OUTPUT ;
 PORT
  LAYER ME4 ;
  RECT 1698.800 0.000 1699.600 1.000 ;
  LAYER ME3 ;
  RECT 1698.800 0.000 1699.600 1.000 ;
  LAYER ME2 ;
  RECT 1698.800 0.000 1699.600 1.000 ;
  LAYER ME1 ;
  RECT 1698.800 0.000 1699.600 1.000 ;
 END
 ANTENNAPARTIALMETALAREA                  4.160 LAYER ME2 ;
 ANTENNADIFFAREA                          5.472 LAYER ME2 ;
 ANTENNADIFFAREA                          5.472 LAYER ME3 ;
 ANTENNADIFFAREA                          5.472 LAYER ME4 ;
END DO79
PIN DI79
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 1684.400 0.000 1685.200 1.000 ;
  LAYER ME3 ;
  RECT 1684.400 0.000 1685.200 1.000 ;
  LAYER ME2 ;
  RECT 1684.400 0.000 1685.200 1.000 ;
  LAYER ME1 ;
  RECT 1684.400 0.000 1685.200 1.000 ;
 END
 ANTENNAPARTIALMETALAREA                  3.142 LAYER ME2 ;
 ANTENNAGATEAREA                          0.086 LAYER ME2 ;
 ANTENNAGATEAREA                          0.086 LAYER ME3 ;
 ANTENNAGATEAREA                          0.086 LAYER ME4 ;
 ANTENNADIFFAREA                          0.160 LAYER ME2 ;
 ANTENNADIFFAREA                          0.160 LAYER ME3 ;
 ANTENNADIFFAREA                          0.160 LAYER ME4 ;
 ANTENNAMAXAREACAR                       48.708 LAYER ME2 ;
 ANTENNAMAXAREACAR                       57.968 LAYER ME3 ;
 ANTENNAMAXAREACAR                       67.227 LAYER ME4 ;
END DI79
PIN DO78
  DIRECTION OUTPUT ;
 PORT
  LAYER ME4 ;
  RECT 1679.200 0.000 1680.000 1.000 ;
  LAYER ME3 ;
  RECT 1679.200 0.000 1680.000 1.000 ;
  LAYER ME2 ;
  RECT 1679.200 0.000 1680.000 1.000 ;
  LAYER ME1 ;
  RECT 1679.200 0.000 1680.000 1.000 ;
 END
 ANTENNAPARTIALMETALAREA                  4.168 LAYER ME2 ;
 ANTENNADIFFAREA                          5.472 LAYER ME2 ;
 ANTENNADIFFAREA                          5.472 LAYER ME3 ;
 ANTENNADIFFAREA                          5.472 LAYER ME4 ;
END DO78
PIN DI78
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 1664.400 0.000 1665.200 1.000 ;
  LAYER ME3 ;
  RECT 1664.400 0.000 1665.200 1.000 ;
  LAYER ME2 ;
  RECT 1664.400 0.000 1665.200 1.000 ;
  LAYER ME1 ;
  RECT 1664.400 0.000 1665.200 1.000 ;
 END
 ANTENNAPARTIALMETALAREA                  3.122 LAYER ME2 ;
 ANTENNAGATEAREA                          0.086 LAYER ME2 ;
 ANTENNAGATEAREA                          0.086 LAYER ME3 ;
 ANTENNAGATEAREA                          0.086 LAYER ME4 ;
 ANTENNADIFFAREA                          0.160 LAYER ME2 ;
 ANTENNADIFFAREA                          0.160 LAYER ME3 ;
 ANTENNADIFFAREA                          0.160 LAYER ME4 ;
 ANTENNAMAXAREACAR                       48.477 LAYER ME2 ;
 ANTENNAMAXAREACAR                       57.736 LAYER ME3 ;
 ANTENNAMAXAREACAR                       66.995 LAYER ME4 ;
END DI78
PIN DO77
  DIRECTION OUTPUT ;
 PORT
  LAYER ME4 ;
  RECT 1658.000 0.000 1658.800 1.000 ;
  LAYER ME3 ;
  RECT 1658.000 0.000 1658.800 1.000 ;
  LAYER ME2 ;
  RECT 1658.000 0.000 1658.800 1.000 ;
  LAYER ME1 ;
  RECT 1658.000 0.000 1658.800 1.000 ;
 END
 ANTENNAPARTIALMETALAREA                  4.144 LAYER ME2 ;
 ANTENNADIFFAREA                          5.472 LAYER ME2 ;
 ANTENNADIFFAREA                          5.472 LAYER ME3 ;
 ANTENNADIFFAREA                          5.472 LAYER ME4 ;
END DO77
PIN DI77
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 1643.200 0.000 1644.000 1.000 ;
  LAYER ME3 ;
  RECT 1643.200 0.000 1644.000 1.000 ;
  LAYER ME2 ;
  RECT 1643.200 0.000 1644.000 1.000 ;
  LAYER ME1 ;
  RECT 1643.200 0.000 1644.000 1.000 ;
 END
 ANTENNAPARTIALMETALAREA                  3.146 LAYER ME2 ;
 ANTENNAGATEAREA                          0.086 LAYER ME2 ;
 ANTENNAGATEAREA                          0.086 LAYER ME3 ;
 ANTENNAGATEAREA                          0.086 LAYER ME4 ;
 ANTENNADIFFAREA                          0.160 LAYER ME2 ;
 ANTENNADIFFAREA                          0.160 LAYER ME3 ;
 ANTENNADIFFAREA                          0.160 LAYER ME4 ;
 ANTENNAMAXAREACAR                       48.755 LAYER ME2 ;
 ANTENNAMAXAREACAR                       58.014 LAYER ME3 ;
 ANTENNAMAXAREACAR                       67.273 LAYER ME4 ;
END DI77
PIN DO76
  DIRECTION OUTPUT ;
 PORT
  LAYER ME4 ;
  RECT 1638.000 0.000 1638.800 1.000 ;
  LAYER ME3 ;
  RECT 1638.000 0.000 1638.800 1.000 ;
  LAYER ME2 ;
  RECT 1638.000 0.000 1638.800 1.000 ;
  LAYER ME1 ;
  RECT 1638.000 0.000 1638.800 1.000 ;
 END
 ANTENNAPARTIALMETALAREA                  4.168 LAYER ME2 ;
 ANTENNADIFFAREA                          5.472 LAYER ME2 ;
 ANTENNADIFFAREA                          5.472 LAYER ME3 ;
 ANTENNADIFFAREA                          5.472 LAYER ME4 ;
END DO76
PIN DI76
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 1623.600 0.000 1624.400 1.000 ;
  LAYER ME3 ;
  RECT 1623.600 0.000 1624.400 1.000 ;
  LAYER ME2 ;
  RECT 1623.600 0.000 1624.400 1.000 ;
  LAYER ME1 ;
  RECT 1623.600 0.000 1624.400 1.000 ;
 END
 ANTENNAPARTIALMETALAREA                  3.134 LAYER ME2 ;
 ANTENNAGATEAREA                          0.086 LAYER ME2 ;
 ANTENNAGATEAREA                          0.086 LAYER ME3 ;
 ANTENNAGATEAREA                          0.086 LAYER ME4 ;
 ANTENNADIFFAREA                          0.160 LAYER ME2 ;
 ANTENNADIFFAREA                          0.160 LAYER ME3 ;
 ANTENNADIFFAREA                          0.160 LAYER ME4 ;
 ANTENNAMAXAREACAR                       48.616 LAYER ME2 ;
 ANTENNAMAXAREACAR                       57.875 LAYER ME3 ;
 ANTENNAMAXAREACAR                       67.134 LAYER ME4 ;
END DI76
PIN DO75
  DIRECTION OUTPUT ;
 PORT
  LAYER ME4 ;
  RECT 1617.200 0.000 1618.000 1.000 ;
  LAYER ME3 ;
  RECT 1617.200 0.000 1618.000 1.000 ;
  LAYER ME2 ;
  RECT 1617.200 0.000 1618.000 1.000 ;
  LAYER ME1 ;
  RECT 1617.200 0.000 1618.000 1.000 ;
 END
 ANTENNAPARTIALMETALAREA                  4.168 LAYER ME2 ;
 ANTENNADIFFAREA                          5.472 LAYER ME2 ;
 ANTENNADIFFAREA                          5.472 LAYER ME3 ;
 ANTENNADIFFAREA                          5.472 LAYER ME4 ;
END DO75
PIN DI75
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 1602.400 0.000 1603.200 1.000 ;
  LAYER ME3 ;
  RECT 1602.400 0.000 1603.200 1.000 ;
  LAYER ME2 ;
  RECT 1602.400 0.000 1603.200 1.000 ;
  LAYER ME1 ;
  RECT 1602.400 0.000 1603.200 1.000 ;
 END
 ANTENNAPARTIALMETALAREA                  3.122 LAYER ME2 ;
 ANTENNAGATEAREA                          0.086 LAYER ME2 ;
 ANTENNAGATEAREA                          0.086 LAYER ME3 ;
 ANTENNAGATEAREA                          0.086 LAYER ME4 ;
 ANTENNADIFFAREA                          0.160 LAYER ME2 ;
 ANTENNADIFFAREA                          0.160 LAYER ME3 ;
 ANTENNADIFFAREA                          0.160 LAYER ME4 ;
 ANTENNAMAXAREACAR                       48.477 LAYER ME2 ;
 ANTENNAMAXAREACAR                       57.736 LAYER ME3 ;
 ANTENNAMAXAREACAR                       66.995 LAYER ME4 ;
END DI75
PIN DO74
  DIRECTION OUTPUT ;
 PORT
  LAYER ME4 ;
  RECT 1597.200 0.000 1598.000 1.000 ;
  LAYER ME3 ;
  RECT 1597.200 0.000 1598.000 1.000 ;
  LAYER ME2 ;
  RECT 1597.200 0.000 1598.000 1.000 ;
  LAYER ME1 ;
  RECT 1597.200 0.000 1598.000 1.000 ;
 END
 ANTENNAPARTIALMETALAREA                  4.144 LAYER ME2 ;
 ANTENNADIFFAREA                          5.472 LAYER ME2 ;
 ANTENNADIFFAREA                          5.472 LAYER ME3 ;
 ANTENNADIFFAREA                          5.472 LAYER ME4 ;
END DO74
PIN DI74
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 1582.400 0.000 1583.200 1.000 ;
  LAYER ME3 ;
  RECT 1582.400 0.000 1583.200 1.000 ;
  LAYER ME2 ;
  RECT 1582.400 0.000 1583.200 1.000 ;
  LAYER ME1 ;
  RECT 1582.400 0.000 1583.200 1.000 ;
 END
 ANTENNAPARTIALMETALAREA                  3.154 LAYER ME2 ;
 ANTENNAGATEAREA                          0.086 LAYER ME2 ;
 ANTENNAGATEAREA                          0.086 LAYER ME3 ;
 ANTENNAGATEAREA                          0.086 LAYER ME4 ;
 ANTENNADIFFAREA                          0.160 LAYER ME2 ;
 ANTENNADIFFAREA                          0.160 LAYER ME3 ;
 ANTENNADIFFAREA                          0.160 LAYER ME4 ;
 ANTENNAMAXAREACAR                       48.847 LAYER ME2 ;
 ANTENNAMAXAREACAR                       58.106 LAYER ME3 ;
 ANTENNAMAXAREACAR                       67.366 LAYER ME4 ;
END DI74
PIN DO73
  DIRECTION OUTPUT ;
 PORT
  LAYER ME4 ;
  RECT 1576.000 0.000 1576.800 1.000 ;
  LAYER ME3 ;
  RECT 1576.000 0.000 1576.800 1.000 ;
  LAYER ME2 ;
  RECT 1576.000 0.000 1576.800 1.000 ;
  LAYER ME1 ;
  RECT 1576.000 0.000 1576.800 1.000 ;
 END
 ANTENNAPARTIALMETALAREA                  4.168 LAYER ME2 ;
 ANTENNADIFFAREA                          5.472 LAYER ME2 ;
 ANTENNADIFFAREA                          5.472 LAYER ME3 ;
 ANTENNADIFFAREA                          5.472 LAYER ME4 ;
END DO73
PIN DI73
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 1561.600 0.000 1562.400 1.000 ;
  LAYER ME3 ;
  RECT 1561.600 0.000 1562.400 1.000 ;
  LAYER ME2 ;
  RECT 1561.600 0.000 1562.400 1.000 ;
  LAYER ME1 ;
  RECT 1561.600 0.000 1562.400 1.000 ;
 END
 ANTENNAPARTIALMETALAREA                  3.134 LAYER ME2 ;
 ANTENNAGATEAREA                          0.086 LAYER ME2 ;
 ANTENNAGATEAREA                          0.086 LAYER ME3 ;
 ANTENNAGATEAREA                          0.086 LAYER ME4 ;
 ANTENNADIFFAREA                          0.160 LAYER ME2 ;
 ANTENNADIFFAREA                          0.160 LAYER ME3 ;
 ANTENNADIFFAREA                          0.160 LAYER ME4 ;
 ANTENNAMAXAREACAR                       48.616 LAYER ME2 ;
 ANTENNAMAXAREACAR                       57.875 LAYER ME3 ;
 ANTENNAMAXAREACAR                       67.134 LAYER ME4 ;
END DI73
PIN DO72
  DIRECTION OUTPUT ;
 PORT
  LAYER ME4 ;
  RECT 1556.400 0.000 1557.200 1.000 ;
  LAYER ME3 ;
  RECT 1556.400 0.000 1557.200 1.000 ;
  LAYER ME2 ;
  RECT 1556.400 0.000 1557.200 1.000 ;
  LAYER ME1 ;
  RECT 1556.400 0.000 1557.200 1.000 ;
 END
 ANTENNAPARTIALMETALAREA                  4.160 LAYER ME2 ;
 ANTENNADIFFAREA                          5.472 LAYER ME2 ;
 ANTENNADIFFAREA                          5.472 LAYER ME3 ;
 ANTENNADIFFAREA                          5.472 LAYER ME4 ;
END DO72
PIN WEB9
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 1543.200 0.000 1544.000 1.000 ;
  LAYER ME3 ;
  RECT 1543.200 0.000 1544.000 1.000 ;
  LAYER ME2 ;
  RECT 1543.200 0.000 1544.000 1.000 ;
  LAYER ME1 ;
  RECT 1543.200 0.000 1544.000 1.000 ;
 END
 ANTENNAPARTIALMETALAREA                  2.868 LAYER ME2 ;
 ANTENNAGATEAREA                          0.072 LAYER ME2 ;
 ANTENNAGATEAREA                          0.072 LAYER ME3 ;
 ANTENNAGATEAREA                          0.072 LAYER ME4 ;
 ANTENNADIFFAREA                          0.160 LAYER ME2 ;
 ANTENNADIFFAREA                          0.160 LAYER ME3 ;
 ANTENNADIFFAREA                          0.160 LAYER ME4 ;
 ANTENNAMAXAREACAR                       54.844 LAYER ME2 ;
 ANTENNAMAXAREACAR                       65.956 LAYER ME3 ;
 ANTENNAMAXAREACAR                       77.067 LAYER ME4 ;
END WEB9
PIN DI72
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 1541.600 0.000 1542.400 1.000 ;
  LAYER ME3 ;
  RECT 1541.600 0.000 1542.400 1.000 ;
  LAYER ME2 ;
  RECT 1541.600 0.000 1542.400 1.000 ;
  LAYER ME1 ;
  RECT 1541.600 0.000 1542.400 1.000 ;
 END
 ANTENNAPARTIALMETALAREA                  3.130 LAYER ME2 ;
 ANTENNAGATEAREA                          0.086 LAYER ME2 ;
 ANTENNAGATEAREA                          0.086 LAYER ME3 ;
 ANTENNAGATEAREA                          0.086 LAYER ME4 ;
 ANTENNADIFFAREA                          0.160 LAYER ME2 ;
 ANTENNADIFFAREA                          0.160 LAYER ME3 ;
 ANTENNADIFFAREA                          0.160 LAYER ME4 ;
 ANTENNAMAXAREACAR                       48.569 LAYER ME2 ;
 ANTENNAMAXAREACAR                       57.829 LAYER ME3 ;
 ANTENNAMAXAREACAR                       67.088 LAYER ME4 ;
END DI72
PIN DO71
  DIRECTION OUTPUT ;
 PORT
  LAYER ME4 ;
  RECT 1535.200 0.000 1536.000 1.000 ;
  LAYER ME3 ;
  RECT 1535.200 0.000 1536.000 1.000 ;
  LAYER ME2 ;
  RECT 1535.200 0.000 1536.000 1.000 ;
  LAYER ME1 ;
  RECT 1535.200 0.000 1536.000 1.000 ;
 END
 ANTENNAPARTIALMETALAREA                  4.144 LAYER ME2 ;
 ANTENNADIFFAREA                          5.472 LAYER ME2 ;
 ANTENNADIFFAREA                          5.472 LAYER ME3 ;
 ANTENNADIFFAREA                          5.472 LAYER ME4 ;
END DO71
PIN DI71
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 1520.400 0.000 1521.200 1.000 ;
  LAYER ME3 ;
  RECT 1520.400 0.000 1521.200 1.000 ;
  LAYER ME2 ;
  RECT 1520.400 0.000 1521.200 1.000 ;
  LAYER ME1 ;
  RECT 1520.400 0.000 1521.200 1.000 ;
 END
 ANTENNAPARTIALMETALAREA                  3.154 LAYER ME2 ;
 ANTENNAGATEAREA                          0.086 LAYER ME2 ;
 ANTENNAGATEAREA                          0.086 LAYER ME3 ;
 ANTENNAGATEAREA                          0.086 LAYER ME4 ;
 ANTENNADIFFAREA                          0.160 LAYER ME2 ;
 ANTENNADIFFAREA                          0.160 LAYER ME3 ;
 ANTENNADIFFAREA                          0.160 LAYER ME4 ;
 ANTENNAMAXAREACAR                       48.847 LAYER ME2 ;
 ANTENNAMAXAREACAR                       58.106 LAYER ME3 ;
 ANTENNAMAXAREACAR                       67.366 LAYER ME4 ;
END DI71
PIN DO70
  DIRECTION OUTPUT ;
 PORT
  LAYER ME4 ;
  RECT 1515.200 0.000 1516.000 1.000 ;
  LAYER ME3 ;
  RECT 1515.200 0.000 1516.000 1.000 ;
  LAYER ME2 ;
  RECT 1515.200 0.000 1516.000 1.000 ;
  LAYER ME1 ;
  RECT 1515.200 0.000 1516.000 1.000 ;
 END
 ANTENNAPARTIALMETALAREA                  4.176 LAYER ME2 ;
 ANTENNADIFFAREA                          5.472 LAYER ME2 ;
 ANTENNADIFFAREA                          5.472 LAYER ME3 ;
 ANTENNADIFFAREA                          5.472 LAYER ME4 ;
END DO70
PIN DI70
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 1500.800 0.000 1501.600 1.000 ;
  LAYER ME3 ;
  RECT 1500.800 0.000 1501.600 1.000 ;
  LAYER ME2 ;
  RECT 1500.800 0.000 1501.600 1.000 ;
  LAYER ME1 ;
  RECT 1500.800 0.000 1501.600 1.000 ;
 END
 ANTENNAPARTIALMETALAREA                  3.126 LAYER ME2 ;
 ANTENNAGATEAREA                          0.086 LAYER ME2 ;
 ANTENNAGATEAREA                          0.086 LAYER ME3 ;
 ANTENNAGATEAREA                          0.086 LAYER ME4 ;
 ANTENNADIFFAREA                          0.160 LAYER ME2 ;
 ANTENNADIFFAREA                          0.160 LAYER ME3 ;
 ANTENNADIFFAREA                          0.160 LAYER ME4 ;
 ANTENNAMAXAREACAR                       48.523 LAYER ME2 ;
 ANTENNAMAXAREACAR                       57.782 LAYER ME3 ;
 ANTENNAMAXAREACAR                       67.042 LAYER ME4 ;
END DI70
PIN DO69
  DIRECTION OUTPUT ;
 PORT
  LAYER ME4 ;
  RECT 1494.400 0.000 1495.200 1.000 ;
  LAYER ME3 ;
  RECT 1494.400 0.000 1495.200 1.000 ;
  LAYER ME2 ;
  RECT 1494.400 0.000 1495.200 1.000 ;
  LAYER ME1 ;
  RECT 1494.400 0.000 1495.200 1.000 ;
 END
 ANTENNAPARTIALMETALAREA                  4.160 LAYER ME2 ;
 ANTENNADIFFAREA                          5.472 LAYER ME2 ;
 ANTENNADIFFAREA                          5.472 LAYER ME3 ;
 ANTENNADIFFAREA                          5.472 LAYER ME4 ;
END DO69
PIN DI69
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 1479.600 0.000 1480.400 1.000 ;
  LAYER ME3 ;
  RECT 1479.600 0.000 1480.400 1.000 ;
  LAYER ME2 ;
  RECT 1479.600 0.000 1480.400 1.000 ;
  LAYER ME1 ;
  RECT 1479.600 0.000 1480.400 1.000 ;
 END
 ANTENNAPARTIALMETALAREA                  3.130 LAYER ME2 ;
 ANTENNAGATEAREA                          0.086 LAYER ME2 ;
 ANTENNAGATEAREA                          0.086 LAYER ME3 ;
 ANTENNAGATEAREA                          0.086 LAYER ME4 ;
 ANTENNADIFFAREA                          0.160 LAYER ME2 ;
 ANTENNADIFFAREA                          0.160 LAYER ME3 ;
 ANTENNADIFFAREA                          0.160 LAYER ME4 ;
 ANTENNAMAXAREACAR                       48.569 LAYER ME2 ;
 ANTENNAMAXAREACAR                       57.829 LAYER ME3 ;
 ANTENNAMAXAREACAR                       67.088 LAYER ME4 ;
END DI69
PIN DO68
  DIRECTION OUTPUT ;
 PORT
  LAYER ME4 ;
  RECT 1474.400 0.000 1475.200 1.000 ;
  LAYER ME3 ;
  RECT 1474.400 0.000 1475.200 1.000 ;
  LAYER ME2 ;
  RECT 1474.400 0.000 1475.200 1.000 ;
  LAYER ME1 ;
  RECT 1474.400 0.000 1475.200 1.000 ;
 END
 ANTENNAPARTIALMETALAREA                  4.152 LAYER ME2 ;
 ANTENNADIFFAREA                          5.472 LAYER ME2 ;
 ANTENNADIFFAREA                          5.472 LAYER ME3 ;
 ANTENNADIFFAREA                          5.472 LAYER ME4 ;
END DO68
PIN DI68
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 1460.000 0.000 1460.800 1.000 ;
  LAYER ME3 ;
  RECT 1460.000 0.000 1460.800 1.000 ;
  LAYER ME2 ;
  RECT 1460.000 0.000 1460.800 1.000 ;
  LAYER ME1 ;
  RECT 1460.000 0.000 1460.800 1.000 ;
 END
 ANTENNAPARTIALMETALAREA                  3.150 LAYER ME2 ;
 ANTENNAGATEAREA                          0.086 LAYER ME2 ;
 ANTENNAGATEAREA                          0.086 LAYER ME3 ;
 ANTENNAGATEAREA                          0.086 LAYER ME4 ;
 ANTENNADIFFAREA                          0.160 LAYER ME2 ;
 ANTENNADIFFAREA                          0.160 LAYER ME3 ;
 ANTENNADIFFAREA                          0.160 LAYER ME4 ;
 ANTENNAMAXAREACAR                       48.801 LAYER ME2 ;
 ANTENNAMAXAREACAR                       58.060 LAYER ME3 ;
 ANTENNAMAXAREACAR                       67.319 LAYER ME4 ;
END DI68
PIN DO67
  DIRECTION OUTPUT ;
 PORT
  LAYER ME4 ;
  RECT 1453.200 0.000 1454.000 1.000 ;
  LAYER ME3 ;
  RECT 1453.200 0.000 1454.000 1.000 ;
  LAYER ME2 ;
  RECT 1453.200 0.000 1454.000 1.000 ;
  LAYER ME1 ;
  RECT 1453.200 0.000 1454.000 1.000 ;
 END
 ANTENNAPARTIALMETALAREA                  4.176 LAYER ME2 ;
 ANTENNADIFFAREA                          5.472 LAYER ME2 ;
 ANTENNADIFFAREA                          5.472 LAYER ME3 ;
 ANTENNADIFFAREA                          5.472 LAYER ME4 ;
END DO67
PIN DI67
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 1438.800 0.000 1439.600 1.000 ;
  LAYER ME3 ;
  RECT 1438.800 0.000 1439.600 1.000 ;
  LAYER ME2 ;
  RECT 1438.800 0.000 1439.600 1.000 ;
  LAYER ME1 ;
  RECT 1438.800 0.000 1439.600 1.000 ;
 END
 ANTENNAPARTIALMETALAREA                  3.126 LAYER ME2 ;
 ANTENNAGATEAREA                          0.086 LAYER ME2 ;
 ANTENNAGATEAREA                          0.086 LAYER ME3 ;
 ANTENNAGATEAREA                          0.086 LAYER ME4 ;
 ANTENNADIFFAREA                          0.160 LAYER ME2 ;
 ANTENNADIFFAREA                          0.160 LAYER ME3 ;
 ANTENNADIFFAREA                          0.160 LAYER ME4 ;
 ANTENNAMAXAREACAR                       48.523 LAYER ME2 ;
 ANTENNAMAXAREACAR                       57.782 LAYER ME3 ;
 ANTENNAMAXAREACAR                       67.042 LAYER ME4 ;
END DI67
PIN DO66
  DIRECTION OUTPUT ;
 PORT
  LAYER ME4 ;
  RECT 1433.600 0.000 1434.400 1.000 ;
  LAYER ME3 ;
  RECT 1433.600 0.000 1434.400 1.000 ;
  LAYER ME2 ;
  RECT 1433.600 0.000 1434.400 1.000 ;
  LAYER ME1 ;
  RECT 1433.600 0.000 1434.400 1.000 ;
 END
 ANTENNAPARTIALMETALAREA                  4.152 LAYER ME2 ;
 ANTENNADIFFAREA                          5.472 LAYER ME2 ;
 ANTENNADIFFAREA                          5.472 LAYER ME3 ;
 ANTENNADIFFAREA                          5.472 LAYER ME4 ;
END DO66
PIN DI66
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 1418.800 0.000 1419.600 1.000 ;
  LAYER ME3 ;
  RECT 1418.800 0.000 1419.600 1.000 ;
  LAYER ME2 ;
  RECT 1418.800 0.000 1419.600 1.000 ;
  LAYER ME1 ;
  RECT 1418.800 0.000 1419.600 1.000 ;
 END
 ANTENNAPARTIALMETALAREA                  3.138 LAYER ME2 ;
 ANTENNAGATEAREA                          0.086 LAYER ME2 ;
 ANTENNAGATEAREA                          0.086 LAYER ME3 ;
 ANTENNAGATEAREA                          0.086 LAYER ME4 ;
 ANTENNADIFFAREA                          0.160 LAYER ME2 ;
 ANTENNADIFFAREA                          0.160 LAYER ME3 ;
 ANTENNADIFFAREA                          0.160 LAYER ME4 ;
 ANTENNAMAXAREACAR                       48.662 LAYER ME2 ;
 ANTENNAMAXAREACAR                       57.921 LAYER ME3 ;
 ANTENNAMAXAREACAR                       67.181 LAYER ME4 ;
END DI66
PIN DO65
  DIRECTION OUTPUT ;
 PORT
  LAYER ME4 ;
  RECT 1412.400 0.000 1413.200 1.000 ;
  LAYER ME3 ;
  RECT 1412.400 0.000 1413.200 1.000 ;
  LAYER ME2 ;
  RECT 1412.400 0.000 1413.200 1.000 ;
  LAYER ME1 ;
  RECT 1412.400 0.000 1413.200 1.000 ;
 END
 ANTENNAPARTIALMETALAREA                  4.152 LAYER ME2 ;
 ANTENNADIFFAREA                          5.472 LAYER ME2 ;
 ANTENNADIFFAREA                          5.472 LAYER ME3 ;
 ANTENNADIFFAREA                          5.472 LAYER ME4 ;
END DO65
PIN DI65
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 1398.000 0.000 1398.800 1.000 ;
  LAYER ME3 ;
  RECT 1398.000 0.000 1398.800 1.000 ;
  LAYER ME2 ;
  RECT 1398.000 0.000 1398.800 1.000 ;
  LAYER ME1 ;
  RECT 1398.000 0.000 1398.800 1.000 ;
 END
 ANTENNAPARTIALMETALAREA                  3.150 LAYER ME2 ;
 ANTENNAGATEAREA                          0.086 LAYER ME2 ;
 ANTENNAGATEAREA                          0.086 LAYER ME3 ;
 ANTENNAGATEAREA                          0.086 LAYER ME4 ;
 ANTENNADIFFAREA                          0.160 LAYER ME2 ;
 ANTENNADIFFAREA                          0.160 LAYER ME3 ;
 ANTENNADIFFAREA                          0.160 LAYER ME4 ;
 ANTENNAMAXAREACAR                       48.801 LAYER ME2 ;
 ANTENNAMAXAREACAR                       58.060 LAYER ME3 ;
 ANTENNAMAXAREACAR                       67.319 LAYER ME4 ;
END DI65
PIN DO64
  DIRECTION OUTPUT ;
 PORT
  LAYER ME4 ;
  RECT 1392.800 0.000 1393.600 1.000 ;
  LAYER ME3 ;
  RECT 1392.800 0.000 1393.600 1.000 ;
  LAYER ME2 ;
  RECT 1392.800 0.000 1393.600 1.000 ;
  LAYER ME1 ;
  RECT 1392.800 0.000 1393.600 1.000 ;
 END
 ANTENNAPARTIALMETALAREA                  4.176 LAYER ME2 ;
 ANTENNADIFFAREA                          5.472 LAYER ME2 ;
 ANTENNADIFFAREA                          5.472 LAYER ME3 ;
 ANTENNADIFFAREA                          5.472 LAYER ME4 ;
END DO64
PIN WEB8
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 1379.600 0.000 1380.400 1.000 ;
  LAYER ME3 ;
  RECT 1379.600 0.000 1380.400 1.000 ;
  LAYER ME2 ;
  RECT 1379.600 0.000 1380.400 1.000 ;
  LAYER ME1 ;
  RECT 1379.600 0.000 1380.400 1.000 ;
 END
 ANTENNAPARTIALMETALAREA                  2.852 LAYER ME2 ;
 ANTENNAGATEAREA                          0.072 LAYER ME2 ;
 ANTENNAGATEAREA                          0.072 LAYER ME3 ;
 ANTENNAGATEAREA                          0.072 LAYER ME4 ;
 ANTENNADIFFAREA                          0.160 LAYER ME2 ;
 ANTENNADIFFAREA                          0.160 LAYER ME3 ;
 ANTENNADIFFAREA                          0.160 LAYER ME4 ;
 ANTENNAMAXAREACAR                       54.622 LAYER ME2 ;
 ANTENNAMAXAREACAR                       65.733 LAYER ME3 ;
 ANTENNAMAXAREACAR                       76.844 LAYER ME4 ;
END WEB8
PIN DI64
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 1378.000 0.000 1378.800 1.000 ;
  LAYER ME3 ;
  RECT 1378.000 0.000 1378.800 1.000 ;
  LAYER ME2 ;
  RECT 1378.000 0.000 1378.800 1.000 ;
  LAYER ME1 ;
  RECT 1378.000 0.000 1378.800 1.000 ;
 END
 ANTENNAPARTIALMETALAREA                  3.118 LAYER ME2 ;
 ANTENNAGATEAREA                          0.086 LAYER ME2 ;
 ANTENNAGATEAREA                          0.086 LAYER ME3 ;
 ANTENNAGATEAREA                          0.086 LAYER ME4 ;
 ANTENNADIFFAREA                          0.160 LAYER ME2 ;
 ANTENNADIFFAREA                          0.160 LAYER ME3 ;
 ANTENNADIFFAREA                          0.160 LAYER ME4 ;
 ANTENNAMAXAREACAR                       48.431 LAYER ME2 ;
 ANTENNAMAXAREACAR                       57.690 LAYER ME3 ;
 ANTENNAMAXAREACAR                       66.949 LAYER ME4 ;
END DI64
PIN A3
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 1357.200 0.000 1358.000 1.000 ;
  LAYER ME3 ;
  RECT 1357.200 0.000 1358.000 1.000 ;
  LAYER ME2 ;
  RECT 1357.200 0.000 1358.000 1.000 ;
  LAYER ME1 ;
  RECT 1357.200 0.000 1358.000 1.000 ;
 END
 ANTENNAPARTIALMETALAREA                  2.028 LAYER ME2 ;
 ANTENNAGATEAREA                          0.180 LAYER ME2 ;
 ANTENNAGATEAREA                          0.180 LAYER ME3 ;
 ANTENNAGATEAREA                          0.180 LAYER ME4 ;
 ANTENNADIFFAREA                          0.160 LAYER ME2 ;
 ANTENNADIFFAREA                          0.160 LAYER ME3 ;
 ANTENNADIFFAREA                          0.160 LAYER ME4 ;
 ANTENNAMAXAREACAR                       17.116 LAYER ME2 ;
 ANTENNAMAXAREACAR                       21.560 LAYER ME3 ;
 ANTENNAMAXAREACAR                       26.004 LAYER ME4 ;
END A3
PIN A1
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 1356.000 0.000 1356.800 1.000 ;
  LAYER ME3 ;
  RECT 1356.000 0.000 1356.800 1.000 ;
  LAYER ME2 ;
  RECT 1356.000 0.000 1356.800 1.000 ;
  LAYER ME1 ;
  RECT 1356.000 0.000 1356.800 1.000 ;
 END
 ANTENNAPARTIALMETALAREA                  7.298 LAYER ME2 ;
 ANTENNAGATEAREA                          0.192 LAYER ME2 ;
 ANTENNAGATEAREA                          0.192 LAYER ME3 ;
 ANTENNAGATEAREA                          0.192 LAYER ME4 ;
 ANTENNADIFFAREA                          0.160 LAYER ME2 ;
 ANTENNADIFFAREA                          0.160 LAYER ME3 ;
 ANTENNADIFFAREA                          0.160 LAYER ME4 ;
 ANTENNAMAXAREACAR                       43.452 LAYER ME2 ;
 ANTENNAMAXAREACAR                       47.619 LAYER ME3 ;
 ANTENNAMAXAREACAR                       51.785 LAYER ME4 ;
END A1
PIN OE
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 1354.800 0.000 1355.600 1.000 ;
  LAYER ME3 ;
  RECT 1354.800 0.000 1355.600 1.000 ;
  LAYER ME2 ;
  RECT 1354.800 0.000 1355.600 1.000 ;
  LAYER ME1 ;
  RECT 1354.800 0.000 1355.600 1.000 ;
 END
 ANTENNAPARTIALMETALAREA                  3.370 LAYER ME2 ;
 ANTENNAGATEAREA                          0.840 LAYER ME2 ;
 ANTENNAGATEAREA                          0.840 LAYER ME3 ;
 ANTENNAGATEAREA                          0.840 LAYER ME4 ;
 ANTENNADIFFAREA                          0.160 LAYER ME2 ;
 ANTENNADIFFAREA                          0.160 LAYER ME3 ;
 ANTENNADIFFAREA                          0.160 LAYER ME4 ;
 ANTENNAMAXAREACAR                        5.336 LAYER ME2 ;
 ANTENNAMAXAREACAR                        6.288 LAYER ME3 ;
 ANTENNAMAXAREACAR                        7.240 LAYER ME4 ;
END OE
PIN CS
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 1353.600 0.000 1354.400 1.000 ;
  LAYER ME3 ;
  RECT 1353.600 0.000 1354.400 1.000 ;
  LAYER ME2 ;
  RECT 1353.600 0.000 1354.400 1.000 ;
  LAYER ME1 ;
  RECT 1353.600 0.000 1354.400 1.000 ;
 END
 ANTENNAPARTIALMETALAREA                  5.076 LAYER ME2 ;
 ANTENNAGATEAREA                          1.680 LAYER ME2 ;
 ANTENNAGATEAREA                          1.680 LAYER ME3 ;
 ANTENNAGATEAREA                          1.680 LAYER ME4 ;
 ANTENNADIFFAREA                          0.160 LAYER ME2 ;
 ANTENNADIFFAREA                          0.160 LAYER ME3 ;
 ANTENNADIFFAREA                          0.160 LAYER ME4 ;
 ANTENNAMAXAREACAR                        3.648 LAYER ME2 ;
 ANTENNAMAXAREACAR                        4.124 LAYER ME3 ;
 ANTENNAMAXAREACAR                        4.600 LAYER ME4 ;
END CS
PIN A2
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 1352.400 0.000 1353.200 1.000 ;
  LAYER ME3 ;
  RECT 1352.400 0.000 1353.200 1.000 ;
  LAYER ME2 ;
  RECT 1352.400 0.000 1353.200 1.000 ;
  LAYER ME1 ;
  RECT 1352.400 0.000 1353.200 1.000 ;
 END
 ANTENNAPARTIALMETALAREA                  7.366 LAYER ME2 ;
 ANTENNAGATEAREA                          0.192 LAYER ME2 ;
 ANTENNAGATEAREA                          0.192 LAYER ME3 ;
 ANTENNAGATEAREA                          0.192 LAYER ME4 ;
 ANTENNADIFFAREA                          0.160 LAYER ME2 ;
 ANTENNADIFFAREA                          0.160 LAYER ME3 ;
 ANTENNADIFFAREA                          0.160 LAYER ME4 ;
 ANTENNAMAXAREACAR                       43.806 LAYER ME2 ;
 ANTENNAMAXAREACAR                       47.973 LAYER ME3 ;
 ANTENNAMAXAREACAR                       52.140 LAYER ME4 ;
END A2
PIN A0
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 1351.200 0.000 1352.000 1.000 ;
  LAYER ME3 ;
  RECT 1351.200 0.000 1352.000 1.000 ;
  LAYER ME2 ;
  RECT 1351.200 0.000 1352.000 1.000 ;
  LAYER ME1 ;
  RECT 1351.200 0.000 1352.000 1.000 ;
 END
 ANTENNAPARTIALMETALAREA                  7.418 LAYER ME2 ;
 ANTENNAGATEAREA                          0.192 LAYER ME2 ;
 ANTENNAGATEAREA                          0.192 LAYER ME3 ;
 ANTENNAGATEAREA                          0.192 LAYER ME4 ;
 ANTENNADIFFAREA                          0.160 LAYER ME2 ;
 ANTENNADIFFAREA                          0.160 LAYER ME3 ;
 ANTENNADIFFAREA                          0.160 LAYER ME4 ;
 ANTENNAMAXAREACAR                       44.077 LAYER ME2 ;
 ANTENNAMAXAREACAR                       48.244 LAYER ME3 ;
 ANTENNAMAXAREACAR                       52.410 LAYER ME4 ;
END A0
PIN CK
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 1345.200 0.000 1346.000 1.000 ;
  LAYER ME3 ;
  RECT 1345.200 0.000 1346.000 1.000 ;
  LAYER ME2 ;
  RECT 1345.200 0.000 1346.000 1.000 ;
  LAYER ME1 ;
  RECT 1345.200 0.000 1346.000 1.000 ;
 END
 ANTENNAPARTIALMETALAREA                  5.506 LAYER ME2 ;
 ANTENNAGATEAREA                          1.908 LAYER ME2 ;
 ANTENNAGATEAREA                          1.908 LAYER ME3 ;
 ANTENNAGATEAREA                          1.908 LAYER ME4 ;
 ANTENNADIFFAREA                          0.160 LAYER ME2 ;
 ANTENNADIFFAREA                          0.160 LAYER ME3 ;
 ANTENNADIFFAREA                          0.160 LAYER ME4 ;
 ANTENNAMAXAREACAR                       59.337 LAYER ME2 ;
 ANTENNAMAXAREACAR                       66.744 LAYER ME3 ;
 ANTENNAMAXAREACAR                       74.152 LAYER ME4 ;
END CK
PIN A4
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 1338.000 0.000 1338.800 1.000 ;
  LAYER ME3 ;
  RECT 1338.000 0.000 1338.800 1.000 ;
  LAYER ME2 ;
  RECT 1338.000 0.000 1338.800 1.000 ;
  LAYER ME1 ;
  RECT 1338.000 0.000 1338.800 1.000 ;
 END
 ANTENNAPARTIALMETALAREA                  2.212 LAYER ME2 ;
 ANTENNAGATEAREA                          0.180 LAYER ME2 ;
 ANTENNAGATEAREA                          0.180 LAYER ME3 ;
 ANTENNAGATEAREA                          0.180 LAYER ME4 ;
 ANTENNADIFFAREA                          0.160 LAYER ME2 ;
 ANTENNADIFFAREA                          0.160 LAYER ME3 ;
 ANTENNADIFFAREA                          0.160 LAYER ME4 ;
 ANTENNAMAXAREACAR                       18.181 LAYER ME2 ;
 ANTENNAMAXAREACAR                       22.626 LAYER ME3 ;
 ANTENNAMAXAREACAR                       27.070 LAYER ME4 ;
END A4
PIN A5
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 1335.200 0.000 1336.000 1.000 ;
  LAYER ME3 ;
  RECT 1335.200 0.000 1336.000 1.000 ;
  LAYER ME2 ;
  RECT 1335.200 0.000 1336.000 1.000 ;
  LAYER ME1 ;
  RECT 1335.200 0.000 1336.000 1.000 ;
 END
 ANTENNAPARTIALMETALAREA                  2.406 LAYER ME2 ;
 ANTENNAGATEAREA                          0.180 LAYER ME2 ;
 ANTENNAGATEAREA                          0.180 LAYER ME3 ;
 ANTENNAGATEAREA                          0.180 LAYER ME4 ;
 ANTENNADIFFAREA                          0.160 LAYER ME2 ;
 ANTENNADIFFAREA                          0.160 LAYER ME3 ;
 ANTENNADIFFAREA                          0.160 LAYER ME4 ;
 ANTENNAMAXAREACAR                       19.319 LAYER ME2 ;
 ANTENNAMAXAREACAR                       23.763 LAYER ME3 ;
 ANTENNAMAXAREACAR                       28.208 LAYER ME4 ;
END A5
PIN A6
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 1332.400 0.000 1333.200 1.000 ;
  LAYER ME3 ;
  RECT 1332.400 0.000 1333.200 1.000 ;
  LAYER ME2 ;
  RECT 1332.400 0.000 1333.200 1.000 ;
  LAYER ME1 ;
  RECT 1332.400 0.000 1333.200 1.000 ;
 END
 ANTENNAPARTIALMETALAREA                  2.394 LAYER ME2 ;
 ANTENNAGATEAREA                          0.180 LAYER ME2 ;
 ANTENNAGATEAREA                          0.180 LAYER ME3 ;
 ANTENNAGATEAREA                          0.180 LAYER ME4 ;
 ANTENNADIFFAREA                          0.160 LAYER ME2 ;
 ANTENNADIFFAREA                          0.160 LAYER ME3 ;
 ANTENNADIFFAREA                          0.160 LAYER ME4 ;
 ANTENNAMAXAREACAR                       19.156 LAYER ME2 ;
 ANTENNAMAXAREACAR                       23.600 LAYER ME3 ;
 ANTENNAMAXAREACAR                       28.044 LAYER ME4 ;
END A6
PIN A7
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 1330.000 0.000 1330.800 1.000 ;
  LAYER ME3 ;
  RECT 1330.000 0.000 1330.800 1.000 ;
  LAYER ME2 ;
  RECT 1330.000 0.000 1330.800 1.000 ;
  LAYER ME1 ;
  RECT 1330.000 0.000 1330.800 1.000 ;
 END
 ANTENNAPARTIALMETALAREA                  2.378 LAYER ME2 ;
 ANTENNAGATEAREA                          0.180 LAYER ME2 ;
 ANTENNAGATEAREA                          0.180 LAYER ME3 ;
 ANTENNAGATEAREA                          0.180 LAYER ME4 ;
 ANTENNADIFFAREA                          0.160 LAYER ME2 ;
 ANTENNADIFFAREA                          0.160 LAYER ME3 ;
 ANTENNADIFFAREA                          0.160 LAYER ME4 ;
 ANTENNAMAXAREACAR                       19.067 LAYER ME2 ;
 ANTENNAMAXAREACAR                       23.511 LAYER ME3 ;
 ANTENNAMAXAREACAR                       27.956 LAYER ME4 ;
END A7
PIN A8
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 1328.400 0.000 1329.200 1.000 ;
  LAYER ME3 ;
  RECT 1328.400 0.000 1329.200 1.000 ;
  LAYER ME2 ;
  RECT 1328.400 0.000 1329.200 1.000 ;
  LAYER ME1 ;
  RECT 1328.400 0.000 1329.200 1.000 ;
 END
 ANTENNAPARTIALMETALAREA                  2.394 LAYER ME2 ;
 ANTENNAGATEAREA                          0.180 LAYER ME2 ;
 ANTENNAGATEAREA                          0.180 LAYER ME3 ;
 ANTENNAGATEAREA                          0.180 LAYER ME4 ;
 ANTENNADIFFAREA                          0.160 LAYER ME2 ;
 ANTENNADIFFAREA                          0.160 LAYER ME3 ;
 ANTENNADIFFAREA                          0.160 LAYER ME4 ;
 ANTENNAMAXAREACAR                       19.156 LAYER ME2 ;
 ANTENNAMAXAREACAR                       23.600 LAYER ME3 ;
 ANTENNAMAXAREACAR                       28.044 LAYER ME4 ;
END A8
PIN A9
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 1326.000 0.000 1326.800 1.000 ;
  LAYER ME3 ;
  RECT 1326.000 0.000 1326.800 1.000 ;
  LAYER ME2 ;
  RECT 1326.000 0.000 1326.800 1.000 ;
  LAYER ME1 ;
  RECT 1326.000 0.000 1326.800 1.000 ;
 END
 ANTENNAPARTIALMETALAREA                  2.378 LAYER ME2 ;
 ANTENNAGATEAREA                          0.180 LAYER ME2 ;
 ANTENNAGATEAREA                          0.180 LAYER ME3 ;
 ANTENNAGATEAREA                          0.180 LAYER ME4 ;
 ANTENNADIFFAREA                          0.160 LAYER ME2 ;
 ANTENNADIFFAREA                          0.160 LAYER ME3 ;
 ANTENNADIFFAREA                          0.160 LAYER ME4 ;
 ANTENNAMAXAREACAR                       19.067 LAYER ME2 ;
 ANTENNAMAXAREACAR                       23.511 LAYER ME3 ;
 ANTENNAMAXAREACAR                       27.956 LAYER ME4 ;
END A9
PIN A10
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 1324.400 0.000 1325.200 1.000 ;
  LAYER ME3 ;
  RECT 1324.400 0.000 1325.200 1.000 ;
  LAYER ME2 ;
  RECT 1324.400 0.000 1325.200 1.000 ;
  LAYER ME1 ;
  RECT 1324.400 0.000 1325.200 1.000 ;
 END
 ANTENNAPARTIALMETALAREA                  2.394 LAYER ME2 ;
 ANTENNAGATEAREA                          0.180 LAYER ME2 ;
 ANTENNAGATEAREA                          0.180 LAYER ME3 ;
 ANTENNAGATEAREA                          0.180 LAYER ME4 ;
 ANTENNADIFFAREA                          0.160 LAYER ME2 ;
 ANTENNADIFFAREA                          0.160 LAYER ME3 ;
 ANTENNADIFFAREA                          0.160 LAYER ME4 ;
 ANTENNAMAXAREACAR                       19.156 LAYER ME2 ;
 ANTENNAMAXAREACAR                       23.600 LAYER ME3 ;
 ANTENNAMAXAREACAR                       28.044 LAYER ME4 ;
END A10
PIN A11
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 1322.000 0.000 1322.800 1.000 ;
  LAYER ME3 ;
  RECT 1322.000 0.000 1322.800 1.000 ;
  LAYER ME2 ;
  RECT 1322.000 0.000 1322.800 1.000 ;
  LAYER ME1 ;
  RECT 1322.000 0.000 1322.800 1.000 ;
 END
 ANTENNAPARTIALMETALAREA                  2.378 LAYER ME2 ;
 ANTENNAGATEAREA                          0.180 LAYER ME2 ;
 ANTENNAGATEAREA                          0.180 LAYER ME3 ;
 ANTENNAGATEAREA                          0.180 LAYER ME4 ;
 ANTENNADIFFAREA                          0.160 LAYER ME2 ;
 ANTENNADIFFAREA                          0.160 LAYER ME3 ;
 ANTENNADIFFAREA                          0.160 LAYER ME4 ;
 ANTENNAMAXAREACAR                       19.067 LAYER ME2 ;
 ANTENNAMAXAREACAR                       23.511 LAYER ME3 ;
 ANTENNAMAXAREACAR                       27.956 LAYER ME4 ;
END A11
PIN A12
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 1320.400 0.000 1321.200 1.000 ;
  LAYER ME3 ;
  RECT 1320.400 0.000 1321.200 1.000 ;
  LAYER ME2 ;
  RECT 1320.400 0.000 1321.200 1.000 ;
  LAYER ME1 ;
  RECT 1320.400 0.000 1321.200 1.000 ;
 END
 ANTENNAPARTIALMETALAREA                  2.394 LAYER ME2 ;
 ANTENNAGATEAREA                          0.180 LAYER ME2 ;
 ANTENNAGATEAREA                          0.180 LAYER ME3 ;
 ANTENNAGATEAREA                          0.180 LAYER ME4 ;
 ANTENNADIFFAREA                          0.160 LAYER ME2 ;
 ANTENNADIFFAREA                          0.160 LAYER ME3 ;
 ANTENNADIFFAREA                          0.160 LAYER ME4 ;
 ANTENNAMAXAREACAR                       19.156 LAYER ME2 ;
 ANTENNAMAXAREACAR                       23.600 LAYER ME3 ;
 ANTENNAMAXAREACAR                       28.044 LAYER ME4 ;
END A12
PIN DO63
  DIRECTION OUTPUT ;
 PORT
  LAYER ME4 ;
  RECT 1311.200 0.000 1312.000 1.000 ;
  LAYER ME3 ;
  RECT 1311.200 0.000 1312.000 1.000 ;
  LAYER ME2 ;
  RECT 1311.200 0.000 1312.000 1.000 ;
  LAYER ME1 ;
  RECT 1311.200 0.000 1312.000 1.000 ;
 END
 ANTENNAPARTIALMETALAREA                  4.148 LAYER ME2 ;
 ANTENNADIFFAREA                          5.472 LAYER ME2 ;
 ANTENNADIFFAREA                          5.472 LAYER ME3 ;
 ANTENNADIFFAREA                          5.472 LAYER ME4 ;
END DO63
PIN DI63
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 1296.400 0.000 1297.200 1.000 ;
  LAYER ME3 ;
  RECT 1296.400 0.000 1297.200 1.000 ;
  LAYER ME2 ;
  RECT 1296.400 0.000 1297.200 1.000 ;
  LAYER ME1 ;
  RECT 1296.400 0.000 1297.200 1.000 ;
 END
 ANTENNAPARTIALMETALAREA                  3.142 LAYER ME2 ;
 ANTENNAGATEAREA                          0.086 LAYER ME2 ;
 ANTENNAGATEAREA                          0.086 LAYER ME3 ;
 ANTENNAGATEAREA                          0.086 LAYER ME4 ;
 ANTENNADIFFAREA                          0.160 LAYER ME2 ;
 ANTENNADIFFAREA                          0.160 LAYER ME3 ;
 ANTENNADIFFAREA                          0.160 LAYER ME4 ;
 ANTENNAMAXAREACAR                       48.708 LAYER ME2 ;
 ANTENNAMAXAREACAR                       57.968 LAYER ME3 ;
 ANTENNAMAXAREACAR                       67.227 LAYER ME4 ;
END DI63
PIN DO62
  DIRECTION OUTPUT ;
 PORT
  LAYER ME4 ;
  RECT 1291.200 0.000 1292.000 1.000 ;
  LAYER ME3 ;
  RECT 1291.200 0.000 1292.000 1.000 ;
  LAYER ME2 ;
  RECT 1291.200 0.000 1292.000 1.000 ;
  LAYER ME1 ;
  RECT 1291.200 0.000 1292.000 1.000 ;
 END
 ANTENNAPARTIALMETALAREA                  4.164 LAYER ME2 ;
 ANTENNADIFFAREA                          5.472 LAYER ME2 ;
 ANTENNADIFFAREA                          5.472 LAYER ME3 ;
 ANTENNADIFFAREA                          5.472 LAYER ME4 ;
END DO62
PIN DI62
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 1276.800 0.000 1277.600 1.000 ;
  LAYER ME3 ;
  RECT 1276.800 0.000 1277.600 1.000 ;
  LAYER ME2 ;
  RECT 1276.800 0.000 1277.600 1.000 ;
  LAYER ME1 ;
  RECT 1276.800 0.000 1277.600 1.000 ;
 END
 ANTENNAPARTIALMETALAREA                  3.138 LAYER ME2 ;
 ANTENNAGATEAREA                          0.086 LAYER ME2 ;
 ANTENNAGATEAREA                          0.086 LAYER ME3 ;
 ANTENNAGATEAREA                          0.086 LAYER ME4 ;
 ANTENNADIFFAREA                          0.160 LAYER ME2 ;
 ANTENNADIFFAREA                          0.160 LAYER ME3 ;
 ANTENNADIFFAREA                          0.160 LAYER ME4 ;
 ANTENNAMAXAREACAR                       48.662 LAYER ME2 ;
 ANTENNAMAXAREACAR                       57.921 LAYER ME3 ;
 ANTENNAMAXAREACAR                       67.181 LAYER ME4 ;
END DI62
PIN DO61
  DIRECTION OUTPUT ;
 PORT
  LAYER ME4 ;
  RECT 1270.400 0.000 1271.200 1.000 ;
  LAYER ME3 ;
  RECT 1270.400 0.000 1271.200 1.000 ;
  LAYER ME2 ;
  RECT 1270.400 0.000 1271.200 1.000 ;
  LAYER ME1 ;
  RECT 1270.400 0.000 1271.200 1.000 ;
 END
 ANTENNAPARTIALMETALAREA                  4.172 LAYER ME2 ;
 ANTENNADIFFAREA                          5.472 LAYER ME2 ;
 ANTENNADIFFAREA                          5.472 LAYER ME3 ;
 ANTENNADIFFAREA                          5.472 LAYER ME4 ;
END DO61
PIN DI61
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 1255.600 0.000 1256.400 1.000 ;
  LAYER ME3 ;
  RECT 1255.600 0.000 1256.400 1.000 ;
  LAYER ME2 ;
  RECT 1255.600 0.000 1256.400 1.000 ;
  LAYER ME1 ;
  RECT 1255.600 0.000 1256.400 1.000 ;
 END
 ANTENNAPARTIALMETALAREA                  3.118 LAYER ME2 ;
 ANTENNAGATEAREA                          0.086 LAYER ME2 ;
 ANTENNAGATEAREA                          0.086 LAYER ME3 ;
 ANTENNAGATEAREA                          0.086 LAYER ME4 ;
 ANTENNADIFFAREA                          0.160 LAYER ME2 ;
 ANTENNADIFFAREA                          0.160 LAYER ME3 ;
 ANTENNADIFFAREA                          0.160 LAYER ME4 ;
 ANTENNAMAXAREACAR                       48.431 LAYER ME2 ;
 ANTENNAMAXAREACAR                       57.690 LAYER ME3 ;
 ANTENNAMAXAREACAR                       66.949 LAYER ME4 ;
END DI61
PIN DO60
  DIRECTION OUTPUT ;
 PORT
  LAYER ME4 ;
  RECT 1250.400 0.000 1251.200 1.000 ;
  LAYER ME3 ;
  RECT 1250.400 0.000 1251.200 1.000 ;
  LAYER ME2 ;
  RECT 1250.400 0.000 1251.200 1.000 ;
  LAYER ME1 ;
  RECT 1250.400 0.000 1251.200 1.000 ;
 END
 ANTENNAPARTIALMETALAREA                  4.140 LAYER ME2 ;
 ANTENNADIFFAREA                          5.472 LAYER ME2 ;
 ANTENNADIFFAREA                          5.472 LAYER ME3 ;
 ANTENNADIFFAREA                          5.472 LAYER ME4 ;
END DO60
PIN DI60
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 1235.600 0.000 1236.400 1.000 ;
  LAYER ME3 ;
  RECT 1235.600 0.000 1236.400 1.000 ;
  LAYER ME2 ;
  RECT 1235.600 0.000 1236.400 1.000 ;
  LAYER ME1 ;
  RECT 1235.600 0.000 1236.400 1.000 ;
 END
 ANTENNAPARTIALMETALAREA                  3.150 LAYER ME2 ;
 ANTENNAGATEAREA                          0.086 LAYER ME2 ;
 ANTENNAGATEAREA                          0.086 LAYER ME3 ;
 ANTENNAGATEAREA                          0.086 LAYER ME4 ;
 ANTENNADIFFAREA                          0.160 LAYER ME2 ;
 ANTENNADIFFAREA                          0.160 LAYER ME3 ;
 ANTENNADIFFAREA                          0.160 LAYER ME4 ;
 ANTENNAMAXAREACAR                       48.801 LAYER ME2 ;
 ANTENNAMAXAREACAR                       58.060 LAYER ME3 ;
 ANTENNAMAXAREACAR                       67.319 LAYER ME4 ;
END DI60
PIN DO59
  DIRECTION OUTPUT ;
 PORT
  LAYER ME4 ;
  RECT 1229.200 0.000 1230.000 1.000 ;
  LAYER ME3 ;
  RECT 1229.200 0.000 1230.000 1.000 ;
  LAYER ME2 ;
  RECT 1229.200 0.000 1230.000 1.000 ;
  LAYER ME1 ;
  RECT 1229.200 0.000 1230.000 1.000 ;
 END
 ANTENNAPARTIALMETALAREA                  4.164 LAYER ME2 ;
 ANTENNADIFFAREA                          5.472 LAYER ME2 ;
 ANTENNADIFFAREA                          5.472 LAYER ME3 ;
 ANTENNADIFFAREA                          5.472 LAYER ME4 ;
END DO59
PIN DI59
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 1214.800 0.000 1215.600 1.000 ;
  LAYER ME3 ;
  RECT 1214.800 0.000 1215.600 1.000 ;
  LAYER ME2 ;
  RECT 1214.800 0.000 1215.600 1.000 ;
  LAYER ME1 ;
  RECT 1214.800 0.000 1215.600 1.000 ;
 END
 ANTENNAPARTIALMETALAREA                  3.138 LAYER ME2 ;
 ANTENNAGATEAREA                          0.086 LAYER ME2 ;
 ANTENNAGATEAREA                          0.086 LAYER ME3 ;
 ANTENNAGATEAREA                          0.086 LAYER ME4 ;
 ANTENNADIFFAREA                          0.160 LAYER ME2 ;
 ANTENNADIFFAREA                          0.160 LAYER ME3 ;
 ANTENNADIFFAREA                          0.160 LAYER ME4 ;
 ANTENNAMAXAREACAR                       48.662 LAYER ME2 ;
 ANTENNAMAXAREACAR                       57.921 LAYER ME3 ;
 ANTENNAMAXAREACAR                       67.181 LAYER ME4 ;
END DI59
PIN DO58
  DIRECTION OUTPUT ;
 PORT
  LAYER ME4 ;
  RECT 1209.600 0.000 1210.400 1.000 ;
  LAYER ME3 ;
  RECT 1209.600 0.000 1210.400 1.000 ;
  LAYER ME2 ;
  RECT 1209.600 0.000 1210.400 1.000 ;
  LAYER ME1 ;
  RECT 1209.600 0.000 1210.400 1.000 ;
 END
 ANTENNAPARTIALMETALAREA                  4.164 LAYER ME2 ;
 ANTENNADIFFAREA                          5.472 LAYER ME2 ;
 ANTENNADIFFAREA                          5.472 LAYER ME3 ;
 ANTENNADIFFAREA                          5.472 LAYER ME4 ;
END DO58
PIN DI58
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 1194.800 0.000 1195.600 1.000 ;
  LAYER ME3 ;
  RECT 1194.800 0.000 1195.600 1.000 ;
  LAYER ME2 ;
  RECT 1194.800 0.000 1195.600 1.000 ;
  LAYER ME1 ;
  RECT 1194.800 0.000 1195.600 1.000 ;
 END
 ANTENNAPARTIALMETALAREA                  3.126 LAYER ME2 ;
 ANTENNAGATEAREA                          0.086 LAYER ME2 ;
 ANTENNAGATEAREA                          0.086 LAYER ME3 ;
 ANTENNAGATEAREA                          0.086 LAYER ME4 ;
 ANTENNADIFFAREA                          0.160 LAYER ME2 ;
 ANTENNADIFFAREA                          0.160 LAYER ME3 ;
 ANTENNADIFFAREA                          0.160 LAYER ME4 ;
 ANTENNAMAXAREACAR                       48.523 LAYER ME2 ;
 ANTENNAMAXAREACAR                       57.782 LAYER ME3 ;
 ANTENNAMAXAREACAR                       67.042 LAYER ME4 ;
END DI58
PIN DO57
  DIRECTION OUTPUT ;
 PORT
  LAYER ME4 ;
  RECT 1188.400 0.000 1189.200 1.000 ;
  LAYER ME3 ;
  RECT 1188.400 0.000 1189.200 1.000 ;
  LAYER ME2 ;
  RECT 1188.400 0.000 1189.200 1.000 ;
  LAYER ME1 ;
  RECT 1188.400 0.000 1189.200 1.000 ;
 END
 ANTENNAPARTIALMETALAREA                  4.140 LAYER ME2 ;
 ANTENNADIFFAREA                          5.472 LAYER ME2 ;
 ANTENNADIFFAREA                          5.472 LAYER ME3 ;
 ANTENNADIFFAREA                          5.472 LAYER ME4 ;
END DO57
PIN DI57
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 1173.600 0.000 1174.400 1.000 ;
  LAYER ME3 ;
  RECT 1173.600 0.000 1174.400 1.000 ;
  LAYER ME2 ;
  RECT 1173.600 0.000 1174.400 1.000 ;
  LAYER ME1 ;
  RECT 1173.600 0.000 1174.400 1.000 ;
 END
 ANTENNAPARTIALMETALAREA                  3.150 LAYER ME2 ;
 ANTENNAGATEAREA                          0.086 LAYER ME2 ;
 ANTENNAGATEAREA                          0.086 LAYER ME3 ;
 ANTENNAGATEAREA                          0.086 LAYER ME4 ;
 ANTENNADIFFAREA                          0.160 LAYER ME2 ;
 ANTENNADIFFAREA                          0.160 LAYER ME3 ;
 ANTENNADIFFAREA                          0.160 LAYER ME4 ;
 ANTENNAMAXAREACAR                       48.801 LAYER ME2 ;
 ANTENNAMAXAREACAR                       58.060 LAYER ME3 ;
 ANTENNAMAXAREACAR                       67.319 LAYER ME4 ;
END DI57
PIN DO56
  DIRECTION OUTPUT ;
 PORT
  LAYER ME4 ;
  RECT 1168.400 0.000 1169.200 1.000 ;
  LAYER ME3 ;
  RECT 1168.400 0.000 1169.200 1.000 ;
  LAYER ME2 ;
  RECT 1168.400 0.000 1169.200 1.000 ;
  LAYER ME1 ;
  RECT 1168.400 0.000 1169.200 1.000 ;
 END
 ANTENNAPARTIALMETALAREA                  4.172 LAYER ME2 ;
 ANTENNADIFFAREA                          5.472 LAYER ME2 ;
 ANTENNADIFFAREA                          5.472 LAYER ME3 ;
 ANTENNADIFFAREA                          5.472 LAYER ME4 ;
END DO56
PIN WEB7
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 1155.600 0.000 1156.400 1.000 ;
  LAYER ME3 ;
  RECT 1155.600 0.000 1156.400 1.000 ;
  LAYER ME2 ;
  RECT 1155.600 0.000 1156.400 1.000 ;
  LAYER ME1 ;
  RECT 1155.600 0.000 1156.400 1.000 ;
 END
 ANTENNAPARTIALMETALAREA                  2.840 LAYER ME2 ;
 ANTENNAGATEAREA                          0.072 LAYER ME2 ;
 ANTENNAGATEAREA                          0.072 LAYER ME3 ;
 ANTENNAGATEAREA                          0.072 LAYER ME4 ;
 ANTENNADIFFAREA                          0.160 LAYER ME2 ;
 ANTENNADIFFAREA                          0.160 LAYER ME3 ;
 ANTENNADIFFAREA                          0.160 LAYER ME4 ;
 ANTENNAMAXAREACAR                       54.456 LAYER ME2 ;
 ANTENNAMAXAREACAR                       65.567 LAYER ME3 ;
 ANTENNAMAXAREACAR                       76.678 LAYER ME4 ;
END WEB7
PIN DI56
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 1154.000 0.000 1154.800 1.000 ;
  LAYER ME3 ;
  RECT 1154.000 0.000 1154.800 1.000 ;
  LAYER ME2 ;
  RECT 1154.000 0.000 1154.800 1.000 ;
  LAYER ME1 ;
  RECT 1154.000 0.000 1154.800 1.000 ;
 END
 ANTENNAPARTIALMETALAREA                  3.130 LAYER ME2 ;
 ANTENNAGATEAREA                          0.086 LAYER ME2 ;
 ANTENNAGATEAREA                          0.086 LAYER ME3 ;
 ANTENNAGATEAREA                          0.086 LAYER ME4 ;
 ANTENNADIFFAREA                          0.160 LAYER ME2 ;
 ANTENNADIFFAREA                          0.160 LAYER ME3 ;
 ANTENNADIFFAREA                          0.160 LAYER ME4 ;
 ANTENNAMAXAREACAR                       48.569 LAYER ME2 ;
 ANTENNAMAXAREACAR                       57.829 LAYER ME3 ;
 ANTENNAMAXAREACAR                       67.088 LAYER ME4 ;
END DI56
PIN DO55
  DIRECTION OUTPUT ;
 PORT
  LAYER ME4 ;
  RECT 1147.600 0.000 1148.400 1.000 ;
  LAYER ME3 ;
  RECT 1147.600 0.000 1148.400 1.000 ;
  LAYER ME2 ;
  RECT 1147.600 0.000 1148.400 1.000 ;
  LAYER ME1 ;
  RECT 1147.600 0.000 1148.400 1.000 ;
 END
 ANTENNAPARTIALMETALAREA                  4.164 LAYER ME2 ;
 ANTENNADIFFAREA                          5.472 LAYER ME2 ;
 ANTENNADIFFAREA                          5.472 LAYER ME3 ;
 ANTENNADIFFAREA                          5.472 LAYER ME4 ;
END DO55
PIN DI55
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 1132.800 0.000 1133.600 1.000 ;
  LAYER ME3 ;
  RECT 1132.800 0.000 1133.600 1.000 ;
  LAYER ME2 ;
  RECT 1132.800 0.000 1133.600 1.000 ;
  LAYER ME1 ;
  RECT 1132.800 0.000 1133.600 1.000 ;
 END
 ANTENNAPARTIALMETALAREA                  3.126 LAYER ME2 ;
 ANTENNAGATEAREA                          0.086 LAYER ME2 ;
 ANTENNAGATEAREA                          0.086 LAYER ME3 ;
 ANTENNAGATEAREA                          0.086 LAYER ME4 ;
 ANTENNADIFFAREA                          0.160 LAYER ME2 ;
 ANTENNADIFFAREA                          0.160 LAYER ME3 ;
 ANTENNADIFFAREA                          0.160 LAYER ME4 ;
 ANTENNAMAXAREACAR                       48.523 LAYER ME2 ;
 ANTENNAMAXAREACAR                       57.782 LAYER ME3 ;
 ANTENNAMAXAREACAR                       67.042 LAYER ME4 ;
END DI55
PIN DO54
  DIRECTION OUTPUT ;
 PORT
  LAYER ME4 ;
  RECT 1127.600 0.000 1128.400 1.000 ;
  LAYER ME3 ;
  RECT 1127.600 0.000 1128.400 1.000 ;
  LAYER ME2 ;
  RECT 1127.600 0.000 1128.400 1.000 ;
  LAYER ME1 ;
  RECT 1127.600 0.000 1128.400 1.000 ;
 END
 ANTENNAPARTIALMETALAREA                  4.148 LAYER ME2 ;
 ANTENNADIFFAREA                          5.472 LAYER ME2 ;
 ANTENNADIFFAREA                          5.472 LAYER ME3 ;
 ANTENNADIFFAREA                          5.472 LAYER ME4 ;
END DO54
PIN DI54
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 1113.200 0.000 1114.000 1.000 ;
  LAYER ME3 ;
  RECT 1113.200 0.000 1114.000 1.000 ;
  LAYER ME2 ;
  RECT 1113.200 0.000 1114.000 1.000 ;
  LAYER ME1 ;
  RECT 1113.200 0.000 1114.000 1.000 ;
 END
 ANTENNAPARTIALMETALAREA                  3.154 LAYER ME2 ;
 ANTENNAGATEAREA                          0.086 LAYER ME2 ;
 ANTENNAGATEAREA                          0.086 LAYER ME3 ;
 ANTENNAGATEAREA                          0.086 LAYER ME4 ;
 ANTENNADIFFAREA                          0.160 LAYER ME2 ;
 ANTENNADIFFAREA                          0.160 LAYER ME3 ;
 ANTENNADIFFAREA                          0.160 LAYER ME4 ;
 ANTENNAMAXAREACAR                       48.847 LAYER ME2 ;
 ANTENNAMAXAREACAR                       58.106 LAYER ME3 ;
 ANTENNAMAXAREACAR                       67.366 LAYER ME4 ;
END DI54
PIN DO53
  DIRECTION OUTPUT ;
 PORT
  LAYER ME4 ;
  RECT 1106.400 0.000 1107.200 1.000 ;
  LAYER ME3 ;
  RECT 1106.400 0.000 1107.200 1.000 ;
  LAYER ME2 ;
  RECT 1106.400 0.000 1107.200 1.000 ;
  LAYER ME1 ;
  RECT 1106.400 0.000 1107.200 1.000 ;
 END
 ANTENNAPARTIALMETALAREA                  4.172 LAYER ME2 ;
 ANTENNADIFFAREA                          5.472 LAYER ME2 ;
 ANTENNADIFFAREA                          5.472 LAYER ME3 ;
 ANTENNADIFFAREA                          5.472 LAYER ME4 ;
END DO53
PIN DI53
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 1092.000 0.000 1092.800 1.000 ;
  LAYER ME3 ;
  RECT 1092.000 0.000 1092.800 1.000 ;
  LAYER ME2 ;
  RECT 1092.000 0.000 1092.800 1.000 ;
  LAYER ME1 ;
  RECT 1092.000 0.000 1092.800 1.000 ;
 END
 ANTENNAPARTIALMETALAREA                  3.130 LAYER ME2 ;
 ANTENNAGATEAREA                          0.086 LAYER ME2 ;
 ANTENNAGATEAREA                          0.086 LAYER ME3 ;
 ANTENNAGATEAREA                          0.086 LAYER ME4 ;
 ANTENNADIFFAREA                          0.160 LAYER ME2 ;
 ANTENNADIFFAREA                          0.160 LAYER ME3 ;
 ANTENNADIFFAREA                          0.160 LAYER ME4 ;
 ANTENNAMAXAREACAR                       48.569 LAYER ME2 ;
 ANTENNAMAXAREACAR                       57.829 LAYER ME3 ;
 ANTENNAMAXAREACAR                       67.088 LAYER ME4 ;
END DI53
PIN DO52
  DIRECTION OUTPUT ;
 PORT
  LAYER ME4 ;
  RECT 1086.800 0.000 1087.600 1.000 ;
  LAYER ME3 ;
  RECT 1086.800 0.000 1087.600 1.000 ;
  LAYER ME2 ;
  RECT 1086.800 0.000 1087.600 1.000 ;
  LAYER ME1 ;
  RECT 1086.800 0.000 1087.600 1.000 ;
 END
 ANTENNAPARTIALMETALAREA                  4.156 LAYER ME2 ;
 ANTENNADIFFAREA                          5.472 LAYER ME2 ;
 ANTENNADIFFAREA                          5.472 LAYER ME3 ;
 ANTENNADIFFAREA                          5.472 LAYER ME4 ;
END DO52
PIN DI52
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 1072.000 0.000 1072.800 1.000 ;
  LAYER ME3 ;
  RECT 1072.000 0.000 1072.800 1.000 ;
  LAYER ME2 ;
  RECT 1072.000 0.000 1072.800 1.000 ;
  LAYER ME1 ;
  RECT 1072.000 0.000 1072.800 1.000 ;
 END
 ANTENNAPARTIALMETALAREA                  3.134 LAYER ME2 ;
 ANTENNAGATEAREA                          0.086 LAYER ME2 ;
 ANTENNAGATEAREA                          0.086 LAYER ME3 ;
 ANTENNAGATEAREA                          0.086 LAYER ME4 ;
 ANTENNADIFFAREA                          0.160 LAYER ME2 ;
 ANTENNADIFFAREA                          0.160 LAYER ME3 ;
 ANTENNADIFFAREA                          0.160 LAYER ME4 ;
 ANTENNAMAXAREACAR                       48.616 LAYER ME2 ;
 ANTENNAMAXAREACAR                       57.875 LAYER ME3 ;
 ANTENNAMAXAREACAR                       67.134 LAYER ME4 ;
END DI52
PIN DO51
  DIRECTION OUTPUT ;
 PORT
  LAYER ME4 ;
  RECT 1065.600 0.000 1066.400 1.000 ;
  LAYER ME3 ;
  RECT 1065.600 0.000 1066.400 1.000 ;
  LAYER ME2 ;
  RECT 1065.600 0.000 1066.400 1.000 ;
  LAYER ME1 ;
  RECT 1065.600 0.000 1066.400 1.000 ;
 END
 ANTENNAPARTIALMETALAREA                  4.148 LAYER ME2 ;
 ANTENNADIFFAREA                          5.472 LAYER ME2 ;
 ANTENNADIFFAREA                          5.472 LAYER ME3 ;
 ANTENNADIFFAREA                          5.472 LAYER ME4 ;
END DO51
PIN DI51
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 1051.200 0.000 1052.000 1.000 ;
  LAYER ME3 ;
  RECT 1051.200 0.000 1052.000 1.000 ;
  LAYER ME2 ;
  RECT 1051.200 0.000 1052.000 1.000 ;
  LAYER ME1 ;
  RECT 1051.200 0.000 1052.000 1.000 ;
 END
 ANTENNAPARTIALMETALAREA                  3.154 LAYER ME2 ;
 ANTENNAGATEAREA                          0.086 LAYER ME2 ;
 ANTENNAGATEAREA                          0.086 LAYER ME3 ;
 ANTENNAGATEAREA                          0.086 LAYER ME4 ;
 ANTENNADIFFAREA                          0.160 LAYER ME2 ;
 ANTENNADIFFAREA                          0.160 LAYER ME3 ;
 ANTENNADIFFAREA                          0.160 LAYER ME4 ;
 ANTENNAMAXAREACAR                       48.847 LAYER ME2 ;
 ANTENNAMAXAREACAR                       58.106 LAYER ME3 ;
 ANTENNAMAXAREACAR                       67.366 LAYER ME4 ;
END DI51
PIN DO50
  DIRECTION OUTPUT ;
 PORT
  LAYER ME4 ;
  RECT 1045.600 0.000 1046.400 1.000 ;
  LAYER ME3 ;
  RECT 1045.600 0.000 1046.400 1.000 ;
  LAYER ME2 ;
  RECT 1045.600 0.000 1046.400 1.000 ;
  LAYER ME1 ;
  RECT 1045.600 0.000 1046.400 1.000 ;
 END
 ANTENNAPARTIALMETALAREA                  4.180 LAYER ME2 ;
 ANTENNADIFFAREA                          5.472 LAYER ME2 ;
 ANTENNADIFFAREA                          5.472 LAYER ME3 ;
 ANTENNADIFFAREA                          5.472 LAYER ME4 ;
END DO50
PIN DI50
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 1031.200 0.000 1032.000 1.000 ;
  LAYER ME3 ;
  RECT 1031.200 0.000 1032.000 1.000 ;
  LAYER ME2 ;
  RECT 1031.200 0.000 1032.000 1.000 ;
  LAYER ME1 ;
  RECT 1031.200 0.000 1032.000 1.000 ;
 END
 ANTENNAPARTIALMETALAREA                  3.122 LAYER ME2 ;
 ANTENNAGATEAREA                          0.086 LAYER ME2 ;
 ANTENNAGATEAREA                          0.086 LAYER ME3 ;
 ANTENNAGATEAREA                          0.086 LAYER ME4 ;
 ANTENNADIFFAREA                          0.160 LAYER ME2 ;
 ANTENNADIFFAREA                          0.160 LAYER ME3 ;
 ANTENNADIFFAREA                          0.160 LAYER ME4 ;
 ANTENNAMAXAREACAR                       48.477 LAYER ME2 ;
 ANTENNAMAXAREACAR                       57.736 LAYER ME3 ;
 ANTENNAMAXAREACAR                       66.995 LAYER ME4 ;
END DI50
PIN DO49
  DIRECTION OUTPUT ;
 PORT
  LAYER ME4 ;
  RECT 1024.800 0.000 1025.600 1.000 ;
  LAYER ME3 ;
  RECT 1024.800 0.000 1025.600 1.000 ;
  LAYER ME2 ;
  RECT 1024.800 0.000 1025.600 1.000 ;
  LAYER ME1 ;
  RECT 1024.800 0.000 1025.600 1.000 ;
 END
 ANTENNAPARTIALMETALAREA                  4.156 LAYER ME2 ;
 ANTENNADIFFAREA                          5.472 LAYER ME2 ;
 ANTENNADIFFAREA                          5.472 LAYER ME3 ;
 ANTENNADIFFAREA                          5.472 LAYER ME4 ;
END DO49
PIN DI49
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 1010.000 0.000 1010.800 1.000 ;
  LAYER ME3 ;
  RECT 1010.000 0.000 1010.800 1.000 ;
  LAYER ME2 ;
  RECT 1010.000 0.000 1010.800 1.000 ;
  LAYER ME1 ;
  RECT 1010.000 0.000 1010.800 1.000 ;
 END
 ANTENNAPARTIALMETALAREA                  3.134 LAYER ME2 ;
 ANTENNAGATEAREA                          0.086 LAYER ME2 ;
 ANTENNAGATEAREA                          0.086 LAYER ME3 ;
 ANTENNAGATEAREA                          0.086 LAYER ME4 ;
 ANTENNADIFFAREA                          0.160 LAYER ME2 ;
 ANTENNADIFFAREA                          0.160 LAYER ME3 ;
 ANTENNADIFFAREA                          0.160 LAYER ME4 ;
 ANTENNAMAXAREACAR                       48.616 LAYER ME2 ;
 ANTENNAMAXAREACAR                       57.875 LAYER ME3 ;
 ANTENNAMAXAREACAR                       67.134 LAYER ME4 ;
END DI49
PIN DO48
  DIRECTION OUTPUT ;
 PORT
  LAYER ME4 ;
  RECT 1004.800 0.000 1005.600 1.000 ;
  LAYER ME3 ;
  RECT 1004.800 0.000 1005.600 1.000 ;
  LAYER ME2 ;
  RECT 1004.800 0.000 1005.600 1.000 ;
  LAYER ME1 ;
  RECT 1004.800 0.000 1005.600 1.000 ;
 END
 ANTENNAPARTIALMETALAREA                  4.156 LAYER ME2 ;
 ANTENNADIFFAREA                          5.472 LAYER ME2 ;
 ANTENNADIFFAREA                          5.472 LAYER ME3 ;
 ANTENNADIFFAREA                          5.472 LAYER ME4 ;
END DO48
PIN WEB6
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 992.000 0.000 992.800 1.000 ;
  LAYER ME3 ;
  RECT 992.000 0.000 992.800 1.000 ;
  LAYER ME2 ;
  RECT 992.000 0.000 992.800 1.000 ;
  LAYER ME1 ;
  RECT 992.000 0.000 992.800 1.000 ;
 END
 ANTENNAPARTIALMETALAREA                  2.836 LAYER ME2 ;
 ANTENNAGATEAREA                          0.072 LAYER ME2 ;
 ANTENNAGATEAREA                          0.072 LAYER ME3 ;
 ANTENNAGATEAREA                          0.072 LAYER ME4 ;
 ANTENNADIFFAREA                          0.160 LAYER ME2 ;
 ANTENNADIFFAREA                          0.160 LAYER ME3 ;
 ANTENNADIFFAREA                          0.160 LAYER ME4 ;
 ANTENNAMAXAREACAR                       54.400 LAYER ME2 ;
 ANTENNAMAXAREACAR                       65.511 LAYER ME3 ;
 ANTENNAMAXAREACAR                       76.622 LAYER ME4 ;
END WEB6
PIN DI48
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 990.400 0.000 991.200 1.000 ;
  LAYER ME3 ;
  RECT 990.400 0.000 991.200 1.000 ;
  LAYER ME2 ;
  RECT 990.400 0.000 991.200 1.000 ;
  LAYER ME1 ;
  RECT 990.400 0.000 991.200 1.000 ;
 END
 ANTENNAPARTIALMETALAREA                  3.146 LAYER ME2 ;
 ANTENNAGATEAREA                          0.086 LAYER ME2 ;
 ANTENNAGATEAREA                          0.086 LAYER ME3 ;
 ANTENNAGATEAREA                          0.086 LAYER ME4 ;
 ANTENNADIFFAREA                          0.160 LAYER ME2 ;
 ANTENNADIFFAREA                          0.160 LAYER ME3 ;
 ANTENNADIFFAREA                          0.160 LAYER ME4 ;
 ANTENNAMAXAREACAR                       48.755 LAYER ME2 ;
 ANTENNAMAXAREACAR                       58.014 LAYER ME3 ;
 ANTENNAMAXAREACAR                       67.273 LAYER ME4 ;
END DI48
PIN DO47
  DIRECTION OUTPUT ;
 PORT
  LAYER ME4 ;
  RECT 983.600 0.000 984.400 1.000 ;
  LAYER ME3 ;
  RECT 983.600 0.000 984.400 1.000 ;
  LAYER ME2 ;
  RECT 983.600 0.000 984.400 1.000 ;
  LAYER ME1 ;
  RECT 983.600 0.000 984.400 1.000 ;
 END
 ANTENNAPARTIALMETALAREA                  4.180 LAYER ME2 ;
 ANTENNADIFFAREA                          5.472 LAYER ME2 ;
 ANTENNADIFFAREA                          5.472 LAYER ME3 ;
 ANTENNADIFFAREA                          5.472 LAYER ME4 ;
END DO47
PIN DI47
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 969.200 0.000 970.000 1.000 ;
  LAYER ME3 ;
  RECT 969.200 0.000 970.000 1.000 ;
  LAYER ME2 ;
  RECT 969.200 0.000 970.000 1.000 ;
  LAYER ME1 ;
  RECT 969.200 0.000 970.000 1.000 ;
 END
 ANTENNAPARTIALMETALAREA                  3.122 LAYER ME2 ;
 ANTENNAGATEAREA                          0.086 LAYER ME2 ;
 ANTENNAGATEAREA                          0.086 LAYER ME3 ;
 ANTENNAGATEAREA                          0.086 LAYER ME4 ;
 ANTENNADIFFAREA                          0.160 LAYER ME2 ;
 ANTENNADIFFAREA                          0.160 LAYER ME3 ;
 ANTENNADIFFAREA                          0.160 LAYER ME4 ;
 ANTENNAMAXAREACAR                       48.477 LAYER ME2 ;
 ANTENNAMAXAREACAR                       57.736 LAYER ME3 ;
 ANTENNAMAXAREACAR                       66.995 LAYER ME4 ;
END DI47
PIN DO46
  DIRECTION OUTPUT ;
 PORT
  LAYER ME4 ;
  RECT 964.000 0.000 964.800 1.000 ;
  LAYER ME3 ;
  RECT 964.000 0.000 964.800 1.000 ;
  LAYER ME2 ;
  RECT 964.000 0.000 964.800 1.000 ;
  LAYER ME1 ;
  RECT 964.000 0.000 964.800 1.000 ;
 END
 ANTENNAPARTIALMETALAREA                  4.148 LAYER ME2 ;
 ANTENNADIFFAREA                          5.472 LAYER ME2 ;
 ANTENNADIFFAREA                          5.472 LAYER ME3 ;
 ANTENNADIFFAREA                          5.472 LAYER ME4 ;
END DO46
PIN DI46
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 949.200 0.000 950.000 1.000 ;
  LAYER ME3 ;
  RECT 949.200 0.000 950.000 1.000 ;
  LAYER ME2 ;
  RECT 949.200 0.000 950.000 1.000 ;
  LAYER ME1 ;
  RECT 949.200 0.000 950.000 1.000 ;
 END
 ANTENNAPARTIALMETALAREA                  3.142 LAYER ME2 ;
 ANTENNAGATEAREA                          0.086 LAYER ME2 ;
 ANTENNAGATEAREA                          0.086 LAYER ME3 ;
 ANTENNAGATEAREA                          0.086 LAYER ME4 ;
 ANTENNADIFFAREA                          0.160 LAYER ME2 ;
 ANTENNADIFFAREA                          0.160 LAYER ME3 ;
 ANTENNADIFFAREA                          0.160 LAYER ME4 ;
 ANTENNAMAXAREACAR                       48.708 LAYER ME2 ;
 ANTENNAMAXAREACAR                       57.968 LAYER ME3 ;
 ANTENNAMAXAREACAR                       67.227 LAYER ME4 ;
END DI46
PIN DO45
  DIRECTION OUTPUT ;
 PORT
  LAYER ME4 ;
  RECT 942.800 0.000 943.600 1.000 ;
  LAYER ME3 ;
  RECT 942.800 0.000 943.600 1.000 ;
  LAYER ME2 ;
  RECT 942.800 0.000 943.600 1.000 ;
  LAYER ME1 ;
  RECT 942.800 0.000 943.600 1.000 ;
 END
 ANTENNAPARTIALMETALAREA                  4.156 LAYER ME2 ;
 ANTENNADIFFAREA                          5.472 LAYER ME2 ;
 ANTENNADIFFAREA                          5.472 LAYER ME3 ;
 ANTENNADIFFAREA                          5.472 LAYER ME4 ;
END DO45
PIN DI45
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 928.400 0.000 929.200 1.000 ;
  LAYER ME3 ;
  RECT 928.400 0.000 929.200 1.000 ;
  LAYER ME2 ;
  RECT 928.400 0.000 929.200 1.000 ;
  LAYER ME1 ;
  RECT 928.400 0.000 929.200 1.000 ;
 END
 ANTENNAPARTIALMETALAREA                  3.146 LAYER ME2 ;
 ANTENNAGATEAREA                          0.086 LAYER ME2 ;
 ANTENNAGATEAREA                          0.086 LAYER ME3 ;
 ANTENNAGATEAREA                          0.086 LAYER ME4 ;
 ANTENNADIFFAREA                          0.160 LAYER ME2 ;
 ANTENNADIFFAREA                          0.160 LAYER ME3 ;
 ANTENNADIFFAREA                          0.160 LAYER ME4 ;
 ANTENNAMAXAREACAR                       48.755 LAYER ME2 ;
 ANTENNAMAXAREACAR                       58.014 LAYER ME3 ;
 ANTENNAMAXAREACAR                       67.273 LAYER ME4 ;
END DI45
PIN DO44
  DIRECTION OUTPUT ;
 PORT
  LAYER ME4 ;
  RECT 923.200 0.000 924.000 1.000 ;
  LAYER ME3 ;
  RECT 923.200 0.000 924.000 1.000 ;
  LAYER ME2 ;
  RECT 923.200 0.000 924.000 1.000 ;
  LAYER ME1 ;
  RECT 923.200 0.000 924.000 1.000 ;
 END
 ANTENNAPARTIALMETALAREA                  4.172 LAYER ME2 ;
 ANTENNADIFFAREA                          5.472 LAYER ME2 ;
 ANTENNADIFFAREA                          5.472 LAYER ME3 ;
 ANTENNADIFFAREA                          5.472 LAYER ME4 ;
END DO44
PIN DI44
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 908.400 0.000 909.200 1.000 ;
  LAYER ME3 ;
  RECT 908.400 0.000 909.200 1.000 ;
  LAYER ME2 ;
  RECT 908.400 0.000 909.200 1.000 ;
  LAYER ME1 ;
  RECT 908.400 0.000 909.200 1.000 ;
 END
 ANTENNAPARTIALMETALAREA                  3.118 LAYER ME2 ;
 ANTENNAGATEAREA                          0.086 LAYER ME2 ;
 ANTENNAGATEAREA                          0.086 LAYER ME3 ;
 ANTENNAGATEAREA                          0.086 LAYER ME4 ;
 ANTENNADIFFAREA                          0.160 LAYER ME2 ;
 ANTENNADIFFAREA                          0.160 LAYER ME3 ;
 ANTENNADIFFAREA                          0.160 LAYER ME4 ;
 ANTENNAMAXAREACAR                       48.431 LAYER ME2 ;
 ANTENNAMAXAREACAR                       57.690 LAYER ME3 ;
 ANTENNAMAXAREACAR                       66.949 LAYER ME4 ;
END DI44
PIN DO43
  DIRECTION OUTPUT ;
 PORT
  LAYER ME4 ;
  RECT 902.000 0.000 902.800 1.000 ;
  LAYER ME3 ;
  RECT 902.000 0.000 902.800 1.000 ;
  LAYER ME2 ;
  RECT 902.000 0.000 902.800 1.000 ;
  LAYER ME1 ;
  RECT 902.000 0.000 902.800 1.000 ;
 END
 ANTENNAPARTIALMETALAREA                  4.148 LAYER ME2 ;
 ANTENNADIFFAREA                          5.472 LAYER ME2 ;
 ANTENNADIFFAREA                          5.472 LAYER ME3 ;
 ANTENNADIFFAREA                          5.472 LAYER ME4 ;
END DO43
PIN DI43
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 887.200 0.000 888.000 1.000 ;
  LAYER ME3 ;
  RECT 887.200 0.000 888.000 1.000 ;
  LAYER ME2 ;
  RECT 887.200 0.000 888.000 1.000 ;
  LAYER ME1 ;
  RECT 887.200 0.000 888.000 1.000 ;
 END
 ANTENNAPARTIALMETALAREA                  3.142 LAYER ME2 ;
 ANTENNAGATEAREA                          0.086 LAYER ME2 ;
 ANTENNAGATEAREA                          0.086 LAYER ME3 ;
 ANTENNAGATEAREA                          0.086 LAYER ME4 ;
 ANTENNADIFFAREA                          0.160 LAYER ME2 ;
 ANTENNADIFFAREA                          0.160 LAYER ME3 ;
 ANTENNADIFFAREA                          0.160 LAYER ME4 ;
 ANTENNAMAXAREACAR                       48.708 LAYER ME2 ;
 ANTENNAMAXAREACAR                       57.968 LAYER ME3 ;
 ANTENNAMAXAREACAR                       67.227 LAYER ME4 ;
END DI43
PIN DO42
  DIRECTION OUTPUT ;
 PORT
  LAYER ME4 ;
  RECT 882.000 0.000 882.800 1.000 ;
  LAYER ME3 ;
  RECT 882.000 0.000 882.800 1.000 ;
  LAYER ME2 ;
  RECT 882.000 0.000 882.800 1.000 ;
  LAYER ME1 ;
  RECT 882.000 0.000 882.800 1.000 ;
 END
 ANTENNAPARTIALMETALAREA                  4.164 LAYER ME2 ;
 ANTENNADIFFAREA                          5.472 LAYER ME2 ;
 ANTENNADIFFAREA                          5.472 LAYER ME3 ;
 ANTENNADIFFAREA                          5.472 LAYER ME4 ;
END DO42
PIN DI42
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 867.600 0.000 868.400 1.000 ;
  LAYER ME3 ;
  RECT 867.600 0.000 868.400 1.000 ;
  LAYER ME2 ;
  RECT 867.600 0.000 868.400 1.000 ;
  LAYER ME1 ;
  RECT 867.600 0.000 868.400 1.000 ;
 END
 ANTENNAPARTIALMETALAREA                  3.138 LAYER ME2 ;
 ANTENNAGATEAREA                          0.086 LAYER ME2 ;
 ANTENNAGATEAREA                          0.086 LAYER ME3 ;
 ANTENNAGATEAREA                          0.086 LAYER ME4 ;
 ANTENNADIFFAREA                          0.160 LAYER ME2 ;
 ANTENNADIFFAREA                          0.160 LAYER ME3 ;
 ANTENNADIFFAREA                          0.160 LAYER ME4 ;
 ANTENNAMAXAREACAR                       48.662 LAYER ME2 ;
 ANTENNAMAXAREACAR                       57.921 LAYER ME3 ;
 ANTENNAMAXAREACAR                       67.181 LAYER ME4 ;
END DI42
PIN DO41
  DIRECTION OUTPUT ;
 PORT
  LAYER ME4 ;
  RECT 861.200 0.000 862.000 1.000 ;
  LAYER ME3 ;
  RECT 861.200 0.000 862.000 1.000 ;
  LAYER ME2 ;
  RECT 861.200 0.000 862.000 1.000 ;
  LAYER ME1 ;
  RECT 861.200 0.000 862.000 1.000 ;
 END
 ANTENNAPARTIALMETALAREA                  4.172 LAYER ME2 ;
 ANTENNADIFFAREA                          5.472 LAYER ME2 ;
 ANTENNADIFFAREA                          5.472 LAYER ME3 ;
 ANTENNADIFFAREA                          5.472 LAYER ME4 ;
END DO41
PIN DI41
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 846.400 0.000 847.200 1.000 ;
  LAYER ME3 ;
  RECT 846.400 0.000 847.200 1.000 ;
  LAYER ME2 ;
  RECT 846.400 0.000 847.200 1.000 ;
  LAYER ME1 ;
  RECT 846.400 0.000 847.200 1.000 ;
 END
 ANTENNAPARTIALMETALAREA                  3.118 LAYER ME2 ;
 ANTENNAGATEAREA                          0.086 LAYER ME2 ;
 ANTENNAGATEAREA                          0.086 LAYER ME3 ;
 ANTENNAGATEAREA                          0.086 LAYER ME4 ;
 ANTENNADIFFAREA                          0.160 LAYER ME2 ;
 ANTENNADIFFAREA                          0.160 LAYER ME3 ;
 ANTENNADIFFAREA                          0.160 LAYER ME4 ;
 ANTENNAMAXAREACAR                       48.431 LAYER ME2 ;
 ANTENNAMAXAREACAR                       57.690 LAYER ME3 ;
 ANTENNAMAXAREACAR                       66.949 LAYER ME4 ;
END DI41
PIN DO40
  DIRECTION OUTPUT ;
 PORT
  LAYER ME4 ;
  RECT 841.200 0.000 842.000 1.000 ;
  LAYER ME3 ;
  RECT 841.200 0.000 842.000 1.000 ;
  LAYER ME2 ;
  RECT 841.200 0.000 842.000 1.000 ;
  LAYER ME1 ;
  RECT 841.200 0.000 842.000 1.000 ;
 END
 ANTENNAPARTIALMETALAREA                  4.140 LAYER ME2 ;
 ANTENNADIFFAREA                          5.472 LAYER ME2 ;
 ANTENNADIFFAREA                          5.472 LAYER ME3 ;
 ANTENNADIFFAREA                          5.472 LAYER ME4 ;
END DO40
PIN WEB5
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 828.400 0.000 829.200 1.000 ;
  LAYER ME3 ;
  RECT 828.400 0.000 829.200 1.000 ;
  LAYER ME2 ;
  RECT 828.400 0.000 829.200 1.000 ;
  LAYER ME1 ;
  RECT 828.400 0.000 829.200 1.000 ;
 END
 ANTENNAPARTIALMETALAREA                  2.852 LAYER ME2 ;
 ANTENNAGATEAREA                          0.072 LAYER ME2 ;
 ANTENNAGATEAREA                          0.072 LAYER ME3 ;
 ANTENNAGATEAREA                          0.072 LAYER ME4 ;
 ANTENNADIFFAREA                          0.160 LAYER ME2 ;
 ANTENNADIFFAREA                          0.160 LAYER ME3 ;
 ANTENNADIFFAREA                          0.160 LAYER ME4 ;
 ANTENNAMAXAREACAR                       54.622 LAYER ME2 ;
 ANTENNAMAXAREACAR                       65.733 LAYER ME3 ;
 ANTENNAMAXAREACAR                       76.844 LAYER ME4 ;
END WEB5
PIN DI40
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 826.400 0.000 827.200 1.000 ;
  LAYER ME3 ;
  RECT 826.400 0.000 827.200 1.000 ;
  LAYER ME2 ;
  RECT 826.400 0.000 827.200 1.000 ;
  LAYER ME1 ;
  RECT 826.400 0.000 827.200 1.000 ;
 END
 ANTENNAPARTIALMETALAREA                  3.150 LAYER ME2 ;
 ANTENNAGATEAREA                          0.086 LAYER ME2 ;
 ANTENNAGATEAREA                          0.086 LAYER ME3 ;
 ANTENNAGATEAREA                          0.086 LAYER ME4 ;
 ANTENNADIFFAREA                          0.160 LAYER ME2 ;
 ANTENNADIFFAREA                          0.160 LAYER ME3 ;
 ANTENNADIFFAREA                          0.160 LAYER ME4 ;
 ANTENNAMAXAREACAR                       48.801 LAYER ME2 ;
 ANTENNAMAXAREACAR                       58.060 LAYER ME3 ;
 ANTENNAMAXAREACAR                       67.319 LAYER ME4 ;
END DI40
PIN DO39
  DIRECTION OUTPUT ;
 PORT
  LAYER ME4 ;
  RECT 820.000 0.000 820.800 1.000 ;
  LAYER ME3 ;
  RECT 820.000 0.000 820.800 1.000 ;
  LAYER ME2 ;
  RECT 820.000 0.000 820.800 1.000 ;
  LAYER ME1 ;
  RECT 820.000 0.000 820.800 1.000 ;
 END
 ANTENNAPARTIALMETALAREA                  4.164 LAYER ME2 ;
 ANTENNADIFFAREA                          5.472 LAYER ME2 ;
 ANTENNADIFFAREA                          5.472 LAYER ME3 ;
 ANTENNADIFFAREA                          5.472 LAYER ME4 ;
END DO39
PIN DI39
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 805.600 0.000 806.400 1.000 ;
  LAYER ME3 ;
  RECT 805.600 0.000 806.400 1.000 ;
  LAYER ME2 ;
  RECT 805.600 0.000 806.400 1.000 ;
  LAYER ME1 ;
  RECT 805.600 0.000 806.400 1.000 ;
 END
 ANTENNAPARTIALMETALAREA                  3.138 LAYER ME2 ;
 ANTENNAGATEAREA                          0.086 LAYER ME2 ;
 ANTENNAGATEAREA                          0.086 LAYER ME3 ;
 ANTENNAGATEAREA                          0.086 LAYER ME4 ;
 ANTENNADIFFAREA                          0.160 LAYER ME2 ;
 ANTENNADIFFAREA                          0.160 LAYER ME3 ;
 ANTENNADIFFAREA                          0.160 LAYER ME4 ;
 ANTENNAMAXAREACAR                       48.662 LAYER ME2 ;
 ANTENNAMAXAREACAR                       57.921 LAYER ME3 ;
 ANTENNAMAXAREACAR                       67.181 LAYER ME4 ;
END DI39
PIN DO38
  DIRECTION OUTPUT ;
 PORT
  LAYER ME4 ;
  RECT 800.400 0.000 801.200 1.000 ;
  LAYER ME3 ;
  RECT 800.400 0.000 801.200 1.000 ;
  LAYER ME2 ;
  RECT 800.400 0.000 801.200 1.000 ;
  LAYER ME1 ;
  RECT 800.400 0.000 801.200 1.000 ;
 END
 ANTENNAPARTIALMETALAREA                  4.164 LAYER ME2 ;
 ANTENNADIFFAREA                          5.472 LAYER ME2 ;
 ANTENNADIFFAREA                          5.472 LAYER ME3 ;
 ANTENNADIFFAREA                          5.472 LAYER ME4 ;
END DO38
PIN DI38
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 785.600 0.000 786.400 1.000 ;
  LAYER ME3 ;
  RECT 785.600 0.000 786.400 1.000 ;
  LAYER ME2 ;
  RECT 785.600 0.000 786.400 1.000 ;
  LAYER ME1 ;
  RECT 785.600 0.000 786.400 1.000 ;
 END
 ANTENNAPARTIALMETALAREA                  3.126 LAYER ME2 ;
 ANTENNAGATEAREA                          0.086 LAYER ME2 ;
 ANTENNAGATEAREA                          0.086 LAYER ME3 ;
 ANTENNAGATEAREA                          0.086 LAYER ME4 ;
 ANTENNADIFFAREA                          0.160 LAYER ME2 ;
 ANTENNADIFFAREA                          0.160 LAYER ME3 ;
 ANTENNADIFFAREA                          0.160 LAYER ME4 ;
 ANTENNAMAXAREACAR                       48.523 LAYER ME2 ;
 ANTENNAMAXAREACAR                       57.782 LAYER ME3 ;
 ANTENNAMAXAREACAR                       67.042 LAYER ME4 ;
END DI38
PIN DO37
  DIRECTION OUTPUT ;
 PORT
  LAYER ME4 ;
  RECT 779.200 0.000 780.000 1.000 ;
  LAYER ME3 ;
  RECT 779.200 0.000 780.000 1.000 ;
  LAYER ME2 ;
  RECT 779.200 0.000 780.000 1.000 ;
  LAYER ME1 ;
  RECT 779.200 0.000 780.000 1.000 ;
 END
 ANTENNAPARTIALMETALAREA                  4.140 LAYER ME2 ;
 ANTENNADIFFAREA                          5.472 LAYER ME2 ;
 ANTENNADIFFAREA                          5.472 LAYER ME3 ;
 ANTENNADIFFAREA                          5.472 LAYER ME4 ;
END DO37
PIN DI37
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 764.400 0.000 765.200 1.000 ;
  LAYER ME3 ;
  RECT 764.400 0.000 765.200 1.000 ;
  LAYER ME2 ;
  RECT 764.400 0.000 765.200 1.000 ;
  LAYER ME1 ;
  RECT 764.400 0.000 765.200 1.000 ;
 END
 ANTENNAPARTIALMETALAREA                  3.150 LAYER ME2 ;
 ANTENNAGATEAREA                          0.086 LAYER ME2 ;
 ANTENNAGATEAREA                          0.086 LAYER ME3 ;
 ANTENNAGATEAREA                          0.086 LAYER ME4 ;
 ANTENNADIFFAREA                          0.160 LAYER ME2 ;
 ANTENNADIFFAREA                          0.160 LAYER ME3 ;
 ANTENNADIFFAREA                          0.160 LAYER ME4 ;
 ANTENNAMAXAREACAR                       48.801 LAYER ME2 ;
 ANTENNAMAXAREACAR                       58.060 LAYER ME3 ;
 ANTENNAMAXAREACAR                       67.319 LAYER ME4 ;
END DI37
PIN DO36
  DIRECTION OUTPUT ;
 PORT
  LAYER ME4 ;
  RECT 759.200 0.000 760.000 1.000 ;
  LAYER ME3 ;
  RECT 759.200 0.000 760.000 1.000 ;
  LAYER ME2 ;
  RECT 759.200 0.000 760.000 1.000 ;
  LAYER ME1 ;
  RECT 759.200 0.000 760.000 1.000 ;
 END
 ANTENNAPARTIALMETALAREA                  4.172 LAYER ME2 ;
 ANTENNADIFFAREA                          5.472 LAYER ME2 ;
 ANTENNADIFFAREA                          5.472 LAYER ME3 ;
 ANTENNADIFFAREA                          5.472 LAYER ME4 ;
END DO36
PIN DI36
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 744.800 0.000 745.600 1.000 ;
  LAYER ME3 ;
  RECT 744.800 0.000 745.600 1.000 ;
  LAYER ME2 ;
  RECT 744.800 0.000 745.600 1.000 ;
  LAYER ME1 ;
  RECT 744.800 0.000 745.600 1.000 ;
 END
 ANTENNAPARTIALMETALAREA                  3.130 LAYER ME2 ;
 ANTENNAGATEAREA                          0.086 LAYER ME2 ;
 ANTENNAGATEAREA                          0.086 LAYER ME3 ;
 ANTENNAGATEAREA                          0.086 LAYER ME4 ;
 ANTENNADIFFAREA                          0.160 LAYER ME2 ;
 ANTENNADIFFAREA                          0.160 LAYER ME3 ;
 ANTENNADIFFAREA                          0.160 LAYER ME4 ;
 ANTENNAMAXAREACAR                       48.569 LAYER ME2 ;
 ANTENNAMAXAREACAR                       57.829 LAYER ME3 ;
 ANTENNAMAXAREACAR                       67.088 LAYER ME4 ;
END DI36
PIN DO35
  DIRECTION OUTPUT ;
 PORT
  LAYER ME4 ;
  RECT 738.400 0.000 739.200 1.000 ;
  LAYER ME3 ;
  RECT 738.400 0.000 739.200 1.000 ;
  LAYER ME2 ;
  RECT 738.400 0.000 739.200 1.000 ;
  LAYER ME1 ;
  RECT 738.400 0.000 739.200 1.000 ;
 END
 ANTENNAPARTIALMETALAREA                  4.164 LAYER ME2 ;
 ANTENNADIFFAREA                          5.472 LAYER ME2 ;
 ANTENNADIFFAREA                          5.472 LAYER ME3 ;
 ANTENNADIFFAREA                          5.472 LAYER ME4 ;
END DO35
PIN DI35
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 723.600 0.000 724.400 1.000 ;
  LAYER ME3 ;
  RECT 723.600 0.000 724.400 1.000 ;
  LAYER ME2 ;
  RECT 723.600 0.000 724.400 1.000 ;
  LAYER ME1 ;
  RECT 723.600 0.000 724.400 1.000 ;
 END
 ANTENNAPARTIALMETALAREA                  3.126 LAYER ME2 ;
 ANTENNAGATEAREA                          0.086 LAYER ME2 ;
 ANTENNAGATEAREA                          0.086 LAYER ME3 ;
 ANTENNAGATEAREA                          0.086 LAYER ME4 ;
 ANTENNADIFFAREA                          0.160 LAYER ME2 ;
 ANTENNADIFFAREA                          0.160 LAYER ME3 ;
 ANTENNADIFFAREA                          0.160 LAYER ME4 ;
 ANTENNAMAXAREACAR                       48.523 LAYER ME2 ;
 ANTENNAMAXAREACAR                       57.782 LAYER ME3 ;
 ANTENNAMAXAREACAR                       67.042 LAYER ME4 ;
END DI35
PIN DO34
  DIRECTION OUTPUT ;
 PORT
  LAYER ME4 ;
  RECT 718.400 0.000 719.200 1.000 ;
  LAYER ME3 ;
  RECT 718.400 0.000 719.200 1.000 ;
  LAYER ME2 ;
  RECT 718.400 0.000 719.200 1.000 ;
  LAYER ME1 ;
  RECT 718.400 0.000 719.200 1.000 ;
 END
 ANTENNAPARTIALMETALAREA                  4.148 LAYER ME2 ;
 ANTENNADIFFAREA                          5.472 LAYER ME2 ;
 ANTENNADIFFAREA                          5.472 LAYER ME3 ;
 ANTENNADIFFAREA                          5.472 LAYER ME4 ;
END DO34
PIN DI34
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 704.000 0.000 704.800 1.000 ;
  LAYER ME3 ;
  RECT 704.000 0.000 704.800 1.000 ;
  LAYER ME2 ;
  RECT 704.000 0.000 704.800 1.000 ;
  LAYER ME1 ;
  RECT 704.000 0.000 704.800 1.000 ;
 END
 ANTENNAPARTIALMETALAREA                  3.154 LAYER ME2 ;
 ANTENNAGATEAREA                          0.086 LAYER ME2 ;
 ANTENNAGATEAREA                          0.086 LAYER ME3 ;
 ANTENNAGATEAREA                          0.086 LAYER ME4 ;
 ANTENNADIFFAREA                          0.160 LAYER ME2 ;
 ANTENNADIFFAREA                          0.160 LAYER ME3 ;
 ANTENNADIFFAREA                          0.160 LAYER ME4 ;
 ANTENNAMAXAREACAR                       48.847 LAYER ME2 ;
 ANTENNAMAXAREACAR                       58.106 LAYER ME3 ;
 ANTENNAMAXAREACAR                       67.366 LAYER ME4 ;
END DI34
PIN DO33
  DIRECTION OUTPUT ;
 PORT
  LAYER ME4 ;
  RECT 697.200 0.000 698.000 1.000 ;
  LAYER ME3 ;
  RECT 697.200 0.000 698.000 1.000 ;
  LAYER ME2 ;
  RECT 697.200 0.000 698.000 1.000 ;
  LAYER ME1 ;
  RECT 697.200 0.000 698.000 1.000 ;
 END
 ANTENNAPARTIALMETALAREA                  4.172 LAYER ME2 ;
 ANTENNADIFFAREA                          5.472 LAYER ME2 ;
 ANTENNADIFFAREA                          5.472 LAYER ME3 ;
 ANTENNADIFFAREA                          5.472 LAYER ME4 ;
END DO33
PIN DI33
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 682.800 0.000 683.600 1.000 ;
  LAYER ME3 ;
  RECT 682.800 0.000 683.600 1.000 ;
  LAYER ME2 ;
  RECT 682.800 0.000 683.600 1.000 ;
  LAYER ME1 ;
  RECT 682.800 0.000 683.600 1.000 ;
 END
 ANTENNAPARTIALMETALAREA                  3.130 LAYER ME2 ;
 ANTENNAGATEAREA                          0.086 LAYER ME2 ;
 ANTENNAGATEAREA                          0.086 LAYER ME3 ;
 ANTENNAGATEAREA                          0.086 LAYER ME4 ;
 ANTENNADIFFAREA                          0.160 LAYER ME2 ;
 ANTENNADIFFAREA                          0.160 LAYER ME3 ;
 ANTENNADIFFAREA                          0.160 LAYER ME4 ;
 ANTENNAMAXAREACAR                       48.569 LAYER ME2 ;
 ANTENNAMAXAREACAR                       57.829 LAYER ME3 ;
 ANTENNAMAXAREACAR                       67.088 LAYER ME4 ;
END DI33
PIN DO32
  DIRECTION OUTPUT ;
 PORT
  LAYER ME4 ;
  RECT 677.600 0.000 678.400 1.000 ;
  LAYER ME3 ;
  RECT 677.600 0.000 678.400 1.000 ;
  LAYER ME2 ;
  RECT 677.600 0.000 678.400 1.000 ;
  LAYER ME1 ;
  RECT 677.600 0.000 678.400 1.000 ;
 END
 ANTENNAPARTIALMETALAREA                  4.156 LAYER ME2 ;
 ANTENNADIFFAREA                          5.472 LAYER ME2 ;
 ANTENNADIFFAREA                          5.472 LAYER ME3 ;
 ANTENNADIFFAREA                          5.472 LAYER ME4 ;
END DO32
PIN WEB4
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 664.800 0.000 665.600 1.000 ;
  LAYER ME3 ;
  RECT 664.800 0.000 665.600 1.000 ;
  LAYER ME2 ;
  RECT 664.800 0.000 665.600 1.000 ;
  LAYER ME1 ;
  RECT 664.800 0.000 665.600 1.000 ;
 END
 ANTENNAPARTIALMETALAREA                  2.868 LAYER ME2 ;
 ANTENNAGATEAREA                          0.072 LAYER ME2 ;
 ANTENNAGATEAREA                          0.072 LAYER ME3 ;
 ANTENNAGATEAREA                          0.072 LAYER ME4 ;
 ANTENNADIFFAREA                          0.160 LAYER ME2 ;
 ANTENNADIFFAREA                          0.160 LAYER ME3 ;
 ANTENNADIFFAREA                          0.160 LAYER ME4 ;
 ANTENNAMAXAREACAR                       54.844 LAYER ME2 ;
 ANTENNAMAXAREACAR                       65.956 LAYER ME3 ;
 ANTENNAMAXAREACAR                       77.067 LAYER ME4 ;
END WEB4
PIN DI32
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 662.800 0.000 663.600 1.000 ;
  LAYER ME3 ;
  RECT 662.800 0.000 663.600 1.000 ;
  LAYER ME2 ;
  RECT 662.800 0.000 663.600 1.000 ;
  LAYER ME1 ;
  RECT 662.800 0.000 663.600 1.000 ;
 END
 ANTENNAPARTIALMETALAREA                  3.134 LAYER ME2 ;
 ANTENNAGATEAREA                          0.086 LAYER ME2 ;
 ANTENNAGATEAREA                          0.086 LAYER ME3 ;
 ANTENNAGATEAREA                          0.086 LAYER ME4 ;
 ANTENNADIFFAREA                          0.160 LAYER ME2 ;
 ANTENNADIFFAREA                          0.160 LAYER ME3 ;
 ANTENNADIFFAREA                          0.160 LAYER ME4 ;
 ANTENNAMAXAREACAR                       48.616 LAYER ME2 ;
 ANTENNAMAXAREACAR                       57.875 LAYER ME3 ;
 ANTENNAMAXAREACAR                       67.134 LAYER ME4 ;
END DI32
PIN DO31
  DIRECTION OUTPUT ;
 PORT
  LAYER ME4 ;
  RECT 656.400 0.000 657.200 1.000 ;
  LAYER ME3 ;
  RECT 656.400 0.000 657.200 1.000 ;
  LAYER ME2 ;
  RECT 656.400 0.000 657.200 1.000 ;
  LAYER ME1 ;
  RECT 656.400 0.000 657.200 1.000 ;
 END
 ANTENNAPARTIALMETALAREA                  4.148 LAYER ME2 ;
 ANTENNADIFFAREA                          5.472 LAYER ME2 ;
 ANTENNADIFFAREA                          5.472 LAYER ME3 ;
 ANTENNADIFFAREA                          5.472 LAYER ME4 ;
END DO31
PIN DI31
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 642.000 0.000 642.800 1.000 ;
  LAYER ME3 ;
  RECT 642.000 0.000 642.800 1.000 ;
  LAYER ME2 ;
  RECT 642.000 0.000 642.800 1.000 ;
  LAYER ME1 ;
  RECT 642.000 0.000 642.800 1.000 ;
 END
 ANTENNAPARTIALMETALAREA                  3.154 LAYER ME2 ;
 ANTENNAGATEAREA                          0.086 LAYER ME2 ;
 ANTENNAGATEAREA                          0.086 LAYER ME3 ;
 ANTENNAGATEAREA                          0.086 LAYER ME4 ;
 ANTENNADIFFAREA                          0.160 LAYER ME2 ;
 ANTENNADIFFAREA                          0.160 LAYER ME3 ;
 ANTENNADIFFAREA                          0.160 LAYER ME4 ;
 ANTENNAMAXAREACAR                       48.847 LAYER ME2 ;
 ANTENNAMAXAREACAR                       58.106 LAYER ME3 ;
 ANTENNAMAXAREACAR                       67.366 LAYER ME4 ;
END DI31
PIN DO30
  DIRECTION OUTPUT ;
 PORT
  LAYER ME4 ;
  RECT 636.400 0.000 637.200 1.000 ;
  LAYER ME3 ;
  RECT 636.400 0.000 637.200 1.000 ;
  LAYER ME2 ;
  RECT 636.400 0.000 637.200 1.000 ;
  LAYER ME1 ;
  RECT 636.400 0.000 637.200 1.000 ;
 END
 ANTENNAPARTIALMETALAREA                  4.180 LAYER ME2 ;
 ANTENNADIFFAREA                          5.472 LAYER ME2 ;
 ANTENNADIFFAREA                          5.472 LAYER ME3 ;
 ANTENNADIFFAREA                          5.472 LAYER ME4 ;
END DO30
PIN DI30
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 622.000 0.000 622.800 1.000 ;
  LAYER ME3 ;
  RECT 622.000 0.000 622.800 1.000 ;
  LAYER ME2 ;
  RECT 622.000 0.000 622.800 1.000 ;
  LAYER ME1 ;
  RECT 622.000 0.000 622.800 1.000 ;
 END
 ANTENNAPARTIALMETALAREA                  3.122 LAYER ME2 ;
 ANTENNAGATEAREA                          0.086 LAYER ME2 ;
 ANTENNAGATEAREA                          0.086 LAYER ME3 ;
 ANTENNAGATEAREA                          0.086 LAYER ME4 ;
 ANTENNADIFFAREA                          0.160 LAYER ME2 ;
 ANTENNADIFFAREA                          0.160 LAYER ME3 ;
 ANTENNADIFFAREA                          0.160 LAYER ME4 ;
 ANTENNAMAXAREACAR                       48.477 LAYER ME2 ;
 ANTENNAMAXAREACAR                       57.736 LAYER ME3 ;
 ANTENNAMAXAREACAR                       66.995 LAYER ME4 ;
END DI30
PIN DO29
  DIRECTION OUTPUT ;
 PORT
  LAYER ME4 ;
  RECT 615.600 0.000 616.400 1.000 ;
  LAYER ME3 ;
  RECT 615.600 0.000 616.400 1.000 ;
  LAYER ME2 ;
  RECT 615.600 0.000 616.400 1.000 ;
  LAYER ME1 ;
  RECT 615.600 0.000 616.400 1.000 ;
 END
 ANTENNAPARTIALMETALAREA                  4.156 LAYER ME2 ;
 ANTENNADIFFAREA                          5.472 LAYER ME2 ;
 ANTENNADIFFAREA                          5.472 LAYER ME3 ;
 ANTENNADIFFAREA                          5.472 LAYER ME4 ;
END DO29
PIN DI29
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 600.800 0.000 601.600 1.000 ;
  LAYER ME3 ;
  RECT 600.800 0.000 601.600 1.000 ;
  LAYER ME2 ;
  RECT 600.800 0.000 601.600 1.000 ;
  LAYER ME1 ;
  RECT 600.800 0.000 601.600 1.000 ;
 END
 ANTENNAPARTIALMETALAREA                  3.134 LAYER ME2 ;
 ANTENNAGATEAREA                          0.086 LAYER ME2 ;
 ANTENNAGATEAREA                          0.086 LAYER ME3 ;
 ANTENNAGATEAREA                          0.086 LAYER ME4 ;
 ANTENNADIFFAREA                          0.160 LAYER ME2 ;
 ANTENNADIFFAREA                          0.160 LAYER ME3 ;
 ANTENNADIFFAREA                          0.160 LAYER ME4 ;
 ANTENNAMAXAREACAR                       48.616 LAYER ME2 ;
 ANTENNAMAXAREACAR                       57.875 LAYER ME3 ;
 ANTENNAMAXAREACAR                       67.134 LAYER ME4 ;
END DI29
PIN DO28
  DIRECTION OUTPUT ;
 PORT
  LAYER ME4 ;
  RECT 595.600 0.000 596.400 1.000 ;
  LAYER ME3 ;
  RECT 595.600 0.000 596.400 1.000 ;
  LAYER ME2 ;
  RECT 595.600 0.000 596.400 1.000 ;
  LAYER ME1 ;
  RECT 595.600 0.000 596.400 1.000 ;
 END
 ANTENNAPARTIALMETALAREA                  4.156 LAYER ME2 ;
 ANTENNADIFFAREA                          5.472 LAYER ME2 ;
 ANTENNADIFFAREA                          5.472 LAYER ME3 ;
 ANTENNADIFFAREA                          5.472 LAYER ME4 ;
END DO28
PIN DI28
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 581.200 0.000 582.000 1.000 ;
  LAYER ME3 ;
  RECT 581.200 0.000 582.000 1.000 ;
  LAYER ME2 ;
  RECT 581.200 0.000 582.000 1.000 ;
  LAYER ME1 ;
  RECT 581.200 0.000 582.000 1.000 ;
 END
 ANTENNAPARTIALMETALAREA                  3.146 LAYER ME2 ;
 ANTENNAGATEAREA                          0.086 LAYER ME2 ;
 ANTENNAGATEAREA                          0.086 LAYER ME3 ;
 ANTENNAGATEAREA                          0.086 LAYER ME4 ;
 ANTENNADIFFAREA                          0.160 LAYER ME2 ;
 ANTENNADIFFAREA                          0.160 LAYER ME3 ;
 ANTENNADIFFAREA                          0.160 LAYER ME4 ;
 ANTENNAMAXAREACAR                       48.755 LAYER ME2 ;
 ANTENNAMAXAREACAR                       58.014 LAYER ME3 ;
 ANTENNAMAXAREACAR                       67.273 LAYER ME4 ;
END DI28
PIN DO27
  DIRECTION OUTPUT ;
 PORT
  LAYER ME4 ;
  RECT 574.400 0.000 575.200 1.000 ;
  LAYER ME3 ;
  RECT 574.400 0.000 575.200 1.000 ;
  LAYER ME2 ;
  RECT 574.400 0.000 575.200 1.000 ;
  LAYER ME1 ;
  RECT 574.400 0.000 575.200 1.000 ;
 END
 ANTENNAPARTIALMETALAREA                  4.180 LAYER ME2 ;
 ANTENNADIFFAREA                          5.472 LAYER ME2 ;
 ANTENNADIFFAREA                          5.472 LAYER ME3 ;
 ANTENNADIFFAREA                          5.472 LAYER ME4 ;
END DO27
PIN DI27
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 560.000 0.000 560.800 1.000 ;
  LAYER ME3 ;
  RECT 560.000 0.000 560.800 1.000 ;
  LAYER ME2 ;
  RECT 560.000 0.000 560.800 1.000 ;
  LAYER ME1 ;
  RECT 560.000 0.000 560.800 1.000 ;
 END
 ANTENNAPARTIALMETALAREA                  3.122 LAYER ME2 ;
 ANTENNAGATEAREA                          0.086 LAYER ME2 ;
 ANTENNAGATEAREA                          0.086 LAYER ME3 ;
 ANTENNAGATEAREA                          0.086 LAYER ME4 ;
 ANTENNADIFFAREA                          0.160 LAYER ME2 ;
 ANTENNADIFFAREA                          0.160 LAYER ME3 ;
 ANTENNADIFFAREA                          0.160 LAYER ME4 ;
 ANTENNAMAXAREACAR                       48.477 LAYER ME2 ;
 ANTENNAMAXAREACAR                       57.736 LAYER ME3 ;
 ANTENNAMAXAREACAR                       66.995 LAYER ME4 ;
END DI27
PIN DO26
  DIRECTION OUTPUT ;
 PORT
  LAYER ME4 ;
  RECT 554.800 0.000 555.600 1.000 ;
  LAYER ME3 ;
  RECT 554.800 0.000 555.600 1.000 ;
  LAYER ME2 ;
  RECT 554.800 0.000 555.600 1.000 ;
  LAYER ME1 ;
  RECT 554.800 0.000 555.600 1.000 ;
 END
 ANTENNAPARTIALMETALAREA                  4.148 LAYER ME2 ;
 ANTENNADIFFAREA                          5.472 LAYER ME2 ;
 ANTENNADIFFAREA                          5.472 LAYER ME3 ;
 ANTENNADIFFAREA                          5.472 LAYER ME4 ;
END DO26
PIN DI26
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 540.000 0.000 540.800 1.000 ;
  LAYER ME3 ;
  RECT 540.000 0.000 540.800 1.000 ;
  LAYER ME2 ;
  RECT 540.000 0.000 540.800 1.000 ;
  LAYER ME1 ;
  RECT 540.000 0.000 540.800 1.000 ;
 END
 ANTENNAPARTIALMETALAREA                  3.142 LAYER ME2 ;
 ANTENNAGATEAREA                          0.086 LAYER ME2 ;
 ANTENNAGATEAREA                          0.086 LAYER ME3 ;
 ANTENNAGATEAREA                          0.086 LAYER ME4 ;
 ANTENNADIFFAREA                          0.160 LAYER ME2 ;
 ANTENNADIFFAREA                          0.160 LAYER ME3 ;
 ANTENNADIFFAREA                          0.160 LAYER ME4 ;
 ANTENNAMAXAREACAR                       48.708 LAYER ME2 ;
 ANTENNAMAXAREACAR                       57.968 LAYER ME3 ;
 ANTENNAMAXAREACAR                       67.227 LAYER ME4 ;
END DI26
PIN DO25
  DIRECTION OUTPUT ;
 PORT
  LAYER ME4 ;
  RECT 533.600 0.000 534.400 1.000 ;
  LAYER ME3 ;
  RECT 533.600 0.000 534.400 1.000 ;
  LAYER ME2 ;
  RECT 533.600 0.000 534.400 1.000 ;
  LAYER ME1 ;
  RECT 533.600 0.000 534.400 1.000 ;
 END
 ANTENNAPARTIALMETALAREA                  4.156 LAYER ME2 ;
 ANTENNADIFFAREA                          5.472 LAYER ME2 ;
 ANTENNADIFFAREA                          5.472 LAYER ME3 ;
 ANTENNADIFFAREA                          5.472 LAYER ME4 ;
END DO25
PIN DI25
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 519.200 0.000 520.000 1.000 ;
  LAYER ME3 ;
  RECT 519.200 0.000 520.000 1.000 ;
  LAYER ME2 ;
  RECT 519.200 0.000 520.000 1.000 ;
  LAYER ME1 ;
  RECT 519.200 0.000 520.000 1.000 ;
 END
 ANTENNAPARTIALMETALAREA                  3.146 LAYER ME2 ;
 ANTENNAGATEAREA                          0.086 LAYER ME2 ;
 ANTENNAGATEAREA                          0.086 LAYER ME3 ;
 ANTENNAGATEAREA                          0.086 LAYER ME4 ;
 ANTENNADIFFAREA                          0.160 LAYER ME2 ;
 ANTENNADIFFAREA                          0.160 LAYER ME3 ;
 ANTENNADIFFAREA                          0.160 LAYER ME4 ;
 ANTENNAMAXAREACAR                       48.755 LAYER ME2 ;
 ANTENNAMAXAREACAR                       58.014 LAYER ME3 ;
 ANTENNAMAXAREACAR                       67.273 LAYER ME4 ;
END DI25
PIN DO24
  DIRECTION OUTPUT ;
 PORT
  LAYER ME4 ;
  RECT 514.000 0.000 514.800 1.000 ;
  LAYER ME3 ;
  RECT 514.000 0.000 514.800 1.000 ;
  LAYER ME2 ;
  RECT 514.000 0.000 514.800 1.000 ;
  LAYER ME1 ;
  RECT 514.000 0.000 514.800 1.000 ;
 END
 ANTENNAPARTIALMETALAREA                  4.172 LAYER ME2 ;
 ANTENNADIFFAREA                          5.472 LAYER ME2 ;
 ANTENNADIFFAREA                          5.472 LAYER ME3 ;
 ANTENNADIFFAREA                          5.472 LAYER ME4 ;
END DO24
PIN WEB3
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 500.800 0.000 501.600 1.000 ;
  LAYER ME3 ;
  RECT 500.800 0.000 501.600 1.000 ;
  LAYER ME2 ;
  RECT 500.800 0.000 501.600 1.000 ;
  LAYER ME1 ;
  RECT 500.800 0.000 501.600 1.000 ;
 END
 ANTENNAPARTIALMETALAREA                  2.856 LAYER ME2 ;
 ANTENNAGATEAREA                          0.072 LAYER ME2 ;
 ANTENNAGATEAREA                          0.072 LAYER ME3 ;
 ANTENNAGATEAREA                          0.072 LAYER ME4 ;
 ANTENNADIFFAREA                          0.160 LAYER ME2 ;
 ANTENNADIFFAREA                          0.160 LAYER ME3 ;
 ANTENNADIFFAREA                          0.160 LAYER ME4 ;
 ANTENNAMAXAREACAR                       54.678 LAYER ME2 ;
 ANTENNAMAXAREACAR                       65.789 LAYER ME3 ;
 ANTENNAMAXAREACAR                       76.900 LAYER ME4 ;
END WEB3
PIN DI24
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 499.200 0.000 500.000 1.000 ;
  LAYER ME3 ;
  RECT 499.200 0.000 500.000 1.000 ;
  LAYER ME2 ;
  RECT 499.200 0.000 500.000 1.000 ;
  LAYER ME1 ;
  RECT 499.200 0.000 500.000 1.000 ;
 END
 ANTENNAPARTIALMETALAREA                  3.118 LAYER ME2 ;
 ANTENNAGATEAREA                          0.086 LAYER ME2 ;
 ANTENNAGATEAREA                          0.086 LAYER ME3 ;
 ANTENNAGATEAREA                          0.086 LAYER ME4 ;
 ANTENNADIFFAREA                          0.160 LAYER ME2 ;
 ANTENNADIFFAREA                          0.160 LAYER ME3 ;
 ANTENNADIFFAREA                          0.160 LAYER ME4 ;
 ANTENNAMAXAREACAR                       48.431 LAYER ME2 ;
 ANTENNAMAXAREACAR                       57.690 LAYER ME3 ;
 ANTENNAMAXAREACAR                       66.949 LAYER ME4 ;
END DI24
PIN DO23
  DIRECTION OUTPUT ;
 PORT
  LAYER ME4 ;
  RECT 492.800 0.000 493.600 1.000 ;
  LAYER ME3 ;
  RECT 492.800 0.000 493.600 1.000 ;
  LAYER ME2 ;
  RECT 492.800 0.000 493.600 1.000 ;
  LAYER ME1 ;
  RECT 492.800 0.000 493.600 1.000 ;
 END
 ANTENNAPARTIALMETALAREA                  4.148 LAYER ME2 ;
 ANTENNADIFFAREA                          5.472 LAYER ME2 ;
 ANTENNADIFFAREA                          5.472 LAYER ME3 ;
 ANTENNADIFFAREA                          5.472 LAYER ME4 ;
END DO23
PIN DI23
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 478.000 0.000 478.800 1.000 ;
  LAYER ME3 ;
  RECT 478.000 0.000 478.800 1.000 ;
  LAYER ME2 ;
  RECT 478.000 0.000 478.800 1.000 ;
  LAYER ME1 ;
  RECT 478.000 0.000 478.800 1.000 ;
 END
 ANTENNAPARTIALMETALAREA                  3.142 LAYER ME2 ;
 ANTENNAGATEAREA                          0.086 LAYER ME2 ;
 ANTENNAGATEAREA                          0.086 LAYER ME3 ;
 ANTENNAGATEAREA                          0.086 LAYER ME4 ;
 ANTENNADIFFAREA                          0.160 LAYER ME2 ;
 ANTENNADIFFAREA                          0.160 LAYER ME3 ;
 ANTENNADIFFAREA                          0.160 LAYER ME4 ;
 ANTENNAMAXAREACAR                       48.708 LAYER ME2 ;
 ANTENNAMAXAREACAR                       57.968 LAYER ME3 ;
 ANTENNAMAXAREACAR                       67.227 LAYER ME4 ;
END DI23
PIN DO22
  DIRECTION OUTPUT ;
 PORT
  LAYER ME4 ;
  RECT 472.800 0.000 473.600 1.000 ;
  LAYER ME3 ;
  RECT 472.800 0.000 473.600 1.000 ;
  LAYER ME2 ;
  RECT 472.800 0.000 473.600 1.000 ;
  LAYER ME1 ;
  RECT 472.800 0.000 473.600 1.000 ;
 END
 ANTENNAPARTIALMETALAREA                  4.164 LAYER ME2 ;
 ANTENNADIFFAREA                          5.472 LAYER ME2 ;
 ANTENNADIFFAREA                          5.472 LAYER ME3 ;
 ANTENNADIFFAREA                          5.472 LAYER ME4 ;
END DO22
PIN DI22
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 458.400 0.000 459.200 1.000 ;
  LAYER ME3 ;
  RECT 458.400 0.000 459.200 1.000 ;
  LAYER ME2 ;
  RECT 458.400 0.000 459.200 1.000 ;
  LAYER ME1 ;
  RECT 458.400 0.000 459.200 1.000 ;
 END
 ANTENNAPARTIALMETALAREA                  3.138 LAYER ME2 ;
 ANTENNAGATEAREA                          0.086 LAYER ME2 ;
 ANTENNAGATEAREA                          0.086 LAYER ME3 ;
 ANTENNAGATEAREA                          0.086 LAYER ME4 ;
 ANTENNADIFFAREA                          0.160 LAYER ME2 ;
 ANTENNADIFFAREA                          0.160 LAYER ME3 ;
 ANTENNADIFFAREA                          0.160 LAYER ME4 ;
 ANTENNAMAXAREACAR                       48.662 LAYER ME2 ;
 ANTENNAMAXAREACAR                       57.921 LAYER ME3 ;
 ANTENNAMAXAREACAR                       67.181 LAYER ME4 ;
END DI22
PIN DO21
  DIRECTION OUTPUT ;
 PORT
  LAYER ME4 ;
  RECT 452.000 0.000 452.800 1.000 ;
  LAYER ME3 ;
  RECT 452.000 0.000 452.800 1.000 ;
  LAYER ME2 ;
  RECT 452.000 0.000 452.800 1.000 ;
  LAYER ME1 ;
  RECT 452.000 0.000 452.800 1.000 ;
 END
 ANTENNAPARTIALMETALAREA                  4.172 LAYER ME2 ;
 ANTENNADIFFAREA                          5.472 LAYER ME2 ;
 ANTENNADIFFAREA                          5.472 LAYER ME3 ;
 ANTENNADIFFAREA                          5.472 LAYER ME4 ;
END DO21
PIN DI21
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 437.200 0.000 438.000 1.000 ;
  LAYER ME3 ;
  RECT 437.200 0.000 438.000 1.000 ;
  LAYER ME2 ;
  RECT 437.200 0.000 438.000 1.000 ;
  LAYER ME1 ;
  RECT 437.200 0.000 438.000 1.000 ;
 END
 ANTENNAPARTIALMETALAREA                  3.118 LAYER ME2 ;
 ANTENNAGATEAREA                          0.086 LAYER ME2 ;
 ANTENNAGATEAREA                          0.086 LAYER ME3 ;
 ANTENNAGATEAREA                          0.086 LAYER ME4 ;
 ANTENNADIFFAREA                          0.160 LAYER ME2 ;
 ANTENNADIFFAREA                          0.160 LAYER ME3 ;
 ANTENNADIFFAREA                          0.160 LAYER ME4 ;
 ANTENNAMAXAREACAR                       48.431 LAYER ME2 ;
 ANTENNAMAXAREACAR                       57.690 LAYER ME3 ;
 ANTENNAMAXAREACAR                       66.949 LAYER ME4 ;
END DI21
PIN DO20
  DIRECTION OUTPUT ;
 PORT
  LAYER ME4 ;
  RECT 432.000 0.000 432.800 1.000 ;
  LAYER ME3 ;
  RECT 432.000 0.000 432.800 1.000 ;
  LAYER ME2 ;
  RECT 432.000 0.000 432.800 1.000 ;
  LAYER ME1 ;
  RECT 432.000 0.000 432.800 1.000 ;
 END
 ANTENNAPARTIALMETALAREA                  4.140 LAYER ME2 ;
 ANTENNADIFFAREA                          5.472 LAYER ME2 ;
 ANTENNADIFFAREA                          5.472 LAYER ME3 ;
 ANTENNADIFFAREA                          5.472 LAYER ME4 ;
END DO20
PIN DI20
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 417.200 0.000 418.000 1.000 ;
  LAYER ME3 ;
  RECT 417.200 0.000 418.000 1.000 ;
  LAYER ME2 ;
  RECT 417.200 0.000 418.000 1.000 ;
  LAYER ME1 ;
  RECT 417.200 0.000 418.000 1.000 ;
 END
 ANTENNAPARTIALMETALAREA                  3.150 LAYER ME2 ;
 ANTENNAGATEAREA                          0.086 LAYER ME2 ;
 ANTENNAGATEAREA                          0.086 LAYER ME3 ;
 ANTENNAGATEAREA                          0.086 LAYER ME4 ;
 ANTENNADIFFAREA                          0.160 LAYER ME2 ;
 ANTENNADIFFAREA                          0.160 LAYER ME3 ;
 ANTENNADIFFAREA                          0.160 LAYER ME4 ;
 ANTENNAMAXAREACAR                       48.801 LAYER ME2 ;
 ANTENNAMAXAREACAR                       58.060 LAYER ME3 ;
 ANTENNAMAXAREACAR                       67.319 LAYER ME4 ;
END DI20
PIN DO19
  DIRECTION OUTPUT ;
 PORT
  LAYER ME4 ;
  RECT 410.800 0.000 411.600 1.000 ;
  LAYER ME3 ;
  RECT 410.800 0.000 411.600 1.000 ;
  LAYER ME2 ;
  RECT 410.800 0.000 411.600 1.000 ;
  LAYER ME1 ;
  RECT 410.800 0.000 411.600 1.000 ;
 END
 ANTENNAPARTIALMETALAREA                  4.164 LAYER ME2 ;
 ANTENNADIFFAREA                          5.472 LAYER ME2 ;
 ANTENNADIFFAREA                          5.472 LAYER ME3 ;
 ANTENNADIFFAREA                          5.472 LAYER ME4 ;
END DO19
PIN DI19
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 396.400 0.000 397.200 1.000 ;
  LAYER ME3 ;
  RECT 396.400 0.000 397.200 1.000 ;
  LAYER ME2 ;
  RECT 396.400 0.000 397.200 1.000 ;
  LAYER ME1 ;
  RECT 396.400 0.000 397.200 1.000 ;
 END
 ANTENNAPARTIALMETALAREA                  3.138 LAYER ME2 ;
 ANTENNAGATEAREA                          0.086 LAYER ME2 ;
 ANTENNAGATEAREA                          0.086 LAYER ME3 ;
 ANTENNAGATEAREA                          0.086 LAYER ME4 ;
 ANTENNADIFFAREA                          0.160 LAYER ME2 ;
 ANTENNADIFFAREA                          0.160 LAYER ME3 ;
 ANTENNADIFFAREA                          0.160 LAYER ME4 ;
 ANTENNAMAXAREACAR                       48.662 LAYER ME2 ;
 ANTENNAMAXAREACAR                       57.921 LAYER ME3 ;
 ANTENNAMAXAREACAR                       67.181 LAYER ME4 ;
END DI19
PIN DO18
  DIRECTION OUTPUT ;
 PORT
  LAYER ME4 ;
  RECT 391.200 0.000 392.000 1.000 ;
  LAYER ME3 ;
  RECT 391.200 0.000 392.000 1.000 ;
  LAYER ME2 ;
  RECT 391.200 0.000 392.000 1.000 ;
  LAYER ME1 ;
  RECT 391.200 0.000 392.000 1.000 ;
 END
 ANTENNAPARTIALMETALAREA                  4.164 LAYER ME2 ;
 ANTENNADIFFAREA                          5.472 LAYER ME2 ;
 ANTENNADIFFAREA                          5.472 LAYER ME3 ;
 ANTENNADIFFAREA                          5.472 LAYER ME4 ;
END DO18
PIN DI18
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 376.400 0.000 377.200 1.000 ;
  LAYER ME3 ;
  RECT 376.400 0.000 377.200 1.000 ;
  LAYER ME2 ;
  RECT 376.400 0.000 377.200 1.000 ;
  LAYER ME1 ;
  RECT 376.400 0.000 377.200 1.000 ;
 END
 ANTENNAPARTIALMETALAREA                  3.126 LAYER ME2 ;
 ANTENNAGATEAREA                          0.086 LAYER ME2 ;
 ANTENNAGATEAREA                          0.086 LAYER ME3 ;
 ANTENNAGATEAREA                          0.086 LAYER ME4 ;
 ANTENNADIFFAREA                          0.160 LAYER ME2 ;
 ANTENNADIFFAREA                          0.160 LAYER ME3 ;
 ANTENNADIFFAREA                          0.160 LAYER ME4 ;
 ANTENNAMAXAREACAR                       48.523 LAYER ME2 ;
 ANTENNAMAXAREACAR                       57.782 LAYER ME3 ;
 ANTENNAMAXAREACAR                       67.042 LAYER ME4 ;
END DI18
PIN DO17
  DIRECTION OUTPUT ;
 PORT
  LAYER ME4 ;
  RECT 370.000 0.000 370.800 1.000 ;
  LAYER ME3 ;
  RECT 370.000 0.000 370.800 1.000 ;
  LAYER ME2 ;
  RECT 370.000 0.000 370.800 1.000 ;
  LAYER ME1 ;
  RECT 370.000 0.000 370.800 1.000 ;
 END
 ANTENNAPARTIALMETALAREA                  4.140 LAYER ME2 ;
 ANTENNADIFFAREA                          5.472 LAYER ME2 ;
 ANTENNADIFFAREA                          5.472 LAYER ME3 ;
 ANTENNADIFFAREA                          5.472 LAYER ME4 ;
END DO17
PIN DI17
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 355.200 0.000 356.000 1.000 ;
  LAYER ME3 ;
  RECT 355.200 0.000 356.000 1.000 ;
  LAYER ME2 ;
  RECT 355.200 0.000 356.000 1.000 ;
  LAYER ME1 ;
  RECT 355.200 0.000 356.000 1.000 ;
 END
 ANTENNAPARTIALMETALAREA                  3.150 LAYER ME2 ;
 ANTENNAGATEAREA                          0.086 LAYER ME2 ;
 ANTENNAGATEAREA                          0.086 LAYER ME3 ;
 ANTENNAGATEAREA                          0.086 LAYER ME4 ;
 ANTENNADIFFAREA                          0.160 LAYER ME2 ;
 ANTENNADIFFAREA                          0.160 LAYER ME3 ;
 ANTENNADIFFAREA                          0.160 LAYER ME4 ;
 ANTENNAMAXAREACAR                       48.801 LAYER ME2 ;
 ANTENNAMAXAREACAR                       58.060 LAYER ME3 ;
 ANTENNAMAXAREACAR                       67.319 LAYER ME4 ;
END DI17
PIN DO16
  DIRECTION OUTPUT ;
 PORT
  LAYER ME4 ;
  RECT 350.000 0.000 350.800 1.000 ;
  LAYER ME3 ;
  RECT 350.000 0.000 350.800 1.000 ;
  LAYER ME2 ;
  RECT 350.000 0.000 350.800 1.000 ;
  LAYER ME1 ;
  RECT 350.000 0.000 350.800 1.000 ;
 END
 ANTENNAPARTIALMETALAREA                  4.172 LAYER ME2 ;
 ANTENNADIFFAREA                          5.472 LAYER ME2 ;
 ANTENNADIFFAREA                          5.472 LAYER ME3 ;
 ANTENNADIFFAREA                          5.472 LAYER ME4 ;
END DO16
PIN WEB2
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 337.200 0.000 338.000 1.000 ;
  LAYER ME3 ;
  RECT 337.200 0.000 338.000 1.000 ;
  LAYER ME2 ;
  RECT 337.200 0.000 338.000 1.000 ;
  LAYER ME1 ;
  RECT 337.200 0.000 338.000 1.000 ;
 END
 ANTENNAPARTIALMETALAREA                  2.840 LAYER ME2 ;
 ANTENNAGATEAREA                          0.072 LAYER ME2 ;
 ANTENNAGATEAREA                          0.072 LAYER ME3 ;
 ANTENNAGATEAREA                          0.072 LAYER ME4 ;
 ANTENNADIFFAREA                          0.160 LAYER ME2 ;
 ANTENNADIFFAREA                          0.160 LAYER ME3 ;
 ANTENNADIFFAREA                          0.160 LAYER ME4 ;
 ANTENNAMAXAREACAR                       54.456 LAYER ME2 ;
 ANTENNAMAXAREACAR                       65.567 LAYER ME3 ;
 ANTENNAMAXAREACAR                       76.678 LAYER ME4 ;
END WEB2
PIN DI16
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 335.600 0.000 336.400 1.000 ;
  LAYER ME3 ;
  RECT 335.600 0.000 336.400 1.000 ;
  LAYER ME2 ;
  RECT 335.600 0.000 336.400 1.000 ;
  LAYER ME1 ;
  RECT 335.600 0.000 336.400 1.000 ;
 END
 ANTENNAPARTIALMETALAREA                  3.130 LAYER ME2 ;
 ANTENNAGATEAREA                          0.086 LAYER ME2 ;
 ANTENNAGATEAREA                          0.086 LAYER ME3 ;
 ANTENNAGATEAREA                          0.086 LAYER ME4 ;
 ANTENNADIFFAREA                          0.160 LAYER ME2 ;
 ANTENNADIFFAREA                          0.160 LAYER ME3 ;
 ANTENNADIFFAREA                          0.160 LAYER ME4 ;
 ANTENNAMAXAREACAR                       48.569 LAYER ME2 ;
 ANTENNAMAXAREACAR                       57.829 LAYER ME3 ;
 ANTENNAMAXAREACAR                       67.088 LAYER ME4 ;
END DI16
PIN DO15
  DIRECTION OUTPUT ;
 PORT
  LAYER ME4 ;
  RECT 329.200 0.000 330.000 1.000 ;
  LAYER ME3 ;
  RECT 329.200 0.000 330.000 1.000 ;
  LAYER ME2 ;
  RECT 329.200 0.000 330.000 1.000 ;
  LAYER ME1 ;
  RECT 329.200 0.000 330.000 1.000 ;
 END
 ANTENNAPARTIALMETALAREA                  4.164 LAYER ME2 ;
 ANTENNADIFFAREA                          5.472 LAYER ME2 ;
 ANTENNADIFFAREA                          5.472 LAYER ME3 ;
 ANTENNADIFFAREA                          5.472 LAYER ME4 ;
END DO15
PIN DI15
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 314.400 0.000 315.200 1.000 ;
  LAYER ME3 ;
  RECT 314.400 0.000 315.200 1.000 ;
  LAYER ME2 ;
  RECT 314.400 0.000 315.200 1.000 ;
  LAYER ME1 ;
  RECT 314.400 0.000 315.200 1.000 ;
 END
 ANTENNAPARTIALMETALAREA                  3.126 LAYER ME2 ;
 ANTENNAGATEAREA                          0.086 LAYER ME2 ;
 ANTENNAGATEAREA                          0.086 LAYER ME3 ;
 ANTENNAGATEAREA                          0.086 LAYER ME4 ;
 ANTENNADIFFAREA                          0.160 LAYER ME2 ;
 ANTENNADIFFAREA                          0.160 LAYER ME3 ;
 ANTENNADIFFAREA                          0.160 LAYER ME4 ;
 ANTENNAMAXAREACAR                       48.523 LAYER ME2 ;
 ANTENNAMAXAREACAR                       57.782 LAYER ME3 ;
 ANTENNAMAXAREACAR                       67.042 LAYER ME4 ;
END DI15
PIN DO14
  DIRECTION OUTPUT ;
 PORT
  LAYER ME4 ;
  RECT 309.200 0.000 310.000 1.000 ;
  LAYER ME3 ;
  RECT 309.200 0.000 310.000 1.000 ;
  LAYER ME2 ;
  RECT 309.200 0.000 310.000 1.000 ;
  LAYER ME1 ;
  RECT 309.200 0.000 310.000 1.000 ;
 END
 ANTENNAPARTIALMETALAREA                  4.148 LAYER ME2 ;
 ANTENNADIFFAREA                          5.472 LAYER ME2 ;
 ANTENNADIFFAREA                          5.472 LAYER ME3 ;
 ANTENNADIFFAREA                          5.472 LAYER ME4 ;
END DO14
PIN DI14
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 294.800 0.000 295.600 1.000 ;
  LAYER ME3 ;
  RECT 294.800 0.000 295.600 1.000 ;
  LAYER ME2 ;
  RECT 294.800 0.000 295.600 1.000 ;
  LAYER ME1 ;
  RECT 294.800 0.000 295.600 1.000 ;
 END
 ANTENNAPARTIALMETALAREA                  3.154 LAYER ME2 ;
 ANTENNAGATEAREA                          0.086 LAYER ME2 ;
 ANTENNAGATEAREA                          0.086 LAYER ME3 ;
 ANTENNAGATEAREA                          0.086 LAYER ME4 ;
 ANTENNADIFFAREA                          0.160 LAYER ME2 ;
 ANTENNADIFFAREA                          0.160 LAYER ME3 ;
 ANTENNADIFFAREA                          0.160 LAYER ME4 ;
 ANTENNAMAXAREACAR                       48.847 LAYER ME2 ;
 ANTENNAMAXAREACAR                       58.106 LAYER ME3 ;
 ANTENNAMAXAREACAR                       67.366 LAYER ME4 ;
END DI14
PIN DO13
  DIRECTION OUTPUT ;
 PORT
  LAYER ME4 ;
  RECT 288.000 0.000 288.800 1.000 ;
  LAYER ME3 ;
  RECT 288.000 0.000 288.800 1.000 ;
  LAYER ME2 ;
  RECT 288.000 0.000 288.800 1.000 ;
  LAYER ME1 ;
  RECT 288.000 0.000 288.800 1.000 ;
 END
 ANTENNAPARTIALMETALAREA                  4.172 LAYER ME2 ;
 ANTENNADIFFAREA                          5.472 LAYER ME2 ;
 ANTENNADIFFAREA                          5.472 LAYER ME3 ;
 ANTENNADIFFAREA                          5.472 LAYER ME4 ;
END DO13
PIN DI13
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 273.600 0.000 274.400 1.000 ;
  LAYER ME3 ;
  RECT 273.600 0.000 274.400 1.000 ;
  LAYER ME2 ;
  RECT 273.600 0.000 274.400 1.000 ;
  LAYER ME1 ;
  RECT 273.600 0.000 274.400 1.000 ;
 END
 ANTENNAPARTIALMETALAREA                  3.130 LAYER ME2 ;
 ANTENNAGATEAREA                          0.086 LAYER ME2 ;
 ANTENNAGATEAREA                          0.086 LAYER ME3 ;
 ANTENNAGATEAREA                          0.086 LAYER ME4 ;
 ANTENNADIFFAREA                          0.160 LAYER ME2 ;
 ANTENNADIFFAREA                          0.160 LAYER ME3 ;
 ANTENNADIFFAREA                          0.160 LAYER ME4 ;
 ANTENNAMAXAREACAR                       48.569 LAYER ME2 ;
 ANTENNAMAXAREACAR                       57.829 LAYER ME3 ;
 ANTENNAMAXAREACAR                       67.088 LAYER ME4 ;
END DI13
PIN DO12
  DIRECTION OUTPUT ;
 PORT
  LAYER ME4 ;
  RECT 268.400 0.000 269.200 1.000 ;
  LAYER ME3 ;
  RECT 268.400 0.000 269.200 1.000 ;
  LAYER ME2 ;
  RECT 268.400 0.000 269.200 1.000 ;
  LAYER ME1 ;
  RECT 268.400 0.000 269.200 1.000 ;
 END
 ANTENNAPARTIALMETALAREA                  4.156 LAYER ME2 ;
 ANTENNADIFFAREA                          5.472 LAYER ME2 ;
 ANTENNADIFFAREA                          5.472 LAYER ME3 ;
 ANTENNADIFFAREA                          5.472 LAYER ME4 ;
END DO12
PIN DI12
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 253.600 0.000 254.400 1.000 ;
  LAYER ME3 ;
  RECT 253.600 0.000 254.400 1.000 ;
  LAYER ME2 ;
  RECT 253.600 0.000 254.400 1.000 ;
  LAYER ME1 ;
  RECT 253.600 0.000 254.400 1.000 ;
 END
 ANTENNAPARTIALMETALAREA                  3.134 LAYER ME2 ;
 ANTENNAGATEAREA                          0.086 LAYER ME2 ;
 ANTENNAGATEAREA                          0.086 LAYER ME3 ;
 ANTENNAGATEAREA                          0.086 LAYER ME4 ;
 ANTENNADIFFAREA                          0.160 LAYER ME2 ;
 ANTENNADIFFAREA                          0.160 LAYER ME3 ;
 ANTENNADIFFAREA                          0.160 LAYER ME4 ;
 ANTENNAMAXAREACAR                       48.616 LAYER ME2 ;
 ANTENNAMAXAREACAR                       57.875 LAYER ME3 ;
 ANTENNAMAXAREACAR                       67.134 LAYER ME4 ;
END DI12
PIN DO11
  DIRECTION OUTPUT ;
 PORT
  LAYER ME4 ;
  RECT 247.200 0.000 248.000 1.000 ;
  LAYER ME3 ;
  RECT 247.200 0.000 248.000 1.000 ;
  LAYER ME2 ;
  RECT 247.200 0.000 248.000 1.000 ;
  LAYER ME1 ;
  RECT 247.200 0.000 248.000 1.000 ;
 END
 ANTENNAPARTIALMETALAREA                  4.148 LAYER ME2 ;
 ANTENNADIFFAREA                          5.472 LAYER ME2 ;
 ANTENNADIFFAREA                          5.472 LAYER ME3 ;
 ANTENNADIFFAREA                          5.472 LAYER ME4 ;
END DO11
PIN DI11
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 232.800 0.000 233.600 1.000 ;
  LAYER ME3 ;
  RECT 232.800 0.000 233.600 1.000 ;
  LAYER ME2 ;
  RECT 232.800 0.000 233.600 1.000 ;
  LAYER ME1 ;
  RECT 232.800 0.000 233.600 1.000 ;
 END
 ANTENNAPARTIALMETALAREA                  3.154 LAYER ME2 ;
 ANTENNAGATEAREA                          0.086 LAYER ME2 ;
 ANTENNAGATEAREA                          0.086 LAYER ME3 ;
 ANTENNAGATEAREA                          0.086 LAYER ME4 ;
 ANTENNADIFFAREA                          0.160 LAYER ME2 ;
 ANTENNADIFFAREA                          0.160 LAYER ME3 ;
 ANTENNADIFFAREA                          0.160 LAYER ME4 ;
 ANTENNAMAXAREACAR                       48.847 LAYER ME2 ;
 ANTENNAMAXAREACAR                       58.106 LAYER ME3 ;
 ANTENNAMAXAREACAR                       67.366 LAYER ME4 ;
END DI11
PIN DO10
  DIRECTION OUTPUT ;
 PORT
  LAYER ME4 ;
  RECT 227.200 0.000 228.000 1.000 ;
  LAYER ME3 ;
  RECT 227.200 0.000 228.000 1.000 ;
  LAYER ME2 ;
  RECT 227.200 0.000 228.000 1.000 ;
  LAYER ME1 ;
  RECT 227.200 0.000 228.000 1.000 ;
 END
 ANTENNAPARTIALMETALAREA                  4.180 LAYER ME2 ;
 ANTENNADIFFAREA                          5.472 LAYER ME2 ;
 ANTENNADIFFAREA                          5.472 LAYER ME3 ;
 ANTENNADIFFAREA                          5.472 LAYER ME4 ;
END DO10
PIN DI10
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 212.800 0.000 213.600 1.000 ;
  LAYER ME3 ;
  RECT 212.800 0.000 213.600 1.000 ;
  LAYER ME2 ;
  RECT 212.800 0.000 213.600 1.000 ;
  LAYER ME1 ;
  RECT 212.800 0.000 213.600 1.000 ;
 END
 ANTENNAPARTIALMETALAREA                  3.122 LAYER ME2 ;
 ANTENNAGATEAREA                          0.086 LAYER ME2 ;
 ANTENNAGATEAREA                          0.086 LAYER ME3 ;
 ANTENNAGATEAREA                          0.086 LAYER ME4 ;
 ANTENNADIFFAREA                          0.160 LAYER ME2 ;
 ANTENNADIFFAREA                          0.160 LAYER ME3 ;
 ANTENNADIFFAREA                          0.160 LAYER ME4 ;
 ANTENNAMAXAREACAR                       48.477 LAYER ME2 ;
 ANTENNAMAXAREACAR                       57.736 LAYER ME3 ;
 ANTENNAMAXAREACAR                       66.995 LAYER ME4 ;
END DI10
PIN DO9
  DIRECTION OUTPUT ;
 PORT
  LAYER ME4 ;
  RECT 206.400 0.000 207.200 1.000 ;
  LAYER ME3 ;
  RECT 206.400 0.000 207.200 1.000 ;
  LAYER ME2 ;
  RECT 206.400 0.000 207.200 1.000 ;
  LAYER ME1 ;
  RECT 206.400 0.000 207.200 1.000 ;
 END
 ANTENNAPARTIALMETALAREA                  4.156 LAYER ME2 ;
 ANTENNADIFFAREA                          5.472 LAYER ME2 ;
 ANTENNADIFFAREA                          5.472 LAYER ME3 ;
 ANTENNADIFFAREA                          5.472 LAYER ME4 ;
END DO9
PIN DI9
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 191.600 0.000 192.400 1.000 ;
  LAYER ME3 ;
  RECT 191.600 0.000 192.400 1.000 ;
  LAYER ME2 ;
  RECT 191.600 0.000 192.400 1.000 ;
  LAYER ME1 ;
  RECT 191.600 0.000 192.400 1.000 ;
 END
 ANTENNAPARTIALMETALAREA                  3.134 LAYER ME2 ;
 ANTENNAGATEAREA                          0.086 LAYER ME2 ;
 ANTENNAGATEAREA                          0.086 LAYER ME3 ;
 ANTENNAGATEAREA                          0.086 LAYER ME4 ;
 ANTENNADIFFAREA                          0.160 LAYER ME2 ;
 ANTENNADIFFAREA                          0.160 LAYER ME3 ;
 ANTENNADIFFAREA                          0.160 LAYER ME4 ;
 ANTENNAMAXAREACAR                       48.616 LAYER ME2 ;
 ANTENNAMAXAREACAR                       57.875 LAYER ME3 ;
 ANTENNAMAXAREACAR                       67.134 LAYER ME4 ;
END DI9
PIN DO8
  DIRECTION OUTPUT ;
 PORT
  LAYER ME4 ;
  RECT 186.400 0.000 187.200 1.000 ;
  LAYER ME3 ;
  RECT 186.400 0.000 187.200 1.000 ;
  LAYER ME2 ;
  RECT 186.400 0.000 187.200 1.000 ;
  LAYER ME1 ;
  RECT 186.400 0.000 187.200 1.000 ;
 END
 ANTENNAPARTIALMETALAREA                  4.156 LAYER ME2 ;
 ANTENNADIFFAREA                          5.472 LAYER ME2 ;
 ANTENNADIFFAREA                          5.472 LAYER ME3 ;
 ANTENNADIFFAREA                          5.472 LAYER ME4 ;
END DO8
PIN WEB1
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 173.600 0.000 174.400 1.000 ;
  LAYER ME3 ;
  RECT 173.600 0.000 174.400 1.000 ;
  LAYER ME2 ;
  RECT 173.600 0.000 174.400 1.000 ;
  LAYER ME1 ;
  RECT 173.600 0.000 174.400 1.000 ;
 END
 ANTENNAPARTIALMETALAREA                  2.836 LAYER ME2 ;
 ANTENNAGATEAREA                          0.072 LAYER ME2 ;
 ANTENNAGATEAREA                          0.072 LAYER ME3 ;
 ANTENNAGATEAREA                          0.072 LAYER ME4 ;
 ANTENNADIFFAREA                          0.160 LAYER ME2 ;
 ANTENNADIFFAREA                          0.160 LAYER ME3 ;
 ANTENNADIFFAREA                          0.160 LAYER ME4 ;
 ANTENNAMAXAREACAR                       54.400 LAYER ME2 ;
 ANTENNAMAXAREACAR                       65.511 LAYER ME3 ;
 ANTENNAMAXAREACAR                       76.622 LAYER ME4 ;
END WEB1
PIN DI8
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 172.000 0.000 172.800 1.000 ;
  LAYER ME3 ;
  RECT 172.000 0.000 172.800 1.000 ;
  LAYER ME2 ;
  RECT 172.000 0.000 172.800 1.000 ;
  LAYER ME1 ;
  RECT 172.000 0.000 172.800 1.000 ;
 END
 ANTENNAPARTIALMETALAREA                  3.146 LAYER ME2 ;
 ANTENNAGATEAREA                          0.086 LAYER ME2 ;
 ANTENNAGATEAREA                          0.086 LAYER ME3 ;
 ANTENNAGATEAREA                          0.086 LAYER ME4 ;
 ANTENNADIFFAREA                          0.160 LAYER ME2 ;
 ANTENNADIFFAREA                          0.160 LAYER ME3 ;
 ANTENNADIFFAREA                          0.160 LAYER ME4 ;
 ANTENNAMAXAREACAR                       48.755 LAYER ME2 ;
 ANTENNAMAXAREACAR                       58.014 LAYER ME3 ;
 ANTENNAMAXAREACAR                       67.273 LAYER ME4 ;
END DI8
PIN DO7
  DIRECTION OUTPUT ;
 PORT
  LAYER ME4 ;
  RECT 165.200 0.000 166.000 1.000 ;
  LAYER ME3 ;
  RECT 165.200 0.000 166.000 1.000 ;
  LAYER ME2 ;
  RECT 165.200 0.000 166.000 1.000 ;
  LAYER ME1 ;
  RECT 165.200 0.000 166.000 1.000 ;
 END
 ANTENNAPARTIALMETALAREA                  4.180 LAYER ME2 ;
 ANTENNADIFFAREA                          5.472 LAYER ME2 ;
 ANTENNADIFFAREA                          5.472 LAYER ME3 ;
 ANTENNADIFFAREA                          5.472 LAYER ME4 ;
END DO7
PIN DI7
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 150.800 0.000 151.600 1.000 ;
  LAYER ME3 ;
  RECT 150.800 0.000 151.600 1.000 ;
  LAYER ME2 ;
  RECT 150.800 0.000 151.600 1.000 ;
  LAYER ME1 ;
  RECT 150.800 0.000 151.600 1.000 ;
 END
 ANTENNAPARTIALMETALAREA                  3.122 LAYER ME2 ;
 ANTENNAGATEAREA                          0.086 LAYER ME2 ;
 ANTENNAGATEAREA                          0.086 LAYER ME3 ;
 ANTENNAGATEAREA                          0.086 LAYER ME4 ;
 ANTENNADIFFAREA                          0.160 LAYER ME2 ;
 ANTENNADIFFAREA                          0.160 LAYER ME3 ;
 ANTENNADIFFAREA                          0.160 LAYER ME4 ;
 ANTENNAMAXAREACAR                       48.477 LAYER ME2 ;
 ANTENNAMAXAREACAR                       57.736 LAYER ME3 ;
 ANTENNAMAXAREACAR                       66.995 LAYER ME4 ;
END DI7
PIN DO6
  DIRECTION OUTPUT ;
 PORT
  LAYER ME4 ;
  RECT 145.600 0.000 146.400 1.000 ;
  LAYER ME3 ;
  RECT 145.600 0.000 146.400 1.000 ;
  LAYER ME2 ;
  RECT 145.600 0.000 146.400 1.000 ;
  LAYER ME1 ;
  RECT 145.600 0.000 146.400 1.000 ;
 END
 ANTENNAPARTIALMETALAREA                  4.148 LAYER ME2 ;
 ANTENNADIFFAREA                          5.472 LAYER ME2 ;
 ANTENNADIFFAREA                          5.472 LAYER ME3 ;
 ANTENNADIFFAREA                          5.472 LAYER ME4 ;
END DO6
PIN DI6
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 130.800 0.000 131.600 1.000 ;
  LAYER ME3 ;
  RECT 130.800 0.000 131.600 1.000 ;
  LAYER ME2 ;
  RECT 130.800 0.000 131.600 1.000 ;
  LAYER ME1 ;
  RECT 130.800 0.000 131.600 1.000 ;
 END
 ANTENNAPARTIALMETALAREA                  3.142 LAYER ME2 ;
 ANTENNAGATEAREA                          0.086 LAYER ME2 ;
 ANTENNAGATEAREA                          0.086 LAYER ME3 ;
 ANTENNAGATEAREA                          0.086 LAYER ME4 ;
 ANTENNADIFFAREA                          0.160 LAYER ME2 ;
 ANTENNADIFFAREA                          0.160 LAYER ME3 ;
 ANTENNADIFFAREA                          0.160 LAYER ME4 ;
 ANTENNAMAXAREACAR                       48.708 LAYER ME2 ;
 ANTENNAMAXAREACAR                       57.968 LAYER ME3 ;
 ANTENNAMAXAREACAR                       67.227 LAYER ME4 ;
END DI6
PIN DO5
  DIRECTION OUTPUT ;
 PORT
  LAYER ME4 ;
  RECT 124.400 0.000 125.200 1.000 ;
  LAYER ME3 ;
  RECT 124.400 0.000 125.200 1.000 ;
  LAYER ME2 ;
  RECT 124.400 0.000 125.200 1.000 ;
  LAYER ME1 ;
  RECT 124.400 0.000 125.200 1.000 ;
 END
 ANTENNAPARTIALMETALAREA                  4.156 LAYER ME2 ;
 ANTENNADIFFAREA                          5.472 LAYER ME2 ;
 ANTENNADIFFAREA                          5.472 LAYER ME3 ;
 ANTENNADIFFAREA                          5.472 LAYER ME4 ;
END DO5
PIN DI5
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 110.000 0.000 110.800 1.000 ;
  LAYER ME3 ;
  RECT 110.000 0.000 110.800 1.000 ;
  LAYER ME2 ;
  RECT 110.000 0.000 110.800 1.000 ;
  LAYER ME1 ;
  RECT 110.000 0.000 110.800 1.000 ;
 END
 ANTENNAPARTIALMETALAREA                  3.146 LAYER ME2 ;
 ANTENNAGATEAREA                          0.086 LAYER ME2 ;
 ANTENNAGATEAREA                          0.086 LAYER ME3 ;
 ANTENNAGATEAREA                          0.086 LAYER ME4 ;
 ANTENNADIFFAREA                          0.160 LAYER ME2 ;
 ANTENNADIFFAREA                          0.160 LAYER ME3 ;
 ANTENNADIFFAREA                          0.160 LAYER ME4 ;
 ANTENNAMAXAREACAR                       48.755 LAYER ME2 ;
 ANTENNAMAXAREACAR                       58.014 LAYER ME3 ;
 ANTENNAMAXAREACAR                       67.273 LAYER ME4 ;
END DI5
PIN DO4
  DIRECTION OUTPUT ;
 PORT
  LAYER ME4 ;
  RECT 104.800 0.000 105.600 1.000 ;
  LAYER ME3 ;
  RECT 104.800 0.000 105.600 1.000 ;
  LAYER ME2 ;
  RECT 104.800 0.000 105.600 1.000 ;
  LAYER ME1 ;
  RECT 104.800 0.000 105.600 1.000 ;
 END
 ANTENNAPARTIALMETALAREA                  4.172 LAYER ME2 ;
 ANTENNADIFFAREA                          5.472 LAYER ME2 ;
 ANTENNADIFFAREA                          5.472 LAYER ME3 ;
 ANTENNADIFFAREA                          5.472 LAYER ME4 ;
END DO4
PIN DI4
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 90.000 0.000 90.800 1.000 ;
  LAYER ME3 ;
  RECT 90.000 0.000 90.800 1.000 ;
  LAYER ME2 ;
  RECT 90.000 0.000 90.800 1.000 ;
  LAYER ME1 ;
  RECT 90.000 0.000 90.800 1.000 ;
 END
 ANTENNAPARTIALMETALAREA                  3.118 LAYER ME2 ;
 ANTENNAGATEAREA                          0.086 LAYER ME2 ;
 ANTENNAGATEAREA                          0.086 LAYER ME3 ;
 ANTENNAGATEAREA                          0.086 LAYER ME4 ;
 ANTENNADIFFAREA                          0.160 LAYER ME2 ;
 ANTENNADIFFAREA                          0.160 LAYER ME3 ;
 ANTENNADIFFAREA                          0.160 LAYER ME4 ;
 ANTENNAMAXAREACAR                       48.431 LAYER ME2 ;
 ANTENNAMAXAREACAR                       57.690 LAYER ME3 ;
 ANTENNAMAXAREACAR                       66.949 LAYER ME4 ;
END DI4
PIN DO3
  DIRECTION OUTPUT ;
 PORT
  LAYER ME4 ;
  RECT 83.600 0.000 84.400 1.000 ;
  LAYER ME3 ;
  RECT 83.600 0.000 84.400 1.000 ;
  LAYER ME2 ;
  RECT 83.600 0.000 84.400 1.000 ;
  LAYER ME1 ;
  RECT 83.600 0.000 84.400 1.000 ;
 END
 ANTENNAPARTIALMETALAREA                  4.148 LAYER ME2 ;
 ANTENNADIFFAREA                          5.472 LAYER ME2 ;
 ANTENNADIFFAREA                          5.472 LAYER ME3 ;
 ANTENNADIFFAREA                          5.472 LAYER ME4 ;
END DO3
PIN DI3
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 68.800 0.000 69.600 1.000 ;
  LAYER ME3 ;
  RECT 68.800 0.000 69.600 1.000 ;
  LAYER ME2 ;
  RECT 68.800 0.000 69.600 1.000 ;
  LAYER ME1 ;
  RECT 68.800 0.000 69.600 1.000 ;
 END
 ANTENNAPARTIALMETALAREA                  3.142 LAYER ME2 ;
 ANTENNAGATEAREA                          0.086 LAYER ME2 ;
 ANTENNAGATEAREA                          0.086 LAYER ME3 ;
 ANTENNAGATEAREA                          0.086 LAYER ME4 ;
 ANTENNADIFFAREA                          0.160 LAYER ME2 ;
 ANTENNADIFFAREA                          0.160 LAYER ME3 ;
 ANTENNADIFFAREA                          0.160 LAYER ME4 ;
 ANTENNAMAXAREACAR                       48.708 LAYER ME2 ;
 ANTENNAMAXAREACAR                       57.968 LAYER ME3 ;
 ANTENNAMAXAREACAR                       67.227 LAYER ME4 ;
END DI3
PIN DO2
  DIRECTION OUTPUT ;
 PORT
  LAYER ME4 ;
  RECT 63.600 0.000 64.400 1.000 ;
  LAYER ME3 ;
  RECT 63.600 0.000 64.400 1.000 ;
  LAYER ME2 ;
  RECT 63.600 0.000 64.400 1.000 ;
  LAYER ME1 ;
  RECT 63.600 0.000 64.400 1.000 ;
 END
 ANTENNAPARTIALMETALAREA                  4.164 LAYER ME2 ;
 ANTENNADIFFAREA                          5.472 LAYER ME2 ;
 ANTENNADIFFAREA                          5.472 LAYER ME3 ;
 ANTENNADIFFAREA                          5.472 LAYER ME4 ;
END DO2
PIN DI2
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 49.200 0.000 50.000 1.000 ;
  LAYER ME3 ;
  RECT 49.200 0.000 50.000 1.000 ;
  LAYER ME2 ;
  RECT 49.200 0.000 50.000 1.000 ;
  LAYER ME1 ;
  RECT 49.200 0.000 50.000 1.000 ;
 END
 ANTENNAPARTIALMETALAREA                  3.138 LAYER ME2 ;
 ANTENNAGATEAREA                          0.086 LAYER ME2 ;
 ANTENNAGATEAREA                          0.086 LAYER ME3 ;
 ANTENNAGATEAREA                          0.086 LAYER ME4 ;
 ANTENNADIFFAREA                          0.160 LAYER ME2 ;
 ANTENNADIFFAREA                          0.160 LAYER ME3 ;
 ANTENNADIFFAREA                          0.160 LAYER ME4 ;
 ANTENNAMAXAREACAR                       48.662 LAYER ME2 ;
 ANTENNAMAXAREACAR                       57.921 LAYER ME3 ;
 ANTENNAMAXAREACAR                       67.181 LAYER ME4 ;
END DI2
PIN DO1
  DIRECTION OUTPUT ;
 PORT
  LAYER ME4 ;
  RECT 42.800 0.000 43.600 1.000 ;
  LAYER ME3 ;
  RECT 42.800 0.000 43.600 1.000 ;
  LAYER ME2 ;
  RECT 42.800 0.000 43.600 1.000 ;
  LAYER ME1 ;
  RECT 42.800 0.000 43.600 1.000 ;
 END
 ANTENNAPARTIALMETALAREA                  4.172 LAYER ME2 ;
 ANTENNADIFFAREA                          5.472 LAYER ME2 ;
 ANTENNADIFFAREA                          5.472 LAYER ME3 ;
 ANTENNADIFFAREA                          5.472 LAYER ME4 ;
END DO1
PIN DI1
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 28.000 0.000 28.800 1.000 ;
  LAYER ME3 ;
  RECT 28.000 0.000 28.800 1.000 ;
  LAYER ME2 ;
  RECT 28.000 0.000 28.800 1.000 ;
  LAYER ME1 ;
  RECT 28.000 0.000 28.800 1.000 ;
 END
 ANTENNAPARTIALMETALAREA                  3.118 LAYER ME2 ;
 ANTENNAGATEAREA                          0.086 LAYER ME2 ;
 ANTENNAGATEAREA                          0.086 LAYER ME3 ;
 ANTENNAGATEAREA                          0.086 LAYER ME4 ;
 ANTENNADIFFAREA                          0.160 LAYER ME2 ;
 ANTENNADIFFAREA                          0.160 LAYER ME3 ;
 ANTENNADIFFAREA                          0.160 LAYER ME4 ;
 ANTENNAMAXAREACAR                       48.431 LAYER ME2 ;
 ANTENNAMAXAREACAR                       57.690 LAYER ME3 ;
 ANTENNAMAXAREACAR                       66.949 LAYER ME4 ;
END DI1
PIN DO0
  DIRECTION OUTPUT ;
 PORT
  LAYER ME4 ;
  RECT 22.800 0.000 23.600 1.000 ;
  LAYER ME3 ;
  RECT 22.800 0.000 23.600 1.000 ;
  LAYER ME2 ;
  RECT 22.800 0.000 23.600 1.000 ;
  LAYER ME1 ;
  RECT 22.800 0.000 23.600 1.000 ;
 END
 ANTENNAPARTIALMETALAREA                  4.140 LAYER ME2 ;
 ANTENNADIFFAREA                          5.472 LAYER ME2 ;
 ANTENNADIFFAREA                          5.472 LAYER ME3 ;
 ANTENNADIFFAREA                          5.472 LAYER ME4 ;
END DO0
PIN WEB0
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 10.000 0.000 10.800 1.000 ;
  LAYER ME3 ;
  RECT 10.000 0.000 10.800 1.000 ;
  LAYER ME2 ;
  RECT 10.000 0.000 10.800 1.000 ;
  LAYER ME1 ;
  RECT 10.000 0.000 10.800 1.000 ;
 END
 ANTENNAPARTIALMETALAREA                  2.852 LAYER ME2 ;
 ANTENNAGATEAREA                          0.072 LAYER ME2 ;
 ANTENNAGATEAREA                          0.072 LAYER ME3 ;
 ANTENNAGATEAREA                          0.072 LAYER ME4 ;
 ANTENNADIFFAREA                          0.160 LAYER ME2 ;
 ANTENNADIFFAREA                          0.160 LAYER ME3 ;
 ANTENNADIFFAREA                          0.160 LAYER ME4 ;
 ANTENNAMAXAREACAR                       54.622 LAYER ME2 ;
 ANTENNAMAXAREACAR                       65.733 LAYER ME3 ;
 ANTENNAMAXAREACAR                       76.844 LAYER ME4 ;
END WEB0
PIN DI0
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 8.000 0.000 8.800 1.000 ;
  LAYER ME3 ;
  RECT 8.000 0.000 8.800 1.000 ;
  LAYER ME2 ;
  RECT 8.000 0.000 8.800 1.000 ;
  LAYER ME1 ;
  RECT 8.000 0.000 8.800 1.000 ;
 END
 ANTENNAPARTIALMETALAREA                  3.150 LAYER ME2 ;
 ANTENNAGATEAREA                          0.086 LAYER ME2 ;
 ANTENNAGATEAREA                          0.086 LAYER ME3 ;
 ANTENNAGATEAREA                          0.086 LAYER ME4 ;
 ANTENNADIFFAREA                          0.160 LAYER ME2 ;
 ANTENNADIFFAREA                          0.160 LAYER ME3 ;
 ANTENNADIFFAREA                          0.160 LAYER ME4 ;
 ANTENNAMAXAREACAR                       48.801 LAYER ME2 ;
 ANTENNAMAXAREACAR                       58.060 LAYER ME3 ;
 ANTENNAMAXAREACAR                       67.319 LAYER ME4 ;
END DI0
PIN VCC
  DIRECTION INOUT ;
  USE POWER ;
  SHAPE RING ;
 PORT
  LAYER ME4 ;
  RECT 2.000 561.930 2690.940 563.930 ;
  RECT 2.000 3.600 2690.940 5.600 ;
  RECT 2688.940 3.600 2690.940 563.930 ;
  RECT 2.000 3.600 4.000 563.930 ;
 END
END VCC
PIN GND
  DIRECTION INOUT ;
  USE GROUND ;
  SHAPE RING ;
 PORT
  LAYER ME3 ;
  RECT 0.000 563.930 2692.940 565.930 ;
  RECT 0.000 1.600 2692.940 3.600 ;
  RECT 2690.940 1.600 2692.940 565.930 ;
  RECT 0.000 1.600 2.000 565.930 ;
 END
END GND
OBS
  LAYER ME4 ;
  RECT 5.420 7.020 2687.520 560.510 ;
  RECT 2688.940 5.600 2690.940 561.930 ;
  RECT 2.000 5.600 4.000 561.930 ;
  RECT 4.000 561.930 2688.940 563.930 ;
  RECT 4.000 3.600 2688.940 5.600 ;
  RECT 2.000 561.930 4.000 563.930 ;
  RECT 2688.940 3.600 2690.940 5.600 ;
  RECT 2688.940 561.930 2690.940 563.930 ;
  RECT 2.000 3.600 4.000 5.600 ;
  RECT 2680.800 0.000 2681.600 1.000 ;
  RECT 2666.400 0.000 2667.200 1.000 ;
  RECT 2661.200 0.000 2662.000 1.000 ;
  RECT 2646.400 0.000 2647.200 1.000 ;
  RECT 2640.000 0.000 2640.800 1.000 ;
  RECT 2625.600 0.000 2626.400 1.000 ;
  RECT 2620.400 0.000 2621.200 1.000 ;
  RECT 2605.600 0.000 2606.400 1.000 ;
  RECT 2599.200 0.000 2600.000 1.000 ;
  RECT 2584.400 0.000 2585.200 1.000 ;
  RECT 2579.200 0.000 2580.000 1.000 ;
  RECT 2564.800 0.000 2565.600 1.000 ;
  RECT 2558.400 0.000 2559.200 1.000 ;
  RECT 2543.600 0.000 2544.400 1.000 ;
  RECT 2538.400 0.000 2539.200 1.000 ;
  RECT 2525.600 0.000 2526.400 1.000 ;
  RECT 2523.600 0.000 2524.400 1.000 ;
  RECT 2517.200 0.000 2518.000 1.000 ;
  RECT 2502.800 0.000 2503.600 1.000 ;
  RECT 2497.600 0.000 2498.400 1.000 ;
  RECT 2482.800 0.000 2483.600 1.000 ;
  RECT 2476.400 0.000 2477.200 1.000 ;
  RECT 2461.600 0.000 2462.400 1.000 ;
  RECT 2456.400 0.000 2457.200 1.000 ;
  RECT 2442.000 0.000 2442.800 1.000 ;
  RECT 2435.600 0.000 2436.400 1.000 ;
  RECT 2420.800 0.000 2421.600 1.000 ;
  RECT 2415.600 0.000 2416.400 1.000 ;
  RECT 2400.800 0.000 2401.600 1.000 ;
  RECT 2394.400 0.000 2395.200 1.000 ;
  RECT 2380.000 0.000 2380.800 1.000 ;
  RECT 2374.800 0.000 2375.600 1.000 ;
  RECT 2361.600 0.000 2362.400 1.000 ;
  RECT 2360.000 0.000 2360.800 1.000 ;
  RECT 2353.600 0.000 2354.400 1.000 ;
  RECT 2338.800 0.000 2339.600 1.000 ;
  RECT 2333.600 0.000 2334.400 1.000 ;
  RECT 2319.200 0.000 2320.000 1.000 ;
  RECT 2312.800 0.000 2313.600 1.000 ;
  RECT 2298.000 0.000 2298.800 1.000 ;
  RECT 2292.800 0.000 2293.600 1.000 ;
  RECT 2278.400 0.000 2279.200 1.000 ;
  RECT 2271.600 0.000 2272.400 1.000 ;
  RECT 2257.200 0.000 2258.000 1.000 ;
  RECT 2252.000 0.000 2252.800 1.000 ;
  RECT 2237.200 0.000 2238.000 1.000 ;
  RECT 2230.800 0.000 2231.600 1.000 ;
  RECT 2216.400 0.000 2217.200 1.000 ;
  RECT 2211.200 0.000 2212.000 1.000 ;
  RECT 2198.000 0.000 2198.800 1.000 ;
  RECT 2196.400 0.000 2197.200 1.000 ;
  RECT 2190.000 0.000 2190.800 1.000 ;
  RECT 2175.200 0.000 2176.000 1.000 ;
  RECT 2170.000 0.000 2170.800 1.000 ;
  RECT 2155.600 0.000 2156.400 1.000 ;
  RECT 2149.200 0.000 2150.000 1.000 ;
  RECT 2134.400 0.000 2135.200 1.000 ;
  RECT 2129.200 0.000 2130.000 1.000 ;
  RECT 2114.400 0.000 2115.200 1.000 ;
  RECT 2108.000 0.000 2108.800 1.000 ;
  RECT 2093.600 0.000 2094.400 1.000 ;
  RECT 2088.400 0.000 2089.200 1.000 ;
  RECT 2073.600 0.000 2074.400 1.000 ;
  RECT 2067.200 0.000 2068.000 1.000 ;
  RECT 2052.400 0.000 2053.200 1.000 ;
  RECT 2047.200 0.000 2048.000 1.000 ;
  RECT 2034.400 0.000 2035.200 1.000 ;
  RECT 2032.800 0.000 2033.600 1.000 ;
  RECT 2026.400 0.000 2027.200 1.000 ;
  RECT 2011.600 0.000 2012.400 1.000 ;
  RECT 2006.400 0.000 2007.200 1.000 ;
  RECT 1991.600 0.000 1992.400 1.000 ;
  RECT 1985.200 0.000 1986.000 1.000 ;
  RECT 1970.800 0.000 1971.600 1.000 ;
  RECT 1965.600 0.000 1966.400 1.000 ;
  RECT 1950.800 0.000 1951.600 1.000 ;
  RECT 1944.400 0.000 1945.200 1.000 ;
  RECT 1929.600 0.000 1930.400 1.000 ;
  RECT 1924.400 0.000 1925.200 1.000 ;
  RECT 1910.000 0.000 1910.800 1.000 ;
  RECT 1903.600 0.000 1904.400 1.000 ;
  RECT 1888.800 0.000 1889.600 1.000 ;
  RECT 1883.600 0.000 1884.400 1.000 ;
  RECT 1870.800 0.000 1871.600 1.000 ;
  RECT 1869.200 0.000 1870.000 1.000 ;
  RECT 1862.400 0.000 1863.200 1.000 ;
  RECT 1848.000 0.000 1848.800 1.000 ;
  RECT 1842.800 0.000 1843.600 1.000 ;
  RECT 1828.000 0.000 1828.800 1.000 ;
  RECT 1821.600 0.000 1822.400 1.000 ;
  RECT 1807.200 0.000 1808.000 1.000 ;
  RECT 1802.000 0.000 1802.800 1.000 ;
  RECT 1787.200 0.000 1788.000 1.000 ;
  RECT 1780.800 0.000 1781.600 1.000 ;
  RECT 1766.000 0.000 1766.800 1.000 ;
  RECT 1760.800 0.000 1761.600 1.000 ;
  RECT 1746.400 0.000 1747.200 1.000 ;
  RECT 1740.000 0.000 1740.800 1.000 ;
  RECT 1725.200 0.000 1726.000 1.000 ;
  RECT 1720.000 0.000 1720.800 1.000 ;
  RECT 1707.200 0.000 1708.000 1.000 ;
  RECT 1705.200 0.000 1706.000 1.000 ;
  RECT 1698.800 0.000 1699.600 1.000 ;
  RECT 1684.400 0.000 1685.200 1.000 ;
  RECT 1679.200 0.000 1680.000 1.000 ;
  RECT 1664.400 0.000 1665.200 1.000 ;
  RECT 1658.000 0.000 1658.800 1.000 ;
  RECT 1643.200 0.000 1644.000 1.000 ;
  RECT 1638.000 0.000 1638.800 1.000 ;
  RECT 1623.600 0.000 1624.400 1.000 ;
  RECT 1617.200 0.000 1618.000 1.000 ;
  RECT 1602.400 0.000 1603.200 1.000 ;
  RECT 1597.200 0.000 1598.000 1.000 ;
  RECT 1582.400 0.000 1583.200 1.000 ;
  RECT 1576.000 0.000 1576.800 1.000 ;
  RECT 1561.600 0.000 1562.400 1.000 ;
  RECT 1556.400 0.000 1557.200 1.000 ;
  RECT 1543.200 0.000 1544.000 1.000 ;
  RECT 1541.600 0.000 1542.400 1.000 ;
  RECT 1535.200 0.000 1536.000 1.000 ;
  RECT 1520.400 0.000 1521.200 1.000 ;
  RECT 1515.200 0.000 1516.000 1.000 ;
  RECT 1500.800 0.000 1501.600 1.000 ;
  RECT 1494.400 0.000 1495.200 1.000 ;
  RECT 1479.600 0.000 1480.400 1.000 ;
  RECT 1474.400 0.000 1475.200 1.000 ;
  RECT 1460.000 0.000 1460.800 1.000 ;
  RECT 1453.200 0.000 1454.000 1.000 ;
  RECT 1438.800 0.000 1439.600 1.000 ;
  RECT 1433.600 0.000 1434.400 1.000 ;
  RECT 1418.800 0.000 1419.600 1.000 ;
  RECT 1412.400 0.000 1413.200 1.000 ;
  RECT 1398.000 0.000 1398.800 1.000 ;
  RECT 1392.800 0.000 1393.600 1.000 ;
  RECT 1379.600 0.000 1380.400 1.000 ;
  RECT 1378.000 0.000 1378.800 1.000 ;
  RECT 1357.200 0.000 1358.000 1.000 ;
  RECT 1356.000 0.000 1356.800 1.000 ;
  RECT 1354.800 0.000 1355.600 1.000 ;
  RECT 1353.600 0.000 1354.400 1.000 ;
  RECT 1352.400 0.000 1353.200 1.000 ;
  RECT 1351.200 0.000 1352.000 1.000 ;
  RECT 1345.200 0.000 1346.000 1.000 ;
  RECT 1338.000 0.000 1338.800 1.000 ;
  RECT 1335.200 0.000 1336.000 1.000 ;
  RECT 1332.400 0.000 1333.200 1.000 ;
  RECT 1330.000 0.000 1330.800 1.000 ;
  RECT 1328.400 0.000 1329.200 1.000 ;
  RECT 1326.000 0.000 1326.800 1.000 ;
  RECT 1324.400 0.000 1325.200 1.000 ;
  RECT 1322.000 0.000 1322.800 1.000 ;
  RECT 1320.400 0.000 1321.200 1.000 ;
  RECT 1311.200 0.000 1312.000 1.000 ;
  RECT 1296.400 0.000 1297.200 1.000 ;
  RECT 1291.200 0.000 1292.000 1.000 ;
  RECT 1276.800 0.000 1277.600 1.000 ;
  RECT 1270.400 0.000 1271.200 1.000 ;
  RECT 1255.600 0.000 1256.400 1.000 ;
  RECT 1250.400 0.000 1251.200 1.000 ;
  RECT 1235.600 0.000 1236.400 1.000 ;
  RECT 1229.200 0.000 1230.000 1.000 ;
  RECT 1214.800 0.000 1215.600 1.000 ;
  RECT 1209.600 0.000 1210.400 1.000 ;
  RECT 1194.800 0.000 1195.600 1.000 ;
  RECT 1188.400 0.000 1189.200 1.000 ;
  RECT 1173.600 0.000 1174.400 1.000 ;
  RECT 1168.400 0.000 1169.200 1.000 ;
  RECT 1155.600 0.000 1156.400 1.000 ;
  RECT 1154.000 0.000 1154.800 1.000 ;
  RECT 1147.600 0.000 1148.400 1.000 ;
  RECT 1132.800 0.000 1133.600 1.000 ;
  RECT 1127.600 0.000 1128.400 1.000 ;
  RECT 1113.200 0.000 1114.000 1.000 ;
  RECT 1106.400 0.000 1107.200 1.000 ;
  RECT 1092.000 0.000 1092.800 1.000 ;
  RECT 1086.800 0.000 1087.600 1.000 ;
  RECT 1072.000 0.000 1072.800 1.000 ;
  RECT 1065.600 0.000 1066.400 1.000 ;
  RECT 1051.200 0.000 1052.000 1.000 ;
  RECT 1045.600 0.000 1046.400 1.000 ;
  RECT 1031.200 0.000 1032.000 1.000 ;
  RECT 1024.800 0.000 1025.600 1.000 ;
  RECT 1010.000 0.000 1010.800 1.000 ;
  RECT 1004.800 0.000 1005.600 1.000 ;
  RECT 992.000 0.000 992.800 1.000 ;
  RECT 990.400 0.000 991.200 1.000 ;
  RECT 983.600 0.000 984.400 1.000 ;
  RECT 969.200 0.000 970.000 1.000 ;
  RECT 964.000 0.000 964.800 1.000 ;
  RECT 949.200 0.000 950.000 1.000 ;
  RECT 942.800 0.000 943.600 1.000 ;
  RECT 928.400 0.000 929.200 1.000 ;
  RECT 923.200 0.000 924.000 1.000 ;
  RECT 908.400 0.000 909.200 1.000 ;
  RECT 902.000 0.000 902.800 1.000 ;
  RECT 887.200 0.000 888.000 1.000 ;
  RECT 882.000 0.000 882.800 1.000 ;
  RECT 867.600 0.000 868.400 1.000 ;
  RECT 861.200 0.000 862.000 1.000 ;
  RECT 846.400 0.000 847.200 1.000 ;
  RECT 841.200 0.000 842.000 1.000 ;
  RECT 828.400 0.000 829.200 1.000 ;
  RECT 826.400 0.000 827.200 1.000 ;
  RECT 820.000 0.000 820.800 1.000 ;
  RECT 805.600 0.000 806.400 1.000 ;
  RECT 800.400 0.000 801.200 1.000 ;
  RECT 785.600 0.000 786.400 1.000 ;
  RECT 779.200 0.000 780.000 1.000 ;
  RECT 764.400 0.000 765.200 1.000 ;
  RECT 759.200 0.000 760.000 1.000 ;
  RECT 744.800 0.000 745.600 1.000 ;
  RECT 738.400 0.000 739.200 1.000 ;
  RECT 723.600 0.000 724.400 1.000 ;
  RECT 718.400 0.000 719.200 1.000 ;
  RECT 704.000 0.000 704.800 1.000 ;
  RECT 697.200 0.000 698.000 1.000 ;
  RECT 682.800 0.000 683.600 1.000 ;
  RECT 677.600 0.000 678.400 1.000 ;
  RECT 664.800 0.000 665.600 1.000 ;
  RECT 662.800 0.000 663.600 1.000 ;
  RECT 656.400 0.000 657.200 1.000 ;
  RECT 642.000 0.000 642.800 1.000 ;
  RECT 636.400 0.000 637.200 1.000 ;
  RECT 622.000 0.000 622.800 1.000 ;
  RECT 615.600 0.000 616.400 1.000 ;
  RECT 600.800 0.000 601.600 1.000 ;
  RECT 595.600 0.000 596.400 1.000 ;
  RECT 581.200 0.000 582.000 1.000 ;
  RECT 574.400 0.000 575.200 1.000 ;
  RECT 560.000 0.000 560.800 1.000 ;
  RECT 554.800 0.000 555.600 1.000 ;
  RECT 540.000 0.000 540.800 1.000 ;
  RECT 533.600 0.000 534.400 1.000 ;
  RECT 519.200 0.000 520.000 1.000 ;
  RECT 514.000 0.000 514.800 1.000 ;
  RECT 500.800 0.000 501.600 1.000 ;
  RECT 499.200 0.000 500.000 1.000 ;
  RECT 492.800 0.000 493.600 1.000 ;
  RECT 478.000 0.000 478.800 1.000 ;
  RECT 472.800 0.000 473.600 1.000 ;
  RECT 458.400 0.000 459.200 1.000 ;
  RECT 452.000 0.000 452.800 1.000 ;
  RECT 437.200 0.000 438.000 1.000 ;
  RECT 432.000 0.000 432.800 1.000 ;
  RECT 417.200 0.000 418.000 1.000 ;
  RECT 410.800 0.000 411.600 1.000 ;
  RECT 396.400 0.000 397.200 1.000 ;
  RECT 391.200 0.000 392.000 1.000 ;
  RECT 376.400 0.000 377.200 1.000 ;
  RECT 370.000 0.000 370.800 1.000 ;
  RECT 355.200 0.000 356.000 1.000 ;
  RECT 350.000 0.000 350.800 1.000 ;
  RECT 337.200 0.000 338.000 1.000 ;
  RECT 335.600 0.000 336.400 1.000 ;
  RECT 329.200 0.000 330.000 1.000 ;
  RECT 314.400 0.000 315.200 1.000 ;
  RECT 309.200 0.000 310.000 1.000 ;
  RECT 294.800 0.000 295.600 1.000 ;
  RECT 288.000 0.000 288.800 1.000 ;
  RECT 273.600 0.000 274.400 1.000 ;
  RECT 268.400 0.000 269.200 1.000 ;
  RECT 253.600 0.000 254.400 1.000 ;
  RECT 247.200 0.000 248.000 1.000 ;
  RECT 232.800 0.000 233.600 1.000 ;
  RECT 227.200 0.000 228.000 1.000 ;
  RECT 212.800 0.000 213.600 1.000 ;
  RECT 206.400 0.000 207.200 1.000 ;
  RECT 191.600 0.000 192.400 1.000 ;
  RECT 186.400 0.000 187.200 1.000 ;
  RECT 173.600 0.000 174.400 1.000 ;
  RECT 172.000 0.000 172.800 1.000 ;
  RECT 165.200 0.000 166.000 1.000 ;
  RECT 150.800 0.000 151.600 1.000 ;
  RECT 145.600 0.000 146.400 1.000 ;
  RECT 130.800 0.000 131.600 1.000 ;
  RECT 124.400 0.000 125.200 1.000 ;
  RECT 110.000 0.000 110.800 1.000 ;
  RECT 104.800 0.000 105.600 1.000 ;
  RECT 90.000 0.000 90.800 1.000 ;
  RECT 83.600 0.000 84.400 1.000 ;
  RECT 68.800 0.000 69.600 1.000 ;
  RECT 63.600 0.000 64.400 1.000 ;
  RECT 49.200 0.000 50.000 1.000 ;
  RECT 42.800 0.000 43.600 1.000 ;
  RECT 28.000 0.000 28.800 1.000 ;
  RECT 22.800 0.000 23.600 1.000 ;
  RECT 10.000 0.000 10.800 1.000 ;
  RECT 8.000 0.000 8.800 1.000 ;
  RECT 2687.800 9.570 2688.940 11.170 ;
  RECT 2687.800 14.200 2688.940 15.200 ;
  RECT 2687.800 18.730 2688.940 19.730 ;
  RECT 2687.800 21.230 2688.940 22.070 ;
  RECT 2687.800 24.170 2688.940 25.170 ;
  RECT 2687.800 36.320 2688.940 37.320 ;
  RECT 2687.800 39.480 2688.940 40.080 ;
  RECT 2687.800 45.560 2688.940 46.160 ;
  RECT 2687.800 57.100 2688.940 61.420 ;
  RECT 2686.380 5.880 2687.520 7.020 ;
  RECT 1388.220 5.600 1396.220 7.020 ;
  RECT 1378.180 5.880 1386.180 7.020 ;
  RECT 1398.020 5.880 1406.020 7.020 ;
  RECT 1408.060 5.600 1416.060 7.020 ;
  RECT 1419.100 5.880 1427.100 7.020 ;
  RECT 1429.140 5.600 1437.140 7.020 ;
  RECT 1438.940 5.880 1446.940 7.020 ;
  RECT 1448.980 5.600 1456.980 7.020 ;
  RECT 1460.020 5.880 1468.020 7.020 ;
  RECT 1470.060 5.600 1478.060 7.020 ;
  RECT 1479.860 5.880 1487.860 7.020 ;
  RECT 1489.900 5.600 1497.900 7.020 ;
  RECT 1500.940 5.880 1508.940 7.020 ;
  RECT 1510.980 5.600 1518.980 7.020 ;
  RECT 1520.780 5.880 1528.780 7.020 ;
  RECT 1530.820 5.600 1538.820 7.020 ;
  RECT 1551.900 5.600 1559.900 7.020 ;
  RECT 1541.860 5.880 1549.860 7.020 ;
  RECT 1561.700 5.880 1569.700 7.020 ;
  RECT 1571.740 5.600 1579.740 7.020 ;
  RECT 1582.780 5.880 1590.780 7.020 ;
  RECT 1592.820 5.600 1600.820 7.020 ;
  RECT 1602.620 5.880 1610.620 7.020 ;
  RECT 1612.660 5.600 1620.660 7.020 ;
  RECT 1623.700 5.880 1631.700 7.020 ;
  RECT 1633.740 5.600 1641.740 7.020 ;
  RECT 1643.540 5.880 1651.540 7.020 ;
  RECT 1653.580 5.600 1661.580 7.020 ;
  RECT 1664.620 5.880 1672.620 7.020 ;
  RECT 1674.660 5.600 1682.660 7.020 ;
  RECT 1684.460 5.880 1692.460 7.020 ;
  RECT 1694.500 5.600 1702.500 7.020 ;
  RECT 1715.580 5.600 1723.580 7.020 ;
  RECT 1705.540 5.880 1713.540 7.020 ;
  RECT 1725.380 5.880 1733.380 7.020 ;
  RECT 1735.420 5.600 1743.420 7.020 ;
  RECT 1746.460 5.880 1754.460 7.020 ;
  RECT 1756.500 5.600 1764.500 7.020 ;
  RECT 1766.300 5.880 1774.300 7.020 ;
  RECT 1776.340 5.600 1784.340 7.020 ;
  RECT 1787.380 5.880 1795.380 7.020 ;
  RECT 1797.420 5.600 1805.420 7.020 ;
  RECT 1807.220 5.880 1815.220 7.020 ;
  RECT 1817.260 5.600 1825.260 7.020 ;
  RECT 1828.300 5.880 1836.300 7.020 ;
  RECT 1838.340 5.600 1846.340 7.020 ;
  RECT 1848.140 5.880 1856.140 7.020 ;
  RECT 1858.180 5.600 1866.180 7.020 ;
  RECT 1879.260 5.600 1887.260 7.020 ;
  RECT 1869.220 5.880 1877.220 7.020 ;
  RECT 1889.060 5.880 1897.060 7.020 ;
  RECT 1899.100 5.600 1907.100 7.020 ;
  RECT 1910.140 5.880 1918.140 7.020 ;
  RECT 1920.180 5.600 1928.180 7.020 ;
  RECT 1929.980 5.880 1937.980 7.020 ;
  RECT 1940.020 5.600 1948.020 7.020 ;
  RECT 1951.060 5.880 1959.060 7.020 ;
  RECT 1961.100 5.600 1969.100 7.020 ;
  RECT 1970.900 5.880 1978.900 7.020 ;
  RECT 1980.940 5.600 1988.940 7.020 ;
  RECT 1991.980 5.880 1999.980 7.020 ;
  RECT 2002.020 5.600 2010.020 7.020 ;
  RECT 2011.820 5.880 2019.820 7.020 ;
  RECT 2021.860 5.600 2029.860 7.020 ;
  RECT 2042.940 5.600 2050.940 7.020 ;
  RECT 2032.900 5.880 2040.900 7.020 ;
  RECT 2052.740 5.880 2060.740 7.020 ;
  RECT 2062.780 5.600 2070.780 7.020 ;
  RECT 2073.820 5.880 2081.820 7.020 ;
  RECT 2083.860 5.600 2091.860 7.020 ;
  RECT 2093.660 5.880 2101.660 7.020 ;
  RECT 2103.700 5.600 2111.700 7.020 ;
  RECT 2114.740 5.880 2122.740 7.020 ;
  RECT 2124.780 5.600 2132.780 7.020 ;
  RECT 2134.580 5.880 2142.580 7.020 ;
  RECT 2144.620 5.600 2152.620 7.020 ;
  RECT 2155.660 5.880 2163.660 7.020 ;
  RECT 2165.700 5.600 2173.700 7.020 ;
  RECT 2175.500 5.880 2183.500 7.020 ;
  RECT 2185.540 5.600 2193.540 7.020 ;
  RECT 2206.620 5.600 2214.620 7.020 ;
  RECT 2196.580 5.880 2204.580 7.020 ;
  RECT 2216.420 5.880 2224.420 7.020 ;
  RECT 2226.460 5.600 2234.460 7.020 ;
  RECT 2237.500 5.880 2245.500 7.020 ;
  RECT 2247.540 5.600 2255.540 7.020 ;
  RECT 2257.340 5.880 2265.340 7.020 ;
  RECT 2267.380 5.600 2275.380 7.020 ;
  RECT 2278.420 5.880 2286.420 7.020 ;
  RECT 2288.460 5.600 2296.460 7.020 ;
  RECT 2298.260 5.880 2306.260 7.020 ;
  RECT 2308.300 5.600 2316.300 7.020 ;
  RECT 2319.340 5.880 2327.340 7.020 ;
  RECT 2329.380 5.600 2337.380 7.020 ;
  RECT 2339.180 5.880 2347.180 7.020 ;
  RECT 2349.220 5.600 2357.220 7.020 ;
  RECT 2370.300 5.600 2378.300 7.020 ;
  RECT 2360.260 5.880 2368.260 7.020 ;
  RECT 2380.100 5.880 2388.100 7.020 ;
  RECT 2390.140 5.600 2398.140 7.020 ;
  RECT 2401.180 5.880 2409.180 7.020 ;
  RECT 2411.220 5.600 2419.220 7.020 ;
  RECT 2421.020 5.880 2429.020 7.020 ;
  RECT 2431.060 5.600 2439.060 7.020 ;
  RECT 2442.100 5.880 2450.100 7.020 ;
  RECT 2452.140 5.600 2460.140 7.020 ;
  RECT 2461.940 5.880 2469.940 7.020 ;
  RECT 2471.980 5.600 2479.980 7.020 ;
  RECT 2483.020 5.880 2491.020 7.020 ;
  RECT 2493.060 5.600 2501.060 7.020 ;
  RECT 2502.860 5.880 2510.860 7.020 ;
  RECT 2512.900 5.600 2520.900 7.020 ;
  RECT 2533.980 5.600 2541.980 7.020 ;
  RECT 2523.940 5.880 2531.940 7.020 ;
  RECT 2543.780 5.880 2551.780 7.020 ;
  RECT 2553.820 5.600 2561.820 7.020 ;
  RECT 2564.860 5.880 2572.860 7.020 ;
  RECT 2574.900 5.600 2582.900 7.020 ;
  RECT 2584.700 5.880 2592.700 7.020 ;
  RECT 2594.740 5.600 2602.740 7.020 ;
  RECT 2605.780 5.880 2613.780 7.020 ;
  RECT 2615.820 5.600 2623.820 7.020 ;
  RECT 2625.620 5.880 2633.620 7.020 ;
  RECT 2635.660 5.600 2643.660 7.020 ;
  RECT 2646.700 5.880 2654.700 7.020 ;
  RECT 2656.740 5.600 2664.740 7.020 ;
  RECT 2666.540 5.880 2674.540 7.020 ;
  RECT 2676.580 5.600 2684.580 7.020 ;
  RECT 1339.880 5.600 1342.940 7.020 ;
  RECT 1343.440 5.880 1346.890 7.020 ;
  RECT 1347.390 5.600 1351.140 7.020 ;
  RECT 1352.290 5.880 1358.210 7.020 ;
  RECT 1359.360 5.600 1363.110 7.020 ;
  RECT 1363.610 5.600 1367.360 7.020 ;
  RECT 1367.860 5.600 1371.610 7.020 ;
  RECT 1337.160 5.600 1338.920 7.020 ;
  RECT 1335.160 5.880 1336.920 7.020 ;
  RECT 1331.820 5.600 1333.580 7.020 ;
  RECT 1329.820 5.880 1331.580 7.020 ;
  RECT 1327.820 5.600 1329.580 7.020 ;
  RECT 1325.820 5.880 1327.580 7.020 ;
  RECT 1323.820 5.600 1325.580 7.020 ;
  RECT 1321.820 5.880 1323.580 7.020 ;
  RECT 1319.820 5.600 1321.580 7.020 ;
  RECT 1317.820 5.880 1319.580 7.020 ;
  RECT 4.000 57.100 5.140 61.420 ;
  RECT 4.000 45.560 5.140 46.160 ;
  RECT 4.000 39.480 5.140 40.080 ;
  RECT 4.000 36.320 5.140 37.320 ;
  RECT 4.000 24.170 5.140 25.170 ;
  RECT 4.000 21.230 5.140 22.070 ;
  RECT 4.000 18.730 5.140 19.730 ;
  RECT 4.000 14.200 5.140 15.200 ;
  RECT 4.000 9.570 5.140 11.170 ;
  RECT 5.420 5.880 6.560 7.020 ;
  RECT 18.400 5.600 26.400 7.020 ;
  RECT 8.360 5.880 16.360 7.020 ;
  RECT 28.200 5.880 36.200 7.020 ;
  RECT 38.240 5.600 46.240 7.020 ;
  RECT 49.280 5.880 57.280 7.020 ;
  RECT 59.320 5.600 67.320 7.020 ;
  RECT 69.120 5.880 77.120 7.020 ;
  RECT 79.160 5.600 87.160 7.020 ;
  RECT 90.200 5.880 98.200 7.020 ;
  RECT 100.240 5.600 108.240 7.020 ;
  RECT 110.040 5.880 118.040 7.020 ;
  RECT 120.080 5.600 128.080 7.020 ;
  RECT 131.120 5.880 139.120 7.020 ;
  RECT 141.160 5.600 149.160 7.020 ;
  RECT 150.960 5.880 158.960 7.020 ;
  RECT 161.000 5.600 169.000 7.020 ;
  RECT 182.080 5.600 190.080 7.020 ;
  RECT 172.040 5.880 180.040 7.020 ;
  RECT 191.880 5.880 199.880 7.020 ;
  RECT 201.920 5.600 209.920 7.020 ;
  RECT 212.960 5.880 220.960 7.020 ;
  RECT 223.000 5.600 231.000 7.020 ;
  RECT 232.800 5.880 240.800 7.020 ;
  RECT 242.840 5.600 250.840 7.020 ;
  RECT 253.880 5.880 261.880 7.020 ;
  RECT 263.920 5.600 271.920 7.020 ;
  RECT 273.720 5.880 281.720 7.020 ;
  RECT 283.760 5.600 291.760 7.020 ;
  RECT 294.800 5.880 302.800 7.020 ;
  RECT 304.840 5.600 312.840 7.020 ;
  RECT 314.640 5.880 322.640 7.020 ;
  RECT 324.680 5.600 332.680 7.020 ;
  RECT 345.760 5.600 353.760 7.020 ;
  RECT 335.720 5.880 343.720 7.020 ;
  RECT 355.560 5.880 363.560 7.020 ;
  RECT 365.600 5.600 373.600 7.020 ;
  RECT 376.640 5.880 384.640 7.020 ;
  RECT 386.680 5.600 394.680 7.020 ;
  RECT 396.480 5.880 404.480 7.020 ;
  RECT 406.520 5.600 414.520 7.020 ;
  RECT 417.560 5.880 425.560 7.020 ;
  RECT 427.600 5.600 435.600 7.020 ;
  RECT 437.400 5.880 445.400 7.020 ;
  RECT 447.440 5.600 455.440 7.020 ;
  RECT 458.480 5.880 466.480 7.020 ;
  RECT 468.520 5.600 476.520 7.020 ;
  RECT 478.320 5.880 486.320 7.020 ;
  RECT 488.360 5.600 496.360 7.020 ;
  RECT 509.440 5.600 517.440 7.020 ;
  RECT 499.400 5.880 507.400 7.020 ;
  RECT 519.240 5.880 527.240 7.020 ;
  RECT 529.280 5.600 537.280 7.020 ;
  RECT 540.320 5.880 548.320 7.020 ;
  RECT 550.360 5.600 558.360 7.020 ;
  RECT 560.160 5.880 568.160 7.020 ;
  RECT 570.200 5.600 578.200 7.020 ;
  RECT 581.240 5.880 589.240 7.020 ;
  RECT 591.280 5.600 599.280 7.020 ;
  RECT 601.080 5.880 609.080 7.020 ;
  RECT 611.120 5.600 619.120 7.020 ;
  RECT 622.160 5.880 630.160 7.020 ;
  RECT 632.200 5.600 640.200 7.020 ;
  RECT 642.000 5.880 650.000 7.020 ;
  RECT 652.040 5.600 660.040 7.020 ;
  RECT 673.120 5.600 681.120 7.020 ;
  RECT 663.080 5.880 671.080 7.020 ;
  RECT 682.920 5.880 690.920 7.020 ;
  RECT 692.960 5.600 700.960 7.020 ;
  RECT 704.000 5.880 712.000 7.020 ;
  RECT 714.040 5.600 722.040 7.020 ;
  RECT 723.840 5.880 731.840 7.020 ;
  RECT 733.880 5.600 741.880 7.020 ;
  RECT 744.920 5.880 752.920 7.020 ;
  RECT 754.960 5.600 762.960 7.020 ;
  RECT 764.760 5.880 772.760 7.020 ;
  RECT 774.800 5.600 782.800 7.020 ;
  RECT 785.840 5.880 793.840 7.020 ;
  RECT 795.880 5.600 803.880 7.020 ;
  RECT 805.680 5.880 813.680 7.020 ;
  RECT 815.720 5.600 823.720 7.020 ;
  RECT 836.800 5.600 844.800 7.020 ;
  RECT 826.760 5.880 834.760 7.020 ;
  RECT 846.600 5.880 854.600 7.020 ;
  RECT 856.640 5.600 864.640 7.020 ;
  RECT 867.680 5.880 875.680 7.020 ;
  RECT 877.720 5.600 885.720 7.020 ;
  RECT 887.520 5.880 895.520 7.020 ;
  RECT 897.560 5.600 905.560 7.020 ;
  RECT 908.600 5.880 916.600 7.020 ;
  RECT 918.640 5.600 926.640 7.020 ;
  RECT 928.440 5.880 936.440 7.020 ;
  RECT 938.480 5.600 946.480 7.020 ;
  RECT 949.520 5.880 957.520 7.020 ;
  RECT 959.560 5.600 967.560 7.020 ;
  RECT 969.360 5.880 977.360 7.020 ;
  RECT 979.400 5.600 987.400 7.020 ;
  RECT 1000.480 5.600 1008.480 7.020 ;
  RECT 990.440 5.880 998.440 7.020 ;
  RECT 1010.280 5.880 1018.280 7.020 ;
  RECT 1020.320 5.600 1028.320 7.020 ;
  RECT 1031.360 5.880 1039.360 7.020 ;
  RECT 1041.400 5.600 1049.400 7.020 ;
  RECT 1051.200 5.880 1059.200 7.020 ;
  RECT 1061.240 5.600 1069.240 7.020 ;
  RECT 1072.280 5.880 1080.280 7.020 ;
  RECT 1082.320 5.600 1090.320 7.020 ;
  RECT 1092.120 5.880 1100.120 7.020 ;
  RECT 1102.160 5.600 1110.160 7.020 ;
  RECT 1113.200 5.880 1121.200 7.020 ;
  RECT 1123.240 5.600 1131.240 7.020 ;
  RECT 1133.040 5.880 1141.040 7.020 ;
  RECT 1143.080 5.600 1151.080 7.020 ;
  RECT 1164.160 5.600 1172.160 7.020 ;
  RECT 1154.120 5.880 1162.120 7.020 ;
  RECT 1173.960 5.880 1181.960 7.020 ;
  RECT 1184.000 5.600 1192.000 7.020 ;
  RECT 1195.040 5.880 1203.040 7.020 ;
  RECT 1205.080 5.600 1213.080 7.020 ;
  RECT 1214.880 5.880 1222.880 7.020 ;
  RECT 1224.920 5.600 1232.920 7.020 ;
  RECT 1235.960 5.880 1243.960 7.020 ;
  RECT 1246.000 5.600 1254.000 7.020 ;
  RECT 1255.800 5.880 1263.800 7.020 ;
  RECT 1265.840 5.600 1273.840 7.020 ;
  RECT 1276.880 5.880 1284.880 7.020 ;
  RECT 1286.920 5.600 1294.920 7.020 ;
  RECT 1296.720 5.880 1304.720 7.020 ;
  RECT 1306.760 5.600 1314.760 7.020 ;
  RECT 2687.800 559.940 2688.940 560.320 ;
  RECT 2687.800 552.020 2688.940 552.300 ;
  RECT 2687.800 548.340 2688.940 548.620 ;
  RECT 2687.800 544.660 2688.940 544.940 ;
  RECT 2687.800 540.980 2688.940 541.260 ;
  RECT 2687.800 537.300 2688.940 537.580 ;
  RECT 2687.800 533.620 2688.940 533.900 ;
  RECT 2687.800 529.940 2688.940 530.220 ;
  RECT 2687.800 526.260 2688.940 526.540 ;
  RECT 2687.800 522.580 2688.940 522.860 ;
  RECT 2687.800 518.900 2688.940 519.180 ;
  RECT 2687.800 515.220 2688.940 515.500 ;
  RECT 2687.800 511.540 2688.940 511.820 ;
  RECT 2687.800 507.860 2688.940 508.140 ;
  RECT 2687.800 504.180 2688.940 504.460 ;
  RECT 2687.800 500.500 2688.940 500.780 ;
  RECT 2687.800 496.820 2688.940 497.100 ;
  RECT 2687.800 493.140 2688.940 493.420 ;
  RECT 2687.800 489.460 2688.940 489.740 ;
  RECT 2687.800 485.780 2688.940 486.060 ;
  RECT 2687.800 482.100 2688.940 482.380 ;
  RECT 2687.800 478.420 2688.940 478.700 ;
  RECT 2687.800 474.740 2688.940 475.020 ;
  RECT 2687.800 471.060 2688.940 471.340 ;
  RECT 2687.800 467.380 2688.940 467.660 ;
  RECT 2687.800 463.700 2688.940 463.980 ;
  RECT 2687.800 460.020 2688.940 460.300 ;
  RECT 2687.800 456.340 2688.940 456.620 ;
  RECT 2687.800 452.660 2688.940 452.940 ;
  RECT 2687.800 448.980 2688.940 449.260 ;
  RECT 2687.800 445.300 2688.940 445.580 ;
  RECT 2687.800 441.620 2688.940 441.900 ;
  RECT 2687.800 437.940 2688.940 438.220 ;
  RECT 2687.800 434.260 2688.940 434.540 ;
  RECT 2687.800 430.580 2688.940 430.860 ;
  RECT 2687.800 426.900 2688.940 427.180 ;
  RECT 2687.800 423.220 2688.940 423.500 ;
  RECT 2687.800 419.540 2688.940 419.820 ;
  RECT 2687.800 415.860 2688.940 416.140 ;
  RECT 2687.800 412.180 2688.940 412.460 ;
  RECT 2687.800 408.500 2688.940 408.780 ;
  RECT 2687.800 404.820 2688.940 405.100 ;
  RECT 2687.800 401.140 2688.940 401.420 ;
  RECT 2687.800 397.460 2688.940 397.740 ;
  RECT 2687.800 393.780 2688.940 394.060 ;
  RECT 2687.800 390.100 2688.940 390.380 ;
  RECT 2687.800 386.420 2688.940 386.700 ;
  RECT 2687.800 382.740 2688.940 383.020 ;
  RECT 2687.800 379.060 2688.940 379.340 ;
  RECT 2687.800 375.380 2688.940 375.660 ;
  RECT 2687.800 371.700 2688.940 371.980 ;
  RECT 2687.800 368.020 2688.940 368.300 ;
  RECT 2687.800 364.340 2688.940 364.620 ;
  RECT 2687.800 360.660 2688.940 360.940 ;
  RECT 2687.800 356.980 2688.940 357.260 ;
  RECT 2687.800 353.300 2688.940 353.580 ;
  RECT 2687.800 349.620 2688.940 349.900 ;
  RECT 2687.800 345.940 2688.940 346.220 ;
  RECT 2687.800 342.260 2688.940 342.540 ;
  RECT 2687.800 338.580 2688.940 338.860 ;
  RECT 2687.800 334.900 2688.940 335.180 ;
  RECT 2687.800 331.220 2688.940 331.500 ;
  RECT 2687.800 327.540 2688.940 327.820 ;
  RECT 2687.800 323.860 2688.940 324.140 ;
  RECT 2687.800 320.180 2688.940 320.460 ;
  RECT 2687.800 316.500 2688.940 316.780 ;
  RECT 2687.800 312.820 2688.940 313.100 ;
  RECT 2687.800 309.140 2688.940 309.420 ;
  RECT 2687.800 305.460 2688.940 305.740 ;
  RECT 2687.800 301.780 2688.940 302.060 ;
  RECT 2687.800 298.100 2688.940 298.380 ;
  RECT 2687.800 294.420 2688.940 294.700 ;
  RECT 2687.800 290.740 2688.940 291.020 ;
  RECT 2687.800 287.060 2688.940 287.340 ;
  RECT 2687.800 283.380 2688.940 283.660 ;
  RECT 2687.800 279.700 2688.940 279.980 ;
  RECT 2687.800 276.020 2688.940 276.300 ;
  RECT 2687.800 272.340 2688.940 272.620 ;
  RECT 2687.800 268.660 2688.940 268.940 ;
  RECT 2687.800 264.980 2688.940 265.260 ;
  RECT 2687.800 261.300 2688.940 261.580 ;
  RECT 2687.800 257.620 2688.940 257.900 ;
  RECT 2687.800 253.940 2688.940 254.220 ;
  RECT 2687.800 250.260 2688.940 250.540 ;
  RECT 2687.800 246.580 2688.940 246.860 ;
  RECT 2687.800 242.900 2688.940 243.180 ;
  RECT 2687.800 239.220 2688.940 239.500 ;
  RECT 2687.800 235.540 2688.940 235.820 ;
  RECT 2687.800 231.860 2688.940 232.140 ;
  RECT 2687.800 228.180 2688.940 228.460 ;
  RECT 2687.800 224.500 2688.940 224.780 ;
  RECT 2687.800 220.820 2688.940 221.100 ;
  RECT 2687.800 217.140 2688.940 217.420 ;
  RECT 2687.800 213.460 2688.940 213.740 ;
  RECT 2687.800 209.780 2688.940 210.060 ;
  RECT 2687.800 206.100 2688.940 206.380 ;
  RECT 2687.800 202.420 2688.940 202.700 ;
  RECT 2687.800 198.740 2688.940 199.020 ;
  RECT 2687.800 195.060 2688.940 195.340 ;
  RECT 2687.800 191.380 2688.940 191.660 ;
  RECT 2687.800 187.700 2688.940 187.980 ;
  RECT 2687.800 184.020 2688.940 184.300 ;
  RECT 2687.800 180.340 2688.940 180.620 ;
  RECT 2687.800 176.660 2688.940 176.940 ;
  RECT 2687.800 172.980 2688.940 173.260 ;
  RECT 2687.800 169.300 2688.940 169.580 ;
  RECT 2687.800 165.620 2688.940 165.900 ;
  RECT 2687.800 161.940 2688.940 162.220 ;
  RECT 2687.800 158.260 2688.940 158.540 ;
  RECT 2687.800 154.580 2688.940 154.860 ;
  RECT 2687.800 150.900 2688.940 151.180 ;
  RECT 2687.800 147.220 2688.940 147.500 ;
  RECT 2687.800 143.540 2688.940 143.820 ;
  RECT 2687.800 139.860 2688.940 140.140 ;
  RECT 2687.800 136.180 2688.940 136.460 ;
  RECT 2687.800 132.500 2688.940 132.780 ;
  RECT 2687.800 128.820 2688.940 129.100 ;
  RECT 2687.800 125.140 2688.940 125.420 ;
  RECT 2687.800 121.460 2688.940 121.740 ;
  RECT 2687.800 117.780 2688.940 118.060 ;
  RECT 2687.800 114.100 2688.940 114.380 ;
  RECT 2687.800 110.420 2688.940 110.700 ;
  RECT 2687.800 106.740 2688.940 107.020 ;
  RECT 2687.800 103.060 2688.940 103.340 ;
  RECT 2687.800 99.380 2688.940 99.660 ;
  RECT 2687.800 95.700 2688.940 95.980 ;
  RECT 2687.800 92.020 2688.940 92.300 ;
  RECT 2687.800 88.340 2688.940 88.620 ;
  RECT 2687.800 84.660 2688.940 84.940 ;
  RECT 2687.800 80.980 2688.940 81.260 ;
  RECT 2687.800 77.300 2688.940 77.580 ;
  RECT 2687.800 73.620 2688.940 73.900 ;
  RECT 2687.800 69.940 2688.940 70.220 ;
  RECT 2687.800 65.600 2688.940 65.980 ;
  RECT 1376.820 560.790 1377.070 561.930 ;
  RECT 1417.740 560.790 1417.990 561.930 ;
  RECT 1458.660 560.790 1458.910 561.930 ;
  RECT 1499.580 560.790 1499.830 561.930 ;
  RECT 1540.500 560.790 1540.750 561.930 ;
  RECT 1581.420 560.790 1581.670 561.930 ;
  RECT 1622.340 560.790 1622.590 561.930 ;
  RECT 1663.260 560.790 1663.510 561.930 ;
  RECT 1704.180 560.790 1704.430 561.930 ;
  RECT 1745.100 560.790 1745.350 561.930 ;
  RECT 1786.020 560.790 1786.270 561.930 ;
  RECT 1826.940 560.790 1827.190 561.930 ;
  RECT 1867.860 560.790 1868.110 561.930 ;
  RECT 1908.780 560.790 1909.030 561.930 ;
  RECT 1949.700 560.790 1949.950 561.930 ;
  RECT 1990.620 560.790 1990.870 561.930 ;
  RECT 2031.540 560.790 2031.790 561.930 ;
  RECT 2072.460 560.790 2072.710 561.930 ;
  RECT 2113.380 560.790 2113.630 561.930 ;
  RECT 2154.300 560.790 2154.550 561.930 ;
  RECT 2195.220 560.790 2195.470 561.930 ;
  RECT 2236.140 560.790 2236.390 561.930 ;
  RECT 2277.060 560.790 2277.310 561.930 ;
  RECT 2317.980 560.790 2318.230 561.930 ;
  RECT 2358.900 560.790 2359.150 561.930 ;
  RECT 2399.820 560.790 2400.070 561.930 ;
  RECT 2440.740 560.790 2440.990 561.930 ;
  RECT 2481.660 560.790 2481.910 561.930 ;
  RECT 2522.580 560.790 2522.830 561.930 ;
  RECT 2563.500 560.790 2563.750 561.930 ;
  RECT 2604.420 560.790 2604.670 561.930 ;
  RECT 2645.340 560.790 2645.590 561.930 ;
  RECT 1359.810 560.790 1362.320 561.930 ;
  RECT 1347.390 560.790 1349.780 561.930 ;
  RECT 1339.880 560.790 1342.940 561.930 ;
  RECT 1364.060 560.790 1366.910 561.930 ;
  RECT 1368.360 560.790 1371.610 561.930 ;
  RECT 1337.160 560.790 1338.920 561.930 ;
  RECT 1319.820 560.790 1321.580 561.930 ;
  RECT 1323.820 560.790 1325.580 561.930 ;
  RECT 1327.820 560.790 1329.580 561.930 ;
  RECT 1331.820 560.790 1333.580 561.930 ;
  RECT 4.000 65.600 5.140 65.980 ;
  RECT 4.000 69.940 5.140 70.220 ;
  RECT 4.000 73.620 5.140 73.900 ;
  RECT 4.000 77.300 5.140 77.580 ;
  RECT 4.000 80.980 5.140 81.260 ;
  RECT 4.000 84.660 5.140 84.940 ;
  RECT 4.000 88.340 5.140 88.620 ;
  RECT 4.000 92.020 5.140 92.300 ;
  RECT 4.000 95.700 5.140 95.980 ;
  RECT 4.000 99.380 5.140 99.660 ;
  RECT 4.000 103.060 5.140 103.340 ;
  RECT 4.000 106.740 5.140 107.020 ;
  RECT 4.000 110.420 5.140 110.700 ;
  RECT 4.000 114.100 5.140 114.380 ;
  RECT 4.000 117.780 5.140 118.060 ;
  RECT 4.000 121.460 5.140 121.740 ;
  RECT 4.000 125.140 5.140 125.420 ;
  RECT 4.000 128.820 5.140 129.100 ;
  RECT 4.000 132.500 5.140 132.780 ;
  RECT 4.000 136.180 5.140 136.460 ;
  RECT 4.000 139.860 5.140 140.140 ;
  RECT 4.000 143.540 5.140 143.820 ;
  RECT 4.000 147.220 5.140 147.500 ;
  RECT 4.000 150.900 5.140 151.180 ;
  RECT 4.000 154.580 5.140 154.860 ;
  RECT 4.000 158.260 5.140 158.540 ;
  RECT 4.000 161.940 5.140 162.220 ;
  RECT 4.000 165.620 5.140 165.900 ;
  RECT 4.000 169.300 5.140 169.580 ;
  RECT 4.000 172.980 5.140 173.260 ;
  RECT 4.000 176.660 5.140 176.940 ;
  RECT 4.000 180.340 5.140 180.620 ;
  RECT 4.000 184.020 5.140 184.300 ;
  RECT 4.000 187.700 5.140 187.980 ;
  RECT 4.000 191.380 5.140 191.660 ;
  RECT 4.000 195.060 5.140 195.340 ;
  RECT 4.000 198.740 5.140 199.020 ;
  RECT 4.000 202.420 5.140 202.700 ;
  RECT 4.000 206.100 5.140 206.380 ;
  RECT 4.000 209.780 5.140 210.060 ;
  RECT 4.000 213.460 5.140 213.740 ;
  RECT 4.000 217.140 5.140 217.420 ;
  RECT 4.000 220.820 5.140 221.100 ;
  RECT 4.000 224.500 5.140 224.780 ;
  RECT 4.000 228.180 5.140 228.460 ;
  RECT 4.000 231.860 5.140 232.140 ;
  RECT 4.000 235.540 5.140 235.820 ;
  RECT 4.000 239.220 5.140 239.500 ;
  RECT 4.000 242.900 5.140 243.180 ;
  RECT 4.000 246.580 5.140 246.860 ;
  RECT 4.000 250.260 5.140 250.540 ;
  RECT 4.000 253.940 5.140 254.220 ;
  RECT 4.000 257.620 5.140 257.900 ;
  RECT 4.000 261.300 5.140 261.580 ;
  RECT 4.000 264.980 5.140 265.260 ;
  RECT 4.000 268.660 5.140 268.940 ;
  RECT 4.000 272.340 5.140 272.620 ;
  RECT 4.000 276.020 5.140 276.300 ;
  RECT 4.000 279.700 5.140 279.980 ;
  RECT 4.000 283.380 5.140 283.660 ;
  RECT 4.000 287.060 5.140 287.340 ;
  RECT 4.000 290.740 5.140 291.020 ;
  RECT 4.000 294.420 5.140 294.700 ;
  RECT 4.000 298.100 5.140 298.380 ;
  RECT 4.000 301.780 5.140 302.060 ;
  RECT 4.000 305.460 5.140 305.740 ;
  RECT 4.000 309.140 5.140 309.420 ;
  RECT 4.000 312.820 5.140 313.100 ;
  RECT 4.000 316.500 5.140 316.780 ;
  RECT 4.000 320.180 5.140 320.460 ;
  RECT 4.000 323.860 5.140 324.140 ;
  RECT 4.000 327.540 5.140 327.820 ;
  RECT 4.000 331.220 5.140 331.500 ;
  RECT 4.000 334.900 5.140 335.180 ;
  RECT 4.000 338.580 5.140 338.860 ;
  RECT 4.000 342.260 5.140 342.540 ;
  RECT 4.000 345.940 5.140 346.220 ;
  RECT 4.000 349.620 5.140 349.900 ;
  RECT 4.000 353.300 5.140 353.580 ;
  RECT 4.000 356.980 5.140 357.260 ;
  RECT 4.000 360.660 5.140 360.940 ;
  RECT 4.000 364.340 5.140 364.620 ;
  RECT 4.000 368.020 5.140 368.300 ;
  RECT 4.000 371.700 5.140 371.980 ;
  RECT 4.000 375.380 5.140 375.660 ;
  RECT 4.000 379.060 5.140 379.340 ;
  RECT 4.000 382.740 5.140 383.020 ;
  RECT 4.000 386.420 5.140 386.700 ;
  RECT 4.000 390.100 5.140 390.380 ;
  RECT 4.000 393.780 5.140 394.060 ;
  RECT 4.000 397.460 5.140 397.740 ;
  RECT 4.000 401.140 5.140 401.420 ;
  RECT 4.000 404.820 5.140 405.100 ;
  RECT 4.000 408.500 5.140 408.780 ;
  RECT 4.000 412.180 5.140 412.460 ;
  RECT 4.000 415.860 5.140 416.140 ;
  RECT 4.000 419.540 5.140 419.820 ;
  RECT 4.000 423.220 5.140 423.500 ;
  RECT 4.000 426.900 5.140 427.180 ;
  RECT 4.000 430.580 5.140 430.860 ;
  RECT 4.000 434.260 5.140 434.540 ;
  RECT 4.000 437.940 5.140 438.220 ;
  RECT 4.000 441.620 5.140 441.900 ;
  RECT 4.000 445.300 5.140 445.580 ;
  RECT 4.000 448.980 5.140 449.260 ;
  RECT 4.000 452.660 5.140 452.940 ;
  RECT 4.000 456.340 5.140 456.620 ;
  RECT 4.000 460.020 5.140 460.300 ;
  RECT 4.000 463.700 5.140 463.980 ;
  RECT 4.000 467.380 5.140 467.660 ;
  RECT 4.000 471.060 5.140 471.340 ;
  RECT 4.000 474.740 5.140 475.020 ;
  RECT 4.000 478.420 5.140 478.700 ;
  RECT 4.000 482.100 5.140 482.380 ;
  RECT 4.000 485.780 5.140 486.060 ;
  RECT 4.000 489.460 5.140 489.740 ;
  RECT 4.000 493.140 5.140 493.420 ;
  RECT 4.000 496.820 5.140 497.100 ;
  RECT 4.000 500.500 5.140 500.780 ;
  RECT 4.000 504.180 5.140 504.460 ;
  RECT 4.000 507.860 5.140 508.140 ;
  RECT 4.000 511.540 5.140 511.820 ;
  RECT 4.000 515.220 5.140 515.500 ;
  RECT 4.000 518.900 5.140 519.180 ;
  RECT 4.000 522.580 5.140 522.860 ;
  RECT 4.000 526.260 5.140 526.540 ;
  RECT 4.000 529.940 5.140 530.220 ;
  RECT 4.000 533.620 5.140 533.900 ;
  RECT 4.000 537.300 5.140 537.580 ;
  RECT 4.000 540.980 5.140 541.260 ;
  RECT 4.000 544.660 5.140 544.940 ;
  RECT 4.000 548.340 5.140 548.620 ;
  RECT 4.000 552.020 5.140 552.300 ;
  RECT 4.000 559.940 5.140 560.320 ;
  RECT 47.350 560.790 47.600 561.930 ;
  RECT 88.270 560.790 88.520 561.930 ;
  RECT 129.190 560.790 129.440 561.930 ;
  RECT 170.110 560.790 170.360 561.930 ;
  RECT 211.030 560.790 211.280 561.930 ;
  RECT 251.950 560.790 252.200 561.930 ;
  RECT 292.870 560.790 293.120 561.930 ;
  RECT 333.790 560.790 334.040 561.930 ;
  RECT 374.710 560.790 374.960 561.930 ;
  RECT 415.630 560.790 415.880 561.930 ;
  RECT 456.550 560.790 456.800 561.930 ;
  RECT 497.470 560.790 497.720 561.930 ;
  RECT 538.390 560.790 538.640 561.930 ;
  RECT 579.310 560.790 579.560 561.930 ;
  RECT 620.230 560.790 620.480 561.930 ;
  RECT 661.150 560.790 661.400 561.930 ;
  RECT 702.070 560.790 702.320 561.930 ;
  RECT 742.990 560.790 743.240 561.930 ;
  RECT 783.910 560.790 784.160 561.930 ;
  RECT 824.830 560.790 825.080 561.930 ;
  RECT 865.750 560.790 866.000 561.930 ;
  RECT 906.670 560.790 906.920 561.930 ;
  RECT 947.590 560.790 947.840 561.930 ;
  RECT 988.510 560.790 988.760 561.930 ;
  RECT 1029.430 560.790 1029.680 561.930 ;
  RECT 1070.350 560.790 1070.600 561.930 ;
  RECT 1111.270 560.790 1111.520 561.930 ;
  RECT 1152.190 560.790 1152.440 561.930 ;
  RECT 1193.110 560.790 1193.360 561.930 ;
  RECT 1234.030 560.790 1234.280 561.930 ;
  RECT 1274.950 560.790 1275.200 561.930 ;
  RECT 2.000 561.930 2690.940 563.930 ;
  RECT 2.000 3.600 2690.940 5.600 ;
  RECT 2688.940 3.600 2690.940 563.930 ;
  RECT 2.000 3.600 4.000 563.930 ;
  LAYER ME3 ;
  RECT 5.420 7.020 2687.520 560.510 ;
  RECT 2690.940 3.600 2692.940 563.930 ;
  RECT 0.000 3.600 2.000 563.930 ;
  RECT 2.000 563.930 2690.940 565.930 ;
  RECT 2.000 1.600 2690.940 3.600 ;
  RECT 2688.940 555.000 2690.660 561.930 ;
  RECT 2688.940 64.930 2690.660 67.240 ;
  RECT 2688.940 44.080 2690.660 61.260 ;
  RECT 2688.940 39.620 2690.660 41.480 ;
  RECT 2688.940 29.870 2690.660 33.520 ;
  RECT 2688.940 24.270 2690.660 26.870 ;
  RECT 2688.940 18.130 2690.660 21.270 ;
  RECT 2688.940 5.600 2690.660 11.230 ;
  RECT 2.280 555.000 4.000 561.930 ;
  RECT 2.280 64.930 4.000 67.240 ;
  RECT 2.280 44.080 4.000 61.260 ;
  RECT 2.280 39.620 4.000 41.480 ;
  RECT 2.280 29.870 4.000 33.520 ;
  RECT 2.280 24.270 4.000 26.870 ;
  RECT 2.280 18.130 4.000 21.270 ;
  RECT 2.280 5.600 4.000 11.230 ;
  RECT 2646.020 561.930 2688.940 563.650 ;
  RECT 2605.100 561.930 2643.770 563.650 ;
  RECT 2564.180 561.930 2602.850 563.650 ;
  RECT 2523.260 561.930 2561.930 563.650 ;
  RECT 2482.340 561.930 2521.010 563.650 ;
  RECT 2441.420 561.930 2480.090 563.650 ;
  RECT 2400.500 561.930 2439.170 563.650 ;
  RECT 2359.580 561.930 2398.250 563.650 ;
  RECT 2318.660 561.930 2357.330 563.650 ;
  RECT 2277.740 561.930 2316.410 563.650 ;
  RECT 2236.820 561.930 2275.490 563.650 ;
  RECT 2195.900 561.930 2234.570 563.650 ;
  RECT 2154.980 561.930 2193.650 563.650 ;
  RECT 2114.060 561.930 2152.730 563.650 ;
  RECT 2073.140 561.930 2111.810 563.650 ;
  RECT 2032.220 561.930 2070.890 563.650 ;
  RECT 1991.300 561.930 2029.970 563.650 ;
  RECT 1950.380 561.930 1989.050 563.650 ;
  RECT 1909.460 561.930 1948.130 563.650 ;
  RECT 1868.540 561.930 1907.210 563.650 ;
  RECT 1827.620 561.930 1866.290 563.650 ;
  RECT 1786.700 561.930 1825.370 563.650 ;
  RECT 1745.780 561.930 1784.450 563.650 ;
  RECT 1704.860 561.930 1743.530 563.650 ;
  RECT 1663.940 561.930 1702.610 563.650 ;
  RECT 1623.020 561.930 1661.690 563.650 ;
  RECT 1582.100 561.930 1620.770 563.650 ;
  RECT 1541.180 561.930 1579.850 563.650 ;
  RECT 1500.260 561.930 1538.930 563.650 ;
  RECT 1459.340 561.930 1498.010 563.650 ;
  RECT 1418.420 561.930 1457.090 563.650 ;
  RECT 1377.500 561.930 1416.170 563.650 ;
  RECT 1358.760 561.930 1371.760 563.650 ;
  RECT 1347.630 561.930 1352.440 563.650 ;
  RECT 1337.920 561.930 1342.440 563.650 ;
  RECT 1332.580 561.930 1334.160 563.650 ;
  RECT 1276.770 561.930 1315.800 563.650 ;
  RECT 1235.850 561.930 1274.520 563.650 ;
  RECT 1194.930 561.930 1233.600 563.650 ;
  RECT 1154.010 561.930 1192.680 563.650 ;
  RECT 1113.090 561.930 1151.760 563.650 ;
  RECT 1072.170 561.930 1110.840 563.650 ;
  RECT 1031.250 561.930 1069.920 563.650 ;
  RECT 990.330 561.930 1029.000 563.650 ;
  RECT 949.410 561.930 988.080 563.650 ;
  RECT 908.490 561.930 947.160 563.650 ;
  RECT 867.570 561.930 906.240 563.650 ;
  RECT 826.650 561.930 865.320 563.650 ;
  RECT 785.730 561.930 824.400 563.650 ;
  RECT 744.810 561.930 783.480 563.650 ;
  RECT 703.890 561.930 742.560 563.650 ;
  RECT 662.970 561.930 701.640 563.650 ;
  RECT 622.050 561.930 660.720 563.650 ;
  RECT 581.130 561.930 619.800 563.650 ;
  RECT 540.210 561.930 578.880 563.650 ;
  RECT 499.290 561.930 537.960 563.650 ;
  RECT 458.370 561.930 497.040 563.650 ;
  RECT 417.450 561.930 456.120 563.650 ;
  RECT 376.530 561.930 415.200 563.650 ;
  RECT 335.610 561.930 374.280 563.650 ;
  RECT 294.690 561.930 333.360 563.650 ;
  RECT 253.770 561.930 292.440 563.650 ;
  RECT 212.850 561.930 251.520 563.650 ;
  RECT 171.930 561.930 210.600 563.650 ;
  RECT 131.010 561.930 169.680 563.650 ;
  RECT 90.090 561.930 128.760 563.650 ;
  RECT 49.170 561.930 87.840 563.650 ;
  RECT 4.000 561.930 46.920 563.650 ;
  RECT 2675.540 3.880 2685.380 5.600 ;
  RECT 2655.700 3.880 2665.540 5.600 ;
  RECT 2634.620 3.880 2645.700 5.600 ;
  RECT 2614.780 3.880 2624.620 5.600 ;
  RECT 2593.700 3.880 2604.780 5.600 ;
  RECT 2573.860 3.880 2583.700 5.600 ;
  RECT 2552.780 3.880 2563.860 5.600 ;
  RECT 2532.940 3.880 2542.780 5.600 ;
  RECT 2511.860 3.880 2522.940 5.600 ;
  RECT 2492.020 3.880 2501.860 5.600 ;
  RECT 2470.940 3.880 2482.020 5.600 ;
  RECT 2451.100 3.880 2460.940 5.600 ;
  RECT 2430.020 3.880 2441.100 5.600 ;
  RECT 2410.180 3.880 2420.020 5.600 ;
  RECT 2389.100 3.880 2400.180 5.600 ;
  RECT 2369.260 3.880 2379.100 5.600 ;
  RECT 2348.180 3.880 2359.260 5.600 ;
  RECT 2328.340 3.880 2338.180 5.600 ;
  RECT 2307.260 3.880 2318.340 5.600 ;
  RECT 2287.420 3.880 2297.260 5.600 ;
  RECT 2266.340 3.880 2277.420 5.600 ;
  RECT 2246.500 3.880 2256.340 5.600 ;
  RECT 2225.420 3.880 2236.500 5.600 ;
  RECT 2205.580 3.880 2215.420 5.600 ;
  RECT 2184.500 3.880 2195.580 5.600 ;
  RECT 2164.660 3.880 2174.500 5.600 ;
  RECT 2143.580 3.880 2154.660 5.600 ;
  RECT 2123.740 3.880 2133.580 5.600 ;
  RECT 2102.660 3.880 2113.740 5.600 ;
  RECT 2082.820 3.880 2092.660 5.600 ;
  RECT 2061.740 3.880 2072.820 5.600 ;
  RECT 2041.900 3.880 2051.740 5.600 ;
  RECT 2020.820 3.880 2031.900 5.600 ;
  RECT 2000.980 3.880 2010.820 5.600 ;
  RECT 1979.900 3.880 1990.980 5.600 ;
  RECT 1960.060 3.880 1969.900 5.600 ;
  RECT 1938.980 3.880 1950.060 5.600 ;
  RECT 1919.140 3.880 1928.980 5.600 ;
  RECT 1898.060 3.880 1909.140 5.600 ;
  RECT 1878.220 3.880 1888.060 5.600 ;
  RECT 1857.140 3.880 1868.220 5.600 ;
  RECT 1837.300 3.880 1847.140 5.600 ;
  RECT 1816.220 3.880 1827.300 5.600 ;
  RECT 1796.380 3.880 1806.220 5.600 ;
  RECT 1775.300 3.880 1786.380 5.600 ;
  RECT 1755.460 3.880 1765.300 5.600 ;
  RECT 1734.380 3.880 1745.460 5.600 ;
  RECT 1714.540 3.880 1724.380 5.600 ;
  RECT 1693.460 3.880 1704.540 5.600 ;
  RECT 1673.620 3.880 1683.460 5.600 ;
  RECT 1652.540 3.880 1663.620 5.600 ;
  RECT 1632.700 3.880 1642.540 5.600 ;
  RECT 1611.620 3.880 1622.700 5.600 ;
  RECT 1591.780 3.880 1601.620 5.600 ;
  RECT 1570.700 3.880 1581.780 5.600 ;
  RECT 1550.860 3.880 1560.700 5.600 ;
  RECT 1529.780 3.880 1540.860 5.600 ;
  RECT 1509.940 3.880 1519.780 5.600 ;
  RECT 1488.860 3.880 1499.940 5.600 ;
  RECT 1469.020 3.880 1478.860 5.600 ;
  RECT 1447.940 3.880 1459.020 5.600 ;
  RECT 1428.100 3.880 1437.940 5.600 ;
  RECT 1407.020 3.880 1418.100 5.600 ;
  RECT 1387.180 3.880 1397.020 5.600 ;
  RECT 1359.210 3.880 1377.180 5.600 ;
  RECT 1347.890 3.880 1351.290 5.600 ;
  RECT 1337.920 3.880 1342.440 5.600 ;
  RECT 1332.580 3.880 1334.160 5.600 ;
  RECT 1305.720 3.880 1316.820 5.600 ;
  RECT 1285.880 3.880 1295.720 5.600 ;
  RECT 1264.800 3.880 1275.880 5.600 ;
  RECT 1244.960 3.880 1254.800 5.600 ;
  RECT 1223.880 3.880 1234.960 5.600 ;
  RECT 1204.040 3.880 1213.880 5.600 ;
  RECT 1182.960 3.880 1194.040 5.600 ;
  RECT 1163.120 3.880 1172.960 5.600 ;
  RECT 1142.040 3.880 1153.120 5.600 ;
  RECT 1122.200 3.880 1132.040 5.600 ;
  RECT 1101.120 3.880 1112.200 5.600 ;
  RECT 1081.280 3.880 1091.120 5.600 ;
  RECT 1060.200 3.880 1071.280 5.600 ;
  RECT 1040.360 3.880 1050.200 5.600 ;
  RECT 1019.280 3.880 1030.360 5.600 ;
  RECT 999.440 3.880 1009.280 5.600 ;
  RECT 978.360 3.880 989.440 5.600 ;
  RECT 958.520 3.880 968.360 5.600 ;
  RECT 937.440 3.880 948.520 5.600 ;
  RECT 917.600 3.880 927.440 5.600 ;
  RECT 896.520 3.880 907.600 5.600 ;
  RECT 876.680 3.880 886.520 5.600 ;
  RECT 855.600 3.880 866.680 5.600 ;
  RECT 835.760 3.880 845.600 5.600 ;
  RECT 814.680 3.880 825.760 5.600 ;
  RECT 794.840 3.880 804.680 5.600 ;
  RECT 773.760 3.880 784.840 5.600 ;
  RECT 753.920 3.880 763.760 5.600 ;
  RECT 732.840 3.880 743.920 5.600 ;
  RECT 713.000 3.880 722.840 5.600 ;
  RECT 691.920 3.880 703.000 5.600 ;
  RECT 672.080 3.880 681.920 5.600 ;
  RECT 651.000 3.880 662.080 5.600 ;
  RECT 631.160 3.880 641.000 5.600 ;
  RECT 610.080 3.880 621.160 5.600 ;
  RECT 590.240 3.880 600.080 5.600 ;
  RECT 569.160 3.880 580.240 5.600 ;
  RECT 549.320 3.880 559.160 5.600 ;
  RECT 528.240 3.880 539.320 5.600 ;
  RECT 508.400 3.880 518.240 5.600 ;
  RECT 487.320 3.880 498.400 5.600 ;
  RECT 467.480 3.880 477.320 5.600 ;
  RECT 446.400 3.880 457.480 5.600 ;
  RECT 426.560 3.880 436.400 5.600 ;
  RECT 405.480 3.880 416.560 5.600 ;
  RECT 385.640 3.880 395.480 5.600 ;
  RECT 364.560 3.880 375.640 5.600 ;
  RECT 344.720 3.880 354.560 5.600 ;
  RECT 323.640 3.880 334.720 5.600 ;
  RECT 303.800 3.880 313.640 5.600 ;
  RECT 282.720 3.880 293.800 5.600 ;
  RECT 262.880 3.880 272.720 5.600 ;
  RECT 241.800 3.880 252.880 5.600 ;
  RECT 221.960 3.880 231.800 5.600 ;
  RECT 200.880 3.880 211.960 5.600 ;
  RECT 181.040 3.880 190.880 5.600 ;
  RECT 159.960 3.880 171.040 5.600 ;
  RECT 140.120 3.880 149.960 5.600 ;
  RECT 119.040 3.880 130.120 5.600 ;
  RECT 99.200 3.880 109.040 5.600 ;
  RECT 78.120 3.880 89.200 5.600 ;
  RECT 58.280 3.880 68.120 5.600 ;
  RECT 37.200 3.880 48.280 5.600 ;
  RECT 17.360 3.880 27.200 5.600 ;
  RECT 2.280 561.930 4.000 563.650 ;
  RECT 0.000 563.930 2.000 565.930 ;
  RECT 2688.940 3.880 2690.660 5.600 ;
  RECT 2690.940 1.600 2692.940 3.600 ;
  RECT 2688.940 561.930 2690.660 563.650 ;
  RECT 2690.940 563.930 2692.940 565.930 ;
  RECT 2.280 3.880 4.000 5.600 ;
  RECT 0.000 1.600 2.000 3.600 ;
  RECT 2680.800 0.000 2681.600 1.000 ;
  RECT 2666.400 0.000 2667.200 1.000 ;
  RECT 2661.200 0.000 2662.000 1.000 ;
  RECT 2646.400 0.000 2647.200 1.000 ;
  RECT 2640.000 0.000 2640.800 1.000 ;
  RECT 2625.600 0.000 2626.400 1.000 ;
  RECT 2620.400 0.000 2621.200 1.000 ;
  RECT 2605.600 0.000 2606.400 1.000 ;
  RECT 2599.200 0.000 2600.000 1.000 ;
  RECT 2584.400 0.000 2585.200 1.000 ;
  RECT 2579.200 0.000 2580.000 1.000 ;
  RECT 2564.800 0.000 2565.600 1.000 ;
  RECT 2558.400 0.000 2559.200 1.000 ;
  RECT 2543.600 0.000 2544.400 1.000 ;
  RECT 2538.400 0.000 2539.200 1.000 ;
  RECT 2525.600 0.000 2526.400 1.000 ;
  RECT 2523.600 0.000 2524.400 1.000 ;
  RECT 2517.200 0.000 2518.000 1.000 ;
  RECT 2502.800 0.000 2503.600 1.000 ;
  RECT 2497.600 0.000 2498.400 1.000 ;
  RECT 2482.800 0.000 2483.600 1.000 ;
  RECT 2476.400 0.000 2477.200 1.000 ;
  RECT 2461.600 0.000 2462.400 1.000 ;
  RECT 2456.400 0.000 2457.200 1.000 ;
  RECT 2442.000 0.000 2442.800 1.000 ;
  RECT 2435.600 0.000 2436.400 1.000 ;
  RECT 2420.800 0.000 2421.600 1.000 ;
  RECT 2415.600 0.000 2416.400 1.000 ;
  RECT 2400.800 0.000 2401.600 1.000 ;
  RECT 2394.400 0.000 2395.200 1.000 ;
  RECT 2380.000 0.000 2380.800 1.000 ;
  RECT 2374.800 0.000 2375.600 1.000 ;
  RECT 2361.600 0.000 2362.400 1.000 ;
  RECT 2360.000 0.000 2360.800 1.000 ;
  RECT 2353.600 0.000 2354.400 1.000 ;
  RECT 2338.800 0.000 2339.600 1.000 ;
  RECT 2333.600 0.000 2334.400 1.000 ;
  RECT 2319.200 0.000 2320.000 1.000 ;
  RECT 2312.800 0.000 2313.600 1.000 ;
  RECT 2298.000 0.000 2298.800 1.000 ;
  RECT 2292.800 0.000 2293.600 1.000 ;
  RECT 2278.400 0.000 2279.200 1.000 ;
  RECT 2271.600 0.000 2272.400 1.000 ;
  RECT 2257.200 0.000 2258.000 1.000 ;
  RECT 2252.000 0.000 2252.800 1.000 ;
  RECT 2237.200 0.000 2238.000 1.000 ;
  RECT 2230.800 0.000 2231.600 1.000 ;
  RECT 2216.400 0.000 2217.200 1.000 ;
  RECT 2211.200 0.000 2212.000 1.000 ;
  RECT 2198.000 0.000 2198.800 1.000 ;
  RECT 2196.400 0.000 2197.200 1.000 ;
  RECT 2190.000 0.000 2190.800 1.000 ;
  RECT 2175.200 0.000 2176.000 1.000 ;
  RECT 2170.000 0.000 2170.800 1.000 ;
  RECT 2155.600 0.000 2156.400 1.000 ;
  RECT 2149.200 0.000 2150.000 1.000 ;
  RECT 2134.400 0.000 2135.200 1.000 ;
  RECT 2129.200 0.000 2130.000 1.000 ;
  RECT 2114.400 0.000 2115.200 1.000 ;
  RECT 2108.000 0.000 2108.800 1.000 ;
  RECT 2093.600 0.000 2094.400 1.000 ;
  RECT 2088.400 0.000 2089.200 1.000 ;
  RECT 2073.600 0.000 2074.400 1.000 ;
  RECT 2067.200 0.000 2068.000 1.000 ;
  RECT 2052.400 0.000 2053.200 1.000 ;
  RECT 2047.200 0.000 2048.000 1.000 ;
  RECT 2034.400 0.000 2035.200 1.000 ;
  RECT 2032.800 0.000 2033.600 1.000 ;
  RECT 2026.400 0.000 2027.200 1.000 ;
  RECT 2011.600 0.000 2012.400 1.000 ;
  RECT 2006.400 0.000 2007.200 1.000 ;
  RECT 1991.600 0.000 1992.400 1.000 ;
  RECT 1985.200 0.000 1986.000 1.000 ;
  RECT 1970.800 0.000 1971.600 1.000 ;
  RECT 1965.600 0.000 1966.400 1.000 ;
  RECT 1950.800 0.000 1951.600 1.000 ;
  RECT 1944.400 0.000 1945.200 1.000 ;
  RECT 1929.600 0.000 1930.400 1.000 ;
  RECT 1924.400 0.000 1925.200 1.000 ;
  RECT 1910.000 0.000 1910.800 1.000 ;
  RECT 1903.600 0.000 1904.400 1.000 ;
  RECT 1888.800 0.000 1889.600 1.000 ;
  RECT 1883.600 0.000 1884.400 1.000 ;
  RECT 1870.800 0.000 1871.600 1.000 ;
  RECT 1869.200 0.000 1870.000 1.000 ;
  RECT 1862.400 0.000 1863.200 1.000 ;
  RECT 1848.000 0.000 1848.800 1.000 ;
  RECT 1842.800 0.000 1843.600 1.000 ;
  RECT 1828.000 0.000 1828.800 1.000 ;
  RECT 1821.600 0.000 1822.400 1.000 ;
  RECT 1807.200 0.000 1808.000 1.000 ;
  RECT 1802.000 0.000 1802.800 1.000 ;
  RECT 1787.200 0.000 1788.000 1.000 ;
  RECT 1780.800 0.000 1781.600 1.000 ;
  RECT 1766.000 0.000 1766.800 1.000 ;
  RECT 1760.800 0.000 1761.600 1.000 ;
  RECT 1746.400 0.000 1747.200 1.000 ;
  RECT 1740.000 0.000 1740.800 1.000 ;
  RECT 1725.200 0.000 1726.000 1.000 ;
  RECT 1720.000 0.000 1720.800 1.000 ;
  RECT 1707.200 0.000 1708.000 1.000 ;
  RECT 1705.200 0.000 1706.000 1.000 ;
  RECT 1698.800 0.000 1699.600 1.000 ;
  RECT 1684.400 0.000 1685.200 1.000 ;
  RECT 1679.200 0.000 1680.000 1.000 ;
  RECT 1664.400 0.000 1665.200 1.000 ;
  RECT 1658.000 0.000 1658.800 1.000 ;
  RECT 1643.200 0.000 1644.000 1.000 ;
  RECT 1638.000 0.000 1638.800 1.000 ;
  RECT 1623.600 0.000 1624.400 1.000 ;
  RECT 1617.200 0.000 1618.000 1.000 ;
  RECT 1602.400 0.000 1603.200 1.000 ;
  RECT 1597.200 0.000 1598.000 1.000 ;
  RECT 1582.400 0.000 1583.200 1.000 ;
  RECT 1576.000 0.000 1576.800 1.000 ;
  RECT 1561.600 0.000 1562.400 1.000 ;
  RECT 1556.400 0.000 1557.200 1.000 ;
  RECT 1543.200 0.000 1544.000 1.000 ;
  RECT 1541.600 0.000 1542.400 1.000 ;
  RECT 1535.200 0.000 1536.000 1.000 ;
  RECT 1520.400 0.000 1521.200 1.000 ;
  RECT 1515.200 0.000 1516.000 1.000 ;
  RECT 1500.800 0.000 1501.600 1.000 ;
  RECT 1494.400 0.000 1495.200 1.000 ;
  RECT 1479.600 0.000 1480.400 1.000 ;
  RECT 1474.400 0.000 1475.200 1.000 ;
  RECT 1460.000 0.000 1460.800 1.000 ;
  RECT 1453.200 0.000 1454.000 1.000 ;
  RECT 1438.800 0.000 1439.600 1.000 ;
  RECT 1433.600 0.000 1434.400 1.000 ;
  RECT 1418.800 0.000 1419.600 1.000 ;
  RECT 1412.400 0.000 1413.200 1.000 ;
  RECT 1398.000 0.000 1398.800 1.000 ;
  RECT 1392.800 0.000 1393.600 1.000 ;
  RECT 1379.600 0.000 1380.400 1.000 ;
  RECT 1378.000 0.000 1378.800 1.000 ;
  RECT 1357.200 0.000 1358.000 1.000 ;
  RECT 1356.000 0.000 1356.800 1.000 ;
  RECT 1354.800 0.000 1355.600 1.000 ;
  RECT 1353.600 0.000 1354.400 1.000 ;
  RECT 1352.400 0.000 1353.200 1.000 ;
  RECT 1351.200 0.000 1352.000 1.000 ;
  RECT 1345.200 0.000 1346.000 1.000 ;
  RECT 1338.000 0.000 1338.800 1.000 ;
  RECT 1335.200 0.000 1336.000 1.000 ;
  RECT 1332.400 0.000 1333.200 1.000 ;
  RECT 1330.000 0.000 1330.800 1.000 ;
  RECT 1328.400 0.000 1329.200 1.000 ;
  RECT 1326.000 0.000 1326.800 1.000 ;
  RECT 1324.400 0.000 1325.200 1.000 ;
  RECT 1322.000 0.000 1322.800 1.000 ;
  RECT 1320.400 0.000 1321.200 1.000 ;
  RECT 1311.200 0.000 1312.000 1.000 ;
  RECT 1296.400 0.000 1297.200 1.000 ;
  RECT 1291.200 0.000 1292.000 1.000 ;
  RECT 1276.800 0.000 1277.600 1.000 ;
  RECT 1270.400 0.000 1271.200 1.000 ;
  RECT 1255.600 0.000 1256.400 1.000 ;
  RECT 1250.400 0.000 1251.200 1.000 ;
  RECT 1235.600 0.000 1236.400 1.000 ;
  RECT 1229.200 0.000 1230.000 1.000 ;
  RECT 1214.800 0.000 1215.600 1.000 ;
  RECT 1209.600 0.000 1210.400 1.000 ;
  RECT 1194.800 0.000 1195.600 1.000 ;
  RECT 1188.400 0.000 1189.200 1.000 ;
  RECT 1173.600 0.000 1174.400 1.000 ;
  RECT 1168.400 0.000 1169.200 1.000 ;
  RECT 1155.600 0.000 1156.400 1.000 ;
  RECT 1154.000 0.000 1154.800 1.000 ;
  RECT 1147.600 0.000 1148.400 1.000 ;
  RECT 1132.800 0.000 1133.600 1.000 ;
  RECT 1127.600 0.000 1128.400 1.000 ;
  RECT 1113.200 0.000 1114.000 1.000 ;
  RECT 1106.400 0.000 1107.200 1.000 ;
  RECT 1092.000 0.000 1092.800 1.000 ;
  RECT 1086.800 0.000 1087.600 1.000 ;
  RECT 1072.000 0.000 1072.800 1.000 ;
  RECT 1065.600 0.000 1066.400 1.000 ;
  RECT 1051.200 0.000 1052.000 1.000 ;
  RECT 1045.600 0.000 1046.400 1.000 ;
  RECT 1031.200 0.000 1032.000 1.000 ;
  RECT 1024.800 0.000 1025.600 1.000 ;
  RECT 1010.000 0.000 1010.800 1.000 ;
  RECT 1004.800 0.000 1005.600 1.000 ;
  RECT 992.000 0.000 992.800 1.000 ;
  RECT 990.400 0.000 991.200 1.000 ;
  RECT 983.600 0.000 984.400 1.000 ;
  RECT 969.200 0.000 970.000 1.000 ;
  RECT 964.000 0.000 964.800 1.000 ;
  RECT 949.200 0.000 950.000 1.000 ;
  RECT 942.800 0.000 943.600 1.000 ;
  RECT 928.400 0.000 929.200 1.000 ;
  RECT 923.200 0.000 924.000 1.000 ;
  RECT 908.400 0.000 909.200 1.000 ;
  RECT 902.000 0.000 902.800 1.000 ;
  RECT 887.200 0.000 888.000 1.000 ;
  RECT 882.000 0.000 882.800 1.000 ;
  RECT 867.600 0.000 868.400 1.000 ;
  RECT 861.200 0.000 862.000 1.000 ;
  RECT 846.400 0.000 847.200 1.000 ;
  RECT 841.200 0.000 842.000 1.000 ;
  RECT 828.400 0.000 829.200 1.000 ;
  RECT 826.400 0.000 827.200 1.000 ;
  RECT 820.000 0.000 820.800 1.000 ;
  RECT 805.600 0.000 806.400 1.000 ;
  RECT 800.400 0.000 801.200 1.000 ;
  RECT 785.600 0.000 786.400 1.000 ;
  RECT 779.200 0.000 780.000 1.000 ;
  RECT 764.400 0.000 765.200 1.000 ;
  RECT 759.200 0.000 760.000 1.000 ;
  RECT 744.800 0.000 745.600 1.000 ;
  RECT 738.400 0.000 739.200 1.000 ;
  RECT 723.600 0.000 724.400 1.000 ;
  RECT 718.400 0.000 719.200 1.000 ;
  RECT 704.000 0.000 704.800 1.000 ;
  RECT 697.200 0.000 698.000 1.000 ;
  RECT 682.800 0.000 683.600 1.000 ;
  RECT 677.600 0.000 678.400 1.000 ;
  RECT 664.800 0.000 665.600 1.000 ;
  RECT 662.800 0.000 663.600 1.000 ;
  RECT 656.400 0.000 657.200 1.000 ;
  RECT 642.000 0.000 642.800 1.000 ;
  RECT 636.400 0.000 637.200 1.000 ;
  RECT 622.000 0.000 622.800 1.000 ;
  RECT 615.600 0.000 616.400 1.000 ;
  RECT 600.800 0.000 601.600 1.000 ;
  RECT 595.600 0.000 596.400 1.000 ;
  RECT 581.200 0.000 582.000 1.000 ;
  RECT 574.400 0.000 575.200 1.000 ;
  RECT 560.000 0.000 560.800 1.000 ;
  RECT 554.800 0.000 555.600 1.000 ;
  RECT 540.000 0.000 540.800 1.000 ;
  RECT 533.600 0.000 534.400 1.000 ;
  RECT 519.200 0.000 520.000 1.000 ;
  RECT 514.000 0.000 514.800 1.000 ;
  RECT 500.800 0.000 501.600 1.000 ;
  RECT 499.200 0.000 500.000 1.000 ;
  RECT 492.800 0.000 493.600 1.000 ;
  RECT 478.000 0.000 478.800 1.000 ;
  RECT 472.800 0.000 473.600 1.000 ;
  RECT 458.400 0.000 459.200 1.000 ;
  RECT 452.000 0.000 452.800 1.000 ;
  RECT 437.200 0.000 438.000 1.000 ;
  RECT 432.000 0.000 432.800 1.000 ;
  RECT 417.200 0.000 418.000 1.000 ;
  RECT 410.800 0.000 411.600 1.000 ;
  RECT 396.400 0.000 397.200 1.000 ;
  RECT 391.200 0.000 392.000 1.000 ;
  RECT 376.400 0.000 377.200 1.000 ;
  RECT 370.000 0.000 370.800 1.000 ;
  RECT 355.200 0.000 356.000 1.000 ;
  RECT 350.000 0.000 350.800 1.000 ;
  RECT 337.200 0.000 338.000 1.000 ;
  RECT 335.600 0.000 336.400 1.000 ;
  RECT 329.200 0.000 330.000 1.000 ;
  RECT 314.400 0.000 315.200 1.000 ;
  RECT 309.200 0.000 310.000 1.000 ;
  RECT 294.800 0.000 295.600 1.000 ;
  RECT 288.000 0.000 288.800 1.000 ;
  RECT 273.600 0.000 274.400 1.000 ;
  RECT 268.400 0.000 269.200 1.000 ;
  RECT 253.600 0.000 254.400 1.000 ;
  RECT 247.200 0.000 248.000 1.000 ;
  RECT 232.800 0.000 233.600 1.000 ;
  RECT 227.200 0.000 228.000 1.000 ;
  RECT 212.800 0.000 213.600 1.000 ;
  RECT 206.400 0.000 207.200 1.000 ;
  RECT 191.600 0.000 192.400 1.000 ;
  RECT 186.400 0.000 187.200 1.000 ;
  RECT 173.600 0.000 174.400 1.000 ;
  RECT 172.000 0.000 172.800 1.000 ;
  RECT 165.200 0.000 166.000 1.000 ;
  RECT 150.800 0.000 151.600 1.000 ;
  RECT 145.600 0.000 146.400 1.000 ;
  RECT 130.800 0.000 131.600 1.000 ;
  RECT 124.400 0.000 125.200 1.000 ;
  RECT 110.000 0.000 110.800 1.000 ;
  RECT 104.800 0.000 105.600 1.000 ;
  RECT 90.000 0.000 90.800 1.000 ;
  RECT 83.600 0.000 84.400 1.000 ;
  RECT 68.800 0.000 69.600 1.000 ;
  RECT 63.600 0.000 64.400 1.000 ;
  RECT 49.200 0.000 50.000 1.000 ;
  RECT 42.800 0.000 43.600 1.000 ;
  RECT 28.000 0.000 28.800 1.000 ;
  RECT 22.800 0.000 23.600 1.000 ;
  RECT 10.000 0.000 10.800 1.000 ;
  RECT 8.000 0.000 8.800 1.000 ;
  RECT 2687.520 62.260 2690.940 63.930 ;
  RECT 2687.520 22.270 2690.940 23.270 ;
  RECT 2687.520 16.130 2690.940 17.130 ;
  RECT 2687.520 12.230 2690.940 13.230 ;
  RECT 2687.520 27.870 2690.940 28.870 ;
  RECT 2687.520 42.480 2690.940 43.080 ;
  RECT 2687.520 37.620 2690.940 38.620 ;
  RECT 2687.520 34.520 2690.940 36.020 ;
  RECT 2687.800 9.570 2688.660 11.170 ;
  RECT 2687.800 14.200 2688.660 15.200 ;
  RECT 2687.800 18.730 2688.660 19.730 ;
  RECT 2687.800 21.230 2688.660 22.070 ;
  RECT 2687.800 24.170 2688.660 25.170 ;
  RECT 2687.800 36.320 2688.660 37.320 ;
  RECT 2687.800 39.480 2688.660 40.080 ;
  RECT 2687.800 45.560 2688.660 46.160 ;
  RECT 2687.800 57.100 2688.660 61.420 ;
  RECT 2686.380 3.600 2687.520 6.740 ;
  RECT 1378.180 3.600 1386.180 6.740 ;
  RECT 1398.020 3.600 1406.020 6.740 ;
  RECT 1419.100 3.600 1427.100 6.740 ;
  RECT 1438.940 3.600 1446.940 6.740 ;
  RECT 1460.020 3.600 1468.020 6.740 ;
  RECT 1479.860 3.600 1487.860 6.740 ;
  RECT 1500.940 3.600 1508.940 6.740 ;
  RECT 1520.780 3.600 1528.780 6.740 ;
  RECT 1541.860 3.600 1549.860 6.740 ;
  RECT 1561.700 3.600 1569.700 6.740 ;
  RECT 1582.780 3.600 1590.780 6.740 ;
  RECT 1602.620 3.600 1610.620 6.740 ;
  RECT 1623.700 3.600 1631.700 6.740 ;
  RECT 1643.540 3.600 1651.540 6.740 ;
  RECT 1664.620 3.600 1672.620 6.740 ;
  RECT 1684.460 3.600 1692.460 6.740 ;
  RECT 1705.540 3.600 1713.540 6.740 ;
  RECT 1725.380 3.600 1733.380 6.740 ;
  RECT 1746.460 3.600 1754.460 6.740 ;
  RECT 1766.300 3.600 1774.300 6.740 ;
  RECT 1787.380 3.600 1795.380 6.740 ;
  RECT 1807.220 3.600 1815.220 6.740 ;
  RECT 1828.300 3.600 1836.300 6.740 ;
  RECT 1848.140 3.600 1856.140 6.740 ;
  RECT 1869.220 3.600 1877.220 6.740 ;
  RECT 1889.060 3.600 1897.060 6.740 ;
  RECT 1910.140 3.600 1918.140 6.740 ;
  RECT 1929.980 3.600 1937.980 6.740 ;
  RECT 1951.060 3.600 1959.060 6.740 ;
  RECT 1970.900 3.600 1978.900 6.740 ;
  RECT 1991.980 3.600 1999.980 6.740 ;
  RECT 2011.820 3.600 2019.820 6.740 ;
  RECT 2032.900 3.600 2040.900 6.740 ;
  RECT 2052.740 3.600 2060.740 6.740 ;
  RECT 2073.820 3.600 2081.820 6.740 ;
  RECT 2093.660 3.600 2101.660 6.740 ;
  RECT 2114.740 3.600 2122.740 6.740 ;
  RECT 2134.580 3.600 2142.580 6.740 ;
  RECT 2155.660 3.600 2163.660 6.740 ;
  RECT 2175.500 3.600 2183.500 6.740 ;
  RECT 2196.580 3.600 2204.580 6.740 ;
  RECT 2216.420 3.600 2224.420 6.740 ;
  RECT 2237.500 3.600 2245.500 6.740 ;
  RECT 2257.340 3.600 2265.340 6.740 ;
  RECT 2278.420 3.600 2286.420 6.740 ;
  RECT 2298.260 3.600 2306.260 6.740 ;
  RECT 2319.340 3.600 2327.340 6.740 ;
  RECT 2339.180 3.600 2347.180 6.740 ;
  RECT 2360.260 3.600 2368.260 6.740 ;
  RECT 2380.100 3.600 2388.100 6.740 ;
  RECT 2401.180 3.600 2409.180 6.740 ;
  RECT 2421.020 3.600 2429.020 6.740 ;
  RECT 2442.100 3.600 2450.100 6.740 ;
  RECT 2461.940 3.600 2469.940 6.740 ;
  RECT 2483.020 3.600 2491.020 6.740 ;
  RECT 2502.860 3.600 2510.860 6.740 ;
  RECT 2523.940 3.600 2531.940 6.740 ;
  RECT 2543.780 3.600 2551.780 6.740 ;
  RECT 2564.860 3.600 2572.860 6.740 ;
  RECT 2584.700 3.600 2592.700 6.740 ;
  RECT 2605.780 3.600 2613.780 6.740 ;
  RECT 2625.620 3.600 2633.620 6.740 ;
  RECT 2646.700 3.600 2654.700 6.740 ;
  RECT 2666.540 3.600 2674.540 6.740 ;
  RECT 1343.440 3.600 1346.890 6.740 ;
  RECT 1352.290 3.600 1358.210 6.740 ;
  RECT 1335.160 3.600 1336.920 6.740 ;
  RECT 1329.820 3.600 1331.580 6.740 ;
  RECT 1325.820 3.600 1327.580 6.740 ;
  RECT 1321.820 3.600 1323.580 6.740 ;
  RECT 1317.820 3.600 1319.580 6.740 ;
  RECT 4.280 57.100 5.140 61.420 ;
  RECT 4.280 45.560 5.140 46.160 ;
  RECT 4.280 39.480 5.140 40.080 ;
  RECT 4.280 36.320 5.140 37.320 ;
  RECT 4.280 24.170 5.140 25.170 ;
  RECT 4.280 21.230 5.140 22.070 ;
  RECT 4.280 18.730 5.140 19.730 ;
  RECT 4.280 14.200 5.140 15.200 ;
  RECT 4.280 9.570 5.140 11.170 ;
  RECT 2.000 34.520 5.420 36.020 ;
  RECT 2.000 37.620 5.420 38.620 ;
  RECT 2.000 42.480 5.420 43.080 ;
  RECT 2.000 27.870 5.420 28.870 ;
  RECT 2.000 12.230 5.420 13.230 ;
  RECT 2.000 16.130 5.420 17.130 ;
  RECT 2.000 22.270 5.420 23.270 ;
  RECT 2.000 62.260 5.420 63.930 ;
  RECT 5.420 3.600 6.560 6.740 ;
  RECT 8.360 3.600 16.360 6.740 ;
  RECT 28.200 3.600 36.200 6.740 ;
  RECT 49.280 3.600 57.280 6.740 ;
  RECT 69.120 3.600 77.120 6.740 ;
  RECT 90.200 3.600 98.200 6.740 ;
  RECT 110.040 3.600 118.040 6.740 ;
  RECT 131.120 3.600 139.120 6.740 ;
  RECT 150.960 3.600 158.960 6.740 ;
  RECT 172.040 3.600 180.040 6.740 ;
  RECT 191.880 3.600 199.880 6.740 ;
  RECT 212.960 3.600 220.960 6.740 ;
  RECT 232.800 3.600 240.800 6.740 ;
  RECT 253.880 3.600 261.880 6.740 ;
  RECT 273.720 3.600 281.720 6.740 ;
  RECT 294.800 3.600 302.800 6.740 ;
  RECT 314.640 3.600 322.640 6.740 ;
  RECT 335.720 3.600 343.720 6.740 ;
  RECT 355.560 3.600 363.560 6.740 ;
  RECT 376.640 3.600 384.640 6.740 ;
  RECT 396.480 3.600 404.480 6.740 ;
  RECT 417.560 3.600 425.560 6.740 ;
  RECT 437.400 3.600 445.400 6.740 ;
  RECT 458.480 3.600 466.480 6.740 ;
  RECT 478.320 3.600 486.320 6.740 ;
  RECT 499.400 3.600 507.400 6.740 ;
  RECT 519.240 3.600 527.240 6.740 ;
  RECT 540.320 3.600 548.320 6.740 ;
  RECT 560.160 3.600 568.160 6.740 ;
  RECT 581.240 3.600 589.240 6.740 ;
  RECT 601.080 3.600 609.080 6.740 ;
  RECT 622.160 3.600 630.160 6.740 ;
  RECT 642.000 3.600 650.000 6.740 ;
  RECT 663.080 3.600 671.080 6.740 ;
  RECT 682.920 3.600 690.920 6.740 ;
  RECT 704.000 3.600 712.000 6.740 ;
  RECT 723.840 3.600 731.840 6.740 ;
  RECT 744.920 3.600 752.920 6.740 ;
  RECT 764.760 3.600 772.760 6.740 ;
  RECT 785.840 3.600 793.840 6.740 ;
  RECT 805.680 3.600 813.680 6.740 ;
  RECT 826.760 3.600 834.760 6.740 ;
  RECT 846.600 3.600 854.600 6.740 ;
  RECT 867.680 3.600 875.680 6.740 ;
  RECT 887.520 3.600 895.520 6.740 ;
  RECT 908.600 3.600 916.600 6.740 ;
  RECT 928.440 3.600 936.440 6.740 ;
  RECT 949.520 3.600 957.520 6.740 ;
  RECT 969.360 3.600 977.360 6.740 ;
  RECT 990.440 3.600 998.440 6.740 ;
  RECT 1010.280 3.600 1018.280 6.740 ;
  RECT 1031.360 3.600 1039.360 6.740 ;
  RECT 1051.200 3.600 1059.200 6.740 ;
  RECT 1072.280 3.600 1080.280 6.740 ;
  RECT 1092.120 3.600 1100.120 6.740 ;
  RECT 1113.200 3.600 1121.200 6.740 ;
  RECT 1133.040 3.600 1141.040 6.740 ;
  RECT 1154.120 3.600 1162.120 6.740 ;
  RECT 1173.960 3.600 1181.960 6.740 ;
  RECT 1195.040 3.600 1203.040 6.740 ;
  RECT 1214.880 3.600 1222.880 6.740 ;
  RECT 1235.960 3.600 1243.960 6.740 ;
  RECT 1255.800 3.600 1263.800 6.740 ;
  RECT 1276.880 3.600 1284.880 6.740 ;
  RECT 1296.720 3.600 1304.720 6.740 ;
  RECT 2687.800 559.940 2688.660 560.320 ;
  RECT 2687.800 552.020 2688.660 552.300 ;
  RECT 2687.520 552.800 2690.940 554.000 ;
  RECT 2687.520 550.320 2690.940 551.520 ;
  RECT 2687.800 548.340 2688.660 548.620 ;
  RECT 2687.520 549.120 2690.940 550.320 ;
  RECT 2687.520 546.640 2690.940 547.840 ;
  RECT 2687.800 544.660 2688.660 544.940 ;
  RECT 2687.520 545.440 2690.940 546.640 ;
  RECT 2687.520 542.960 2690.940 544.160 ;
  RECT 2687.800 540.980 2688.660 541.260 ;
  RECT 2687.520 541.760 2690.940 542.960 ;
  RECT 2687.520 539.280 2690.940 540.480 ;
  RECT 2687.800 537.300 2688.660 537.580 ;
  RECT 2687.520 538.080 2690.940 539.280 ;
  RECT 2687.520 535.600 2690.940 536.800 ;
  RECT 2687.800 533.620 2688.660 533.900 ;
  RECT 2687.520 534.400 2690.940 535.600 ;
  RECT 2687.520 531.920 2690.940 533.120 ;
  RECT 2687.800 529.940 2688.660 530.220 ;
  RECT 2687.520 530.720 2690.940 531.920 ;
  RECT 2687.520 528.240 2690.940 529.440 ;
  RECT 2687.800 526.260 2688.660 526.540 ;
  RECT 2687.520 527.040 2690.940 528.240 ;
  RECT 2687.520 524.560 2690.940 525.760 ;
  RECT 2687.800 522.580 2688.660 522.860 ;
  RECT 2687.520 523.360 2690.940 524.560 ;
  RECT 2687.520 520.880 2690.940 522.080 ;
  RECT 2687.800 518.900 2688.660 519.180 ;
  RECT 2687.520 519.680 2690.940 520.880 ;
  RECT 2687.520 517.200 2690.940 518.400 ;
  RECT 2687.800 515.220 2688.660 515.500 ;
  RECT 2687.520 516.000 2690.940 517.200 ;
  RECT 2687.520 513.520 2690.940 514.720 ;
  RECT 2687.800 511.540 2688.660 511.820 ;
  RECT 2687.520 512.320 2690.940 513.520 ;
  RECT 2687.520 509.840 2690.940 511.040 ;
  RECT 2687.800 507.860 2688.660 508.140 ;
  RECT 2687.520 508.640 2690.940 509.840 ;
  RECT 2687.520 506.160 2690.940 507.360 ;
  RECT 2687.800 504.180 2688.660 504.460 ;
  RECT 2687.520 504.960 2690.940 506.160 ;
  RECT 2687.520 502.480 2690.940 503.680 ;
  RECT 2687.800 500.500 2688.660 500.780 ;
  RECT 2687.520 501.280 2690.940 502.480 ;
  RECT 2687.520 498.800 2690.940 500.000 ;
  RECT 2687.800 496.820 2688.660 497.100 ;
  RECT 2687.520 497.600 2690.940 498.800 ;
  RECT 2687.520 495.120 2690.940 496.320 ;
  RECT 2687.800 493.140 2688.660 493.420 ;
  RECT 2687.520 493.920 2690.940 495.120 ;
  RECT 2687.520 491.440 2690.940 492.640 ;
  RECT 2687.800 489.460 2688.660 489.740 ;
  RECT 2687.520 490.240 2690.940 491.440 ;
  RECT 2687.520 487.760 2690.940 488.960 ;
  RECT 2687.800 485.780 2688.660 486.060 ;
  RECT 2687.520 486.560 2690.940 487.760 ;
  RECT 2687.520 484.080 2690.940 485.280 ;
  RECT 2687.800 482.100 2688.660 482.380 ;
  RECT 2687.520 482.880 2690.940 484.080 ;
  RECT 2687.520 480.400 2690.940 481.600 ;
  RECT 2687.800 478.420 2688.660 478.700 ;
  RECT 2687.520 479.200 2690.940 480.400 ;
  RECT 2687.520 476.720 2690.940 477.920 ;
  RECT 2687.800 474.740 2688.660 475.020 ;
  RECT 2687.520 475.520 2690.940 476.720 ;
  RECT 2687.520 473.040 2690.940 474.240 ;
  RECT 2687.800 471.060 2688.660 471.340 ;
  RECT 2687.520 471.840 2690.940 473.040 ;
  RECT 2687.520 469.360 2690.940 470.560 ;
  RECT 2687.800 467.380 2688.660 467.660 ;
  RECT 2687.520 468.160 2690.940 469.360 ;
  RECT 2687.520 465.680 2690.940 466.880 ;
  RECT 2687.800 463.700 2688.660 463.980 ;
  RECT 2687.520 464.480 2690.940 465.680 ;
  RECT 2687.520 462.000 2690.940 463.200 ;
  RECT 2687.800 460.020 2688.660 460.300 ;
  RECT 2687.520 460.800 2690.940 462.000 ;
  RECT 2687.520 458.320 2690.940 459.520 ;
  RECT 2687.800 456.340 2688.660 456.620 ;
  RECT 2687.520 457.120 2690.940 458.320 ;
  RECT 2687.520 454.640 2690.940 455.840 ;
  RECT 2687.800 452.660 2688.660 452.940 ;
  RECT 2687.520 453.440 2690.940 454.640 ;
  RECT 2687.520 450.960 2690.940 452.160 ;
  RECT 2687.800 448.980 2688.660 449.260 ;
  RECT 2687.520 449.760 2690.940 450.960 ;
  RECT 2687.520 447.280 2690.940 448.480 ;
  RECT 2687.800 445.300 2688.660 445.580 ;
  RECT 2687.520 446.080 2690.940 447.280 ;
  RECT 2687.520 443.600 2690.940 444.800 ;
  RECT 2687.800 441.620 2688.660 441.900 ;
  RECT 2687.520 442.400 2690.940 443.600 ;
  RECT 2687.520 439.920 2690.940 441.120 ;
  RECT 2687.800 437.940 2688.660 438.220 ;
  RECT 2687.520 438.720 2690.940 439.920 ;
  RECT 2687.520 436.240 2690.940 437.440 ;
  RECT 2687.800 434.260 2688.660 434.540 ;
  RECT 2687.520 435.040 2690.940 436.240 ;
  RECT 2687.520 432.560 2690.940 433.760 ;
  RECT 2687.800 430.580 2688.660 430.860 ;
  RECT 2687.520 431.360 2690.940 432.560 ;
  RECT 2687.520 428.880 2690.940 430.080 ;
  RECT 2687.800 426.900 2688.660 427.180 ;
  RECT 2687.520 427.680 2690.940 428.880 ;
  RECT 2687.520 425.200 2690.940 426.400 ;
  RECT 2687.800 423.220 2688.660 423.500 ;
  RECT 2687.520 424.000 2690.940 425.200 ;
  RECT 2687.520 421.520 2690.940 422.720 ;
  RECT 2687.800 419.540 2688.660 419.820 ;
  RECT 2687.520 420.320 2690.940 421.520 ;
  RECT 2687.520 417.840 2690.940 419.040 ;
  RECT 2687.800 415.860 2688.660 416.140 ;
  RECT 2687.520 416.640 2690.940 417.840 ;
  RECT 2687.520 414.160 2690.940 415.360 ;
  RECT 2687.800 412.180 2688.660 412.460 ;
  RECT 2687.520 412.960 2690.940 414.160 ;
  RECT 2687.520 410.480 2690.940 411.680 ;
  RECT 2687.800 408.500 2688.660 408.780 ;
  RECT 2687.520 409.280 2690.940 410.480 ;
  RECT 2687.520 406.800 2690.940 408.000 ;
  RECT 2687.800 404.820 2688.660 405.100 ;
  RECT 2687.520 405.600 2690.940 406.800 ;
  RECT 2687.520 403.120 2690.940 404.320 ;
  RECT 2687.800 401.140 2688.660 401.420 ;
  RECT 2687.520 401.920 2690.940 403.120 ;
  RECT 2687.520 399.440 2690.940 400.640 ;
  RECT 2687.800 397.460 2688.660 397.740 ;
  RECT 2687.520 398.240 2690.940 399.440 ;
  RECT 2687.520 395.760 2690.940 396.960 ;
  RECT 2687.800 393.780 2688.660 394.060 ;
  RECT 2687.520 394.560 2690.940 395.760 ;
  RECT 2687.520 392.080 2690.940 393.280 ;
  RECT 2687.800 390.100 2688.660 390.380 ;
  RECT 2687.520 390.880 2690.940 392.080 ;
  RECT 2687.520 388.400 2690.940 389.600 ;
  RECT 2687.800 386.420 2688.660 386.700 ;
  RECT 2687.520 387.200 2690.940 388.400 ;
  RECT 2687.520 384.720 2690.940 385.920 ;
  RECT 2687.800 382.740 2688.660 383.020 ;
  RECT 2687.520 383.520 2690.940 384.720 ;
  RECT 2687.520 381.040 2690.940 382.240 ;
  RECT 2687.800 379.060 2688.660 379.340 ;
  RECT 2687.520 379.840 2690.940 381.040 ;
  RECT 2687.520 377.360 2690.940 378.560 ;
  RECT 2687.800 375.380 2688.660 375.660 ;
  RECT 2687.520 376.160 2690.940 377.360 ;
  RECT 2687.520 373.680 2690.940 374.880 ;
  RECT 2687.800 371.700 2688.660 371.980 ;
  RECT 2687.520 372.480 2690.940 373.680 ;
  RECT 2687.520 370.000 2690.940 371.200 ;
  RECT 2687.800 368.020 2688.660 368.300 ;
  RECT 2687.520 368.800 2690.940 370.000 ;
  RECT 2687.520 366.320 2690.940 367.520 ;
  RECT 2687.800 364.340 2688.660 364.620 ;
  RECT 2687.520 365.120 2690.940 366.320 ;
  RECT 2687.520 362.640 2690.940 363.840 ;
  RECT 2687.800 360.660 2688.660 360.940 ;
  RECT 2687.520 361.440 2690.940 362.640 ;
  RECT 2687.520 358.960 2690.940 360.160 ;
  RECT 2687.800 356.980 2688.660 357.260 ;
  RECT 2687.520 357.760 2690.940 358.960 ;
  RECT 2687.520 355.280 2690.940 356.480 ;
  RECT 2687.800 353.300 2688.660 353.580 ;
  RECT 2687.520 354.080 2690.940 355.280 ;
  RECT 2687.520 351.600 2690.940 352.800 ;
  RECT 2687.800 349.620 2688.660 349.900 ;
  RECT 2687.520 350.400 2690.940 351.600 ;
  RECT 2687.520 347.920 2690.940 349.120 ;
  RECT 2687.800 345.940 2688.660 346.220 ;
  RECT 2687.520 346.720 2690.940 347.920 ;
  RECT 2687.520 344.240 2690.940 345.440 ;
  RECT 2687.800 342.260 2688.660 342.540 ;
  RECT 2687.520 343.040 2690.940 344.240 ;
  RECT 2687.520 340.560 2690.940 341.760 ;
  RECT 2687.800 338.580 2688.660 338.860 ;
  RECT 2687.520 339.360 2690.940 340.560 ;
  RECT 2687.520 336.880 2690.940 338.080 ;
  RECT 2687.800 334.900 2688.660 335.180 ;
  RECT 2687.520 335.680 2690.940 336.880 ;
  RECT 2687.520 333.200 2690.940 334.400 ;
  RECT 2687.800 331.220 2688.660 331.500 ;
  RECT 2687.520 332.000 2690.940 333.200 ;
  RECT 2687.520 329.520 2690.940 330.720 ;
  RECT 2687.800 327.540 2688.660 327.820 ;
  RECT 2687.520 328.320 2690.940 329.520 ;
  RECT 2687.520 325.840 2690.940 327.040 ;
  RECT 2687.800 323.860 2688.660 324.140 ;
  RECT 2687.520 324.640 2690.940 325.840 ;
  RECT 2687.520 322.160 2690.940 323.360 ;
  RECT 2687.800 320.180 2688.660 320.460 ;
  RECT 2687.520 320.960 2690.940 322.160 ;
  RECT 2687.520 318.480 2690.940 319.680 ;
  RECT 2687.800 316.500 2688.660 316.780 ;
  RECT 2687.520 317.280 2690.940 318.480 ;
  RECT 2687.520 314.800 2690.940 316.000 ;
  RECT 2687.800 312.820 2688.660 313.100 ;
  RECT 2687.520 313.600 2690.940 314.800 ;
  RECT 2687.520 311.120 2690.940 312.320 ;
  RECT 2687.800 309.140 2688.660 309.420 ;
  RECT 2687.520 309.920 2690.940 311.120 ;
  RECT 2687.520 307.440 2690.940 308.640 ;
  RECT 2687.800 305.460 2688.660 305.740 ;
  RECT 2687.520 306.240 2690.940 307.440 ;
  RECT 2687.520 303.760 2690.940 304.960 ;
  RECT 2687.800 301.780 2688.660 302.060 ;
  RECT 2687.520 302.560 2690.940 303.760 ;
  RECT 2687.520 300.080 2690.940 301.280 ;
  RECT 2687.800 298.100 2688.660 298.380 ;
  RECT 2687.520 298.880 2690.940 300.080 ;
  RECT 2687.520 296.400 2690.940 297.600 ;
  RECT 2687.800 294.420 2688.660 294.700 ;
  RECT 2687.520 295.200 2690.940 296.400 ;
  RECT 2687.520 292.720 2690.940 293.920 ;
  RECT 2687.800 290.740 2688.660 291.020 ;
  RECT 2687.520 291.520 2690.940 292.720 ;
  RECT 2687.520 289.040 2690.940 290.240 ;
  RECT 2687.800 287.060 2688.660 287.340 ;
  RECT 2687.520 287.840 2690.940 289.040 ;
  RECT 2687.520 285.360 2690.940 286.560 ;
  RECT 2687.800 283.380 2688.660 283.660 ;
  RECT 2687.520 284.160 2690.940 285.360 ;
  RECT 2687.520 281.680 2690.940 282.880 ;
  RECT 2687.800 279.700 2688.660 279.980 ;
  RECT 2687.520 280.480 2690.940 281.680 ;
  RECT 2687.520 278.000 2690.940 279.200 ;
  RECT 2687.800 276.020 2688.660 276.300 ;
  RECT 2687.520 276.800 2690.940 278.000 ;
  RECT 2687.520 274.320 2690.940 275.520 ;
  RECT 2687.800 272.340 2688.660 272.620 ;
  RECT 2687.520 273.120 2690.940 274.320 ;
  RECT 2687.520 270.640 2690.940 271.840 ;
  RECT 2687.800 268.660 2688.660 268.940 ;
  RECT 2687.520 269.440 2690.940 270.640 ;
  RECT 2687.520 266.960 2690.940 268.160 ;
  RECT 2687.800 264.980 2688.660 265.260 ;
  RECT 2687.520 265.760 2690.940 266.960 ;
  RECT 2687.520 263.280 2690.940 264.480 ;
  RECT 2687.800 261.300 2688.660 261.580 ;
  RECT 2687.520 262.080 2690.940 263.280 ;
  RECT 2687.520 259.600 2690.940 260.800 ;
  RECT 2687.800 257.620 2688.660 257.900 ;
  RECT 2687.520 258.400 2690.940 259.600 ;
  RECT 2687.520 255.920 2690.940 257.120 ;
  RECT 2687.800 253.940 2688.660 254.220 ;
  RECT 2687.520 254.720 2690.940 255.920 ;
  RECT 2687.520 252.240 2690.940 253.440 ;
  RECT 2687.800 250.260 2688.660 250.540 ;
  RECT 2687.520 251.040 2690.940 252.240 ;
  RECT 2687.520 248.560 2690.940 249.760 ;
  RECT 2687.800 246.580 2688.660 246.860 ;
  RECT 2687.520 247.360 2690.940 248.560 ;
  RECT 2687.520 244.880 2690.940 246.080 ;
  RECT 2687.800 242.900 2688.660 243.180 ;
  RECT 2687.520 243.680 2690.940 244.880 ;
  RECT 2687.520 241.200 2690.940 242.400 ;
  RECT 2687.800 239.220 2688.660 239.500 ;
  RECT 2687.520 240.000 2690.940 241.200 ;
  RECT 2687.520 237.520 2690.940 238.720 ;
  RECT 2687.800 235.540 2688.660 235.820 ;
  RECT 2687.520 236.320 2690.940 237.520 ;
  RECT 2687.520 233.840 2690.940 235.040 ;
  RECT 2687.800 231.860 2688.660 232.140 ;
  RECT 2687.520 232.640 2690.940 233.840 ;
  RECT 2687.520 230.160 2690.940 231.360 ;
  RECT 2687.800 228.180 2688.660 228.460 ;
  RECT 2687.520 228.960 2690.940 230.160 ;
  RECT 2687.520 226.480 2690.940 227.680 ;
  RECT 2687.800 224.500 2688.660 224.780 ;
  RECT 2687.520 225.280 2690.940 226.480 ;
  RECT 2687.520 222.800 2690.940 224.000 ;
  RECT 2687.800 220.820 2688.660 221.100 ;
  RECT 2687.520 221.600 2690.940 222.800 ;
  RECT 2687.520 219.120 2690.940 220.320 ;
  RECT 2687.800 217.140 2688.660 217.420 ;
  RECT 2687.520 217.920 2690.940 219.120 ;
  RECT 2687.520 215.440 2690.940 216.640 ;
  RECT 2687.800 213.460 2688.660 213.740 ;
  RECT 2687.520 214.240 2690.940 215.440 ;
  RECT 2687.520 211.760 2690.940 212.960 ;
  RECT 2687.800 209.780 2688.660 210.060 ;
  RECT 2687.520 210.560 2690.940 211.760 ;
  RECT 2687.520 208.080 2690.940 209.280 ;
  RECT 2687.800 206.100 2688.660 206.380 ;
  RECT 2687.520 206.880 2690.940 208.080 ;
  RECT 2687.520 204.400 2690.940 205.600 ;
  RECT 2687.800 202.420 2688.660 202.700 ;
  RECT 2687.520 203.200 2690.940 204.400 ;
  RECT 2687.520 200.720 2690.940 201.920 ;
  RECT 2687.800 198.740 2688.660 199.020 ;
  RECT 2687.520 199.520 2690.940 200.720 ;
  RECT 2687.520 197.040 2690.940 198.240 ;
  RECT 2687.800 195.060 2688.660 195.340 ;
  RECT 2687.520 195.840 2690.940 197.040 ;
  RECT 2687.520 193.360 2690.940 194.560 ;
  RECT 2687.800 191.380 2688.660 191.660 ;
  RECT 2687.520 192.160 2690.940 193.360 ;
  RECT 2687.520 189.680 2690.940 190.880 ;
  RECT 2687.800 187.700 2688.660 187.980 ;
  RECT 2687.520 188.480 2690.940 189.680 ;
  RECT 2687.520 186.000 2690.940 187.200 ;
  RECT 2687.800 184.020 2688.660 184.300 ;
  RECT 2687.520 184.800 2690.940 186.000 ;
  RECT 2687.520 182.320 2690.940 183.520 ;
  RECT 2687.800 180.340 2688.660 180.620 ;
  RECT 2687.520 181.120 2690.940 182.320 ;
  RECT 2687.520 178.640 2690.940 179.840 ;
  RECT 2687.800 176.660 2688.660 176.940 ;
  RECT 2687.520 177.440 2690.940 178.640 ;
  RECT 2687.520 174.960 2690.940 176.160 ;
  RECT 2687.800 172.980 2688.660 173.260 ;
  RECT 2687.520 173.760 2690.940 174.960 ;
  RECT 2687.520 171.280 2690.940 172.480 ;
  RECT 2687.800 169.300 2688.660 169.580 ;
  RECT 2687.520 170.080 2690.940 171.280 ;
  RECT 2687.520 167.600 2690.940 168.800 ;
  RECT 2687.800 165.620 2688.660 165.900 ;
  RECT 2687.520 166.400 2690.940 167.600 ;
  RECT 2687.520 163.920 2690.940 165.120 ;
  RECT 2687.800 161.940 2688.660 162.220 ;
  RECT 2687.520 162.720 2690.940 163.920 ;
  RECT 2687.520 160.240 2690.940 161.440 ;
  RECT 2687.800 158.260 2688.660 158.540 ;
  RECT 2687.520 159.040 2690.940 160.240 ;
  RECT 2687.520 156.560 2690.940 157.760 ;
  RECT 2687.800 154.580 2688.660 154.860 ;
  RECT 2687.520 155.360 2690.940 156.560 ;
  RECT 2687.520 152.880 2690.940 154.080 ;
  RECT 2687.800 150.900 2688.660 151.180 ;
  RECT 2687.520 151.680 2690.940 152.880 ;
  RECT 2687.520 149.200 2690.940 150.400 ;
  RECT 2687.800 147.220 2688.660 147.500 ;
  RECT 2687.520 148.000 2690.940 149.200 ;
  RECT 2687.520 145.520 2690.940 146.720 ;
  RECT 2687.800 143.540 2688.660 143.820 ;
  RECT 2687.520 144.320 2690.940 145.520 ;
  RECT 2687.520 141.840 2690.940 143.040 ;
  RECT 2687.800 139.860 2688.660 140.140 ;
  RECT 2687.520 140.640 2690.940 141.840 ;
  RECT 2687.520 138.160 2690.940 139.360 ;
  RECT 2687.800 136.180 2688.660 136.460 ;
  RECT 2687.520 136.960 2690.940 138.160 ;
  RECT 2687.520 134.480 2690.940 135.680 ;
  RECT 2687.800 132.500 2688.660 132.780 ;
  RECT 2687.520 133.280 2690.940 134.480 ;
  RECT 2687.520 130.800 2690.940 132.000 ;
  RECT 2687.800 128.820 2688.660 129.100 ;
  RECT 2687.520 129.600 2690.940 130.800 ;
  RECT 2687.520 127.120 2690.940 128.320 ;
  RECT 2687.800 125.140 2688.660 125.420 ;
  RECT 2687.520 125.920 2690.940 127.120 ;
  RECT 2687.520 123.440 2690.940 124.640 ;
  RECT 2687.800 121.460 2688.660 121.740 ;
  RECT 2687.520 122.240 2690.940 123.440 ;
  RECT 2687.520 119.760 2690.940 120.960 ;
  RECT 2687.800 117.780 2688.660 118.060 ;
  RECT 2687.520 118.560 2690.940 119.760 ;
  RECT 2687.520 116.080 2690.940 117.280 ;
  RECT 2687.800 114.100 2688.660 114.380 ;
  RECT 2687.520 114.880 2690.940 116.080 ;
  RECT 2687.520 112.400 2690.940 113.600 ;
  RECT 2687.800 110.420 2688.660 110.700 ;
  RECT 2687.520 111.200 2690.940 112.400 ;
  RECT 2687.520 108.720 2690.940 109.920 ;
  RECT 2687.800 106.740 2688.660 107.020 ;
  RECT 2687.520 107.520 2690.940 108.720 ;
  RECT 2687.520 105.040 2690.940 106.240 ;
  RECT 2687.800 103.060 2688.660 103.340 ;
  RECT 2687.520 103.840 2690.940 105.040 ;
  RECT 2687.520 101.360 2690.940 102.560 ;
  RECT 2687.800 99.380 2688.660 99.660 ;
  RECT 2687.520 100.160 2690.940 101.360 ;
  RECT 2687.520 97.680 2690.940 98.880 ;
  RECT 2687.800 95.700 2688.660 95.980 ;
  RECT 2687.520 96.480 2690.940 97.680 ;
  RECT 2687.520 94.000 2690.940 95.200 ;
  RECT 2687.800 92.020 2688.660 92.300 ;
  RECT 2687.520 92.800 2690.940 94.000 ;
  RECT 2687.520 90.320 2690.940 91.520 ;
  RECT 2687.800 88.340 2688.660 88.620 ;
  RECT 2687.520 89.120 2690.940 90.320 ;
  RECT 2687.520 86.640 2690.940 87.840 ;
  RECT 2687.800 84.660 2688.660 84.940 ;
  RECT 2687.520 85.440 2690.940 86.640 ;
  RECT 2687.520 82.960 2690.940 84.160 ;
  RECT 2687.800 80.980 2688.660 81.260 ;
  RECT 2687.520 81.760 2690.940 82.960 ;
  RECT 2687.520 79.280 2690.940 80.480 ;
  RECT 2687.800 77.300 2688.660 77.580 ;
  RECT 2687.520 78.080 2690.940 79.280 ;
  RECT 2687.520 75.600 2690.940 76.800 ;
  RECT 2687.800 73.620 2688.660 73.900 ;
  RECT 2687.520 74.400 2690.940 75.600 ;
  RECT 2687.520 71.920 2690.940 73.120 ;
  RECT 2687.800 69.940 2688.660 70.220 ;
  RECT 2687.520 70.720 2690.940 71.920 ;
  RECT 2687.520 68.240 2690.940 69.440 ;
  RECT 2687.800 65.600 2688.660 65.980 ;
  RECT 1376.250 560.510 1376.500 563.930 ;
  RECT 1376.820 560.790 1377.070 561.650 ;
  RECT 1417.170 560.510 1417.420 563.930 ;
  RECT 1417.740 560.790 1417.990 561.650 ;
  RECT 1458.090 560.510 1458.340 563.930 ;
  RECT 1458.660 560.790 1458.910 561.650 ;
  RECT 1499.010 560.510 1499.260 563.930 ;
  RECT 1499.580 560.790 1499.830 561.650 ;
  RECT 1539.930 560.510 1540.180 563.930 ;
  RECT 1540.500 560.790 1540.750 561.650 ;
  RECT 1580.850 560.510 1581.100 563.930 ;
  RECT 1581.420 560.790 1581.670 561.650 ;
  RECT 1621.770 560.510 1622.020 563.930 ;
  RECT 1622.340 560.790 1622.590 561.650 ;
  RECT 1662.690 560.510 1662.940 563.930 ;
  RECT 1663.260 560.790 1663.510 561.650 ;
  RECT 1703.610 560.510 1703.860 563.930 ;
  RECT 1704.180 560.790 1704.430 561.650 ;
  RECT 1744.530 560.510 1744.780 563.930 ;
  RECT 1745.100 560.790 1745.350 561.650 ;
  RECT 1785.450 560.510 1785.700 563.930 ;
  RECT 1786.020 560.790 1786.270 561.650 ;
  RECT 1826.370 560.510 1826.620 563.930 ;
  RECT 1826.940 560.790 1827.190 561.650 ;
  RECT 1867.290 560.510 1867.540 563.930 ;
  RECT 1867.860 560.790 1868.110 561.650 ;
  RECT 1908.210 560.510 1908.460 563.930 ;
  RECT 1908.780 560.790 1909.030 561.650 ;
  RECT 1949.130 560.510 1949.380 563.930 ;
  RECT 1949.700 560.790 1949.950 561.650 ;
  RECT 1990.050 560.510 1990.300 563.930 ;
  RECT 1990.620 560.790 1990.870 561.650 ;
  RECT 2030.970 560.510 2031.220 563.930 ;
  RECT 2031.540 560.790 2031.790 561.650 ;
  RECT 2071.890 560.510 2072.140 563.930 ;
  RECT 2072.460 560.790 2072.710 561.650 ;
  RECT 2112.810 560.510 2113.060 563.930 ;
  RECT 2113.380 560.790 2113.630 561.650 ;
  RECT 2153.730 560.510 2153.980 563.930 ;
  RECT 2154.300 560.790 2154.550 561.650 ;
  RECT 2194.650 560.510 2194.900 563.930 ;
  RECT 2195.220 560.790 2195.470 561.650 ;
  RECT 2235.570 560.510 2235.820 563.930 ;
  RECT 2236.140 560.790 2236.390 561.650 ;
  RECT 2276.490 560.510 2276.740 563.930 ;
  RECT 2277.060 560.790 2277.310 561.650 ;
  RECT 2317.410 560.510 2317.660 563.930 ;
  RECT 2317.980 560.790 2318.230 561.650 ;
  RECT 2358.330 560.510 2358.580 563.930 ;
  RECT 2358.900 560.790 2359.150 561.650 ;
  RECT 2399.250 560.510 2399.500 563.930 ;
  RECT 2399.820 560.790 2400.070 561.650 ;
  RECT 2440.170 560.510 2440.420 563.930 ;
  RECT 2440.740 560.790 2440.990 561.650 ;
  RECT 2481.090 560.510 2481.340 563.930 ;
  RECT 2481.660 560.790 2481.910 561.650 ;
  RECT 2522.010 560.510 2522.260 563.930 ;
  RECT 2522.580 560.790 2522.830 561.650 ;
  RECT 2562.930 560.510 2563.180 563.930 ;
  RECT 2563.500 560.790 2563.750 561.650 ;
  RECT 2603.850 560.510 2604.100 563.930 ;
  RECT 2604.420 560.790 2604.670 561.650 ;
  RECT 2644.770 560.510 2645.020 563.930 ;
  RECT 2645.340 560.790 2645.590 561.650 ;
  RECT 1372.760 560.510 1373.660 563.930 ;
  RECT 1343.440 560.510 1346.630 563.930 ;
  RECT 1353.440 560.510 1357.760 563.930 ;
  RECT 1359.810 560.790 1362.320 561.650 ;
  RECT 1347.390 560.790 1349.780 561.650 ;
  RECT 1339.880 560.790 1342.940 561.650 ;
  RECT 1364.060 560.790 1366.910 561.650 ;
  RECT 1368.360 560.790 1371.610 561.650 ;
  RECT 1335.160 560.510 1336.920 563.930 ;
  RECT 1337.160 560.790 1338.920 561.650 ;
  RECT 1317.900 560.510 1319.580 563.930 ;
  RECT 1321.820 560.510 1323.580 563.930 ;
  RECT 1325.820 560.510 1327.580 563.930 ;
  RECT 1329.820 560.510 1331.580 563.930 ;
  RECT 1319.820 560.790 1321.580 561.650 ;
  RECT 1323.820 560.790 1325.580 561.650 ;
  RECT 1327.820 560.790 1329.580 561.650 ;
  RECT 1331.820 560.790 1333.580 561.650 ;
  RECT 1316.800 560.510 1317.700 563.930 ;
  RECT 4.280 65.600 5.140 65.980 ;
  RECT 2.000 68.240 5.420 69.440 ;
  RECT 2.000 70.720 5.420 71.920 ;
  RECT 4.280 69.940 5.140 70.220 ;
  RECT 2.000 71.920 5.420 73.120 ;
  RECT 2.000 74.400 5.420 75.600 ;
  RECT 4.280 73.620 5.140 73.900 ;
  RECT 2.000 75.600 5.420 76.800 ;
  RECT 2.000 78.080 5.420 79.280 ;
  RECT 4.280 77.300 5.140 77.580 ;
  RECT 2.000 79.280 5.420 80.480 ;
  RECT 2.000 81.760 5.420 82.960 ;
  RECT 4.280 80.980 5.140 81.260 ;
  RECT 2.000 82.960 5.420 84.160 ;
  RECT 2.000 85.440 5.420 86.640 ;
  RECT 4.280 84.660 5.140 84.940 ;
  RECT 2.000 86.640 5.420 87.840 ;
  RECT 2.000 89.120 5.420 90.320 ;
  RECT 4.280 88.340 5.140 88.620 ;
  RECT 2.000 90.320 5.420 91.520 ;
  RECT 2.000 92.800 5.420 94.000 ;
  RECT 4.280 92.020 5.140 92.300 ;
  RECT 2.000 94.000 5.420 95.200 ;
  RECT 2.000 96.480 5.420 97.680 ;
  RECT 4.280 95.700 5.140 95.980 ;
  RECT 2.000 97.680 5.420 98.880 ;
  RECT 2.000 100.160 5.420 101.360 ;
  RECT 4.280 99.380 5.140 99.660 ;
  RECT 2.000 101.360 5.420 102.560 ;
  RECT 2.000 103.840 5.420 105.040 ;
  RECT 4.280 103.060 5.140 103.340 ;
  RECT 2.000 105.040 5.420 106.240 ;
  RECT 2.000 107.520 5.420 108.720 ;
  RECT 4.280 106.740 5.140 107.020 ;
  RECT 2.000 108.720 5.420 109.920 ;
  RECT 2.000 111.200 5.420 112.400 ;
  RECT 4.280 110.420 5.140 110.700 ;
  RECT 2.000 112.400 5.420 113.600 ;
  RECT 2.000 114.880 5.420 116.080 ;
  RECT 4.280 114.100 5.140 114.380 ;
  RECT 2.000 116.080 5.420 117.280 ;
  RECT 2.000 118.560 5.420 119.760 ;
  RECT 4.280 117.780 5.140 118.060 ;
  RECT 2.000 119.760 5.420 120.960 ;
  RECT 2.000 122.240 5.420 123.440 ;
  RECT 4.280 121.460 5.140 121.740 ;
  RECT 2.000 123.440 5.420 124.640 ;
  RECT 2.000 125.920 5.420 127.120 ;
  RECT 4.280 125.140 5.140 125.420 ;
  RECT 2.000 127.120 5.420 128.320 ;
  RECT 2.000 129.600 5.420 130.800 ;
  RECT 4.280 128.820 5.140 129.100 ;
  RECT 2.000 130.800 5.420 132.000 ;
  RECT 2.000 133.280 5.420 134.480 ;
  RECT 4.280 132.500 5.140 132.780 ;
  RECT 2.000 134.480 5.420 135.680 ;
  RECT 2.000 136.960 5.420 138.160 ;
  RECT 4.280 136.180 5.140 136.460 ;
  RECT 2.000 138.160 5.420 139.360 ;
  RECT 2.000 140.640 5.420 141.840 ;
  RECT 4.280 139.860 5.140 140.140 ;
  RECT 2.000 141.840 5.420 143.040 ;
  RECT 2.000 144.320 5.420 145.520 ;
  RECT 4.280 143.540 5.140 143.820 ;
  RECT 2.000 145.520 5.420 146.720 ;
  RECT 2.000 148.000 5.420 149.200 ;
  RECT 4.280 147.220 5.140 147.500 ;
  RECT 2.000 149.200 5.420 150.400 ;
  RECT 2.000 151.680 5.420 152.880 ;
  RECT 4.280 150.900 5.140 151.180 ;
  RECT 2.000 152.880 5.420 154.080 ;
  RECT 2.000 155.360 5.420 156.560 ;
  RECT 4.280 154.580 5.140 154.860 ;
  RECT 2.000 156.560 5.420 157.760 ;
  RECT 2.000 159.040 5.420 160.240 ;
  RECT 4.280 158.260 5.140 158.540 ;
  RECT 2.000 160.240 5.420 161.440 ;
  RECT 2.000 162.720 5.420 163.920 ;
  RECT 4.280 161.940 5.140 162.220 ;
  RECT 2.000 163.920 5.420 165.120 ;
  RECT 2.000 166.400 5.420 167.600 ;
  RECT 4.280 165.620 5.140 165.900 ;
  RECT 2.000 167.600 5.420 168.800 ;
  RECT 2.000 170.080 5.420 171.280 ;
  RECT 4.280 169.300 5.140 169.580 ;
  RECT 2.000 171.280 5.420 172.480 ;
  RECT 2.000 173.760 5.420 174.960 ;
  RECT 4.280 172.980 5.140 173.260 ;
  RECT 2.000 174.960 5.420 176.160 ;
  RECT 2.000 177.440 5.420 178.640 ;
  RECT 4.280 176.660 5.140 176.940 ;
  RECT 2.000 178.640 5.420 179.840 ;
  RECT 2.000 181.120 5.420 182.320 ;
  RECT 4.280 180.340 5.140 180.620 ;
  RECT 2.000 182.320 5.420 183.520 ;
  RECT 2.000 184.800 5.420 186.000 ;
  RECT 4.280 184.020 5.140 184.300 ;
  RECT 2.000 186.000 5.420 187.200 ;
  RECT 2.000 188.480 5.420 189.680 ;
  RECT 4.280 187.700 5.140 187.980 ;
  RECT 2.000 189.680 5.420 190.880 ;
  RECT 2.000 192.160 5.420 193.360 ;
  RECT 4.280 191.380 5.140 191.660 ;
  RECT 2.000 193.360 5.420 194.560 ;
  RECT 2.000 195.840 5.420 197.040 ;
  RECT 4.280 195.060 5.140 195.340 ;
  RECT 2.000 197.040 5.420 198.240 ;
  RECT 2.000 199.520 5.420 200.720 ;
  RECT 4.280 198.740 5.140 199.020 ;
  RECT 2.000 200.720 5.420 201.920 ;
  RECT 2.000 203.200 5.420 204.400 ;
  RECT 4.280 202.420 5.140 202.700 ;
  RECT 2.000 204.400 5.420 205.600 ;
  RECT 2.000 206.880 5.420 208.080 ;
  RECT 4.280 206.100 5.140 206.380 ;
  RECT 2.000 208.080 5.420 209.280 ;
  RECT 2.000 210.560 5.420 211.760 ;
  RECT 4.280 209.780 5.140 210.060 ;
  RECT 2.000 211.760 5.420 212.960 ;
  RECT 2.000 214.240 5.420 215.440 ;
  RECT 4.280 213.460 5.140 213.740 ;
  RECT 2.000 215.440 5.420 216.640 ;
  RECT 2.000 217.920 5.420 219.120 ;
  RECT 4.280 217.140 5.140 217.420 ;
  RECT 2.000 219.120 5.420 220.320 ;
  RECT 2.000 221.600 5.420 222.800 ;
  RECT 4.280 220.820 5.140 221.100 ;
  RECT 2.000 222.800 5.420 224.000 ;
  RECT 2.000 225.280 5.420 226.480 ;
  RECT 4.280 224.500 5.140 224.780 ;
  RECT 2.000 226.480 5.420 227.680 ;
  RECT 2.000 228.960 5.420 230.160 ;
  RECT 4.280 228.180 5.140 228.460 ;
  RECT 2.000 230.160 5.420 231.360 ;
  RECT 2.000 232.640 5.420 233.840 ;
  RECT 4.280 231.860 5.140 232.140 ;
  RECT 2.000 233.840 5.420 235.040 ;
  RECT 2.000 236.320 5.420 237.520 ;
  RECT 4.280 235.540 5.140 235.820 ;
  RECT 2.000 237.520 5.420 238.720 ;
  RECT 2.000 240.000 5.420 241.200 ;
  RECT 4.280 239.220 5.140 239.500 ;
  RECT 2.000 241.200 5.420 242.400 ;
  RECT 2.000 243.680 5.420 244.880 ;
  RECT 4.280 242.900 5.140 243.180 ;
  RECT 2.000 244.880 5.420 246.080 ;
  RECT 2.000 247.360 5.420 248.560 ;
  RECT 4.280 246.580 5.140 246.860 ;
  RECT 2.000 248.560 5.420 249.760 ;
  RECT 2.000 251.040 5.420 252.240 ;
  RECT 4.280 250.260 5.140 250.540 ;
  RECT 2.000 252.240 5.420 253.440 ;
  RECT 2.000 254.720 5.420 255.920 ;
  RECT 4.280 253.940 5.140 254.220 ;
  RECT 2.000 255.920 5.420 257.120 ;
  RECT 2.000 258.400 5.420 259.600 ;
  RECT 4.280 257.620 5.140 257.900 ;
  RECT 2.000 259.600 5.420 260.800 ;
  RECT 2.000 262.080 5.420 263.280 ;
  RECT 4.280 261.300 5.140 261.580 ;
  RECT 2.000 263.280 5.420 264.480 ;
  RECT 2.000 265.760 5.420 266.960 ;
  RECT 4.280 264.980 5.140 265.260 ;
  RECT 2.000 266.960 5.420 268.160 ;
  RECT 2.000 269.440 5.420 270.640 ;
  RECT 4.280 268.660 5.140 268.940 ;
  RECT 2.000 270.640 5.420 271.840 ;
  RECT 2.000 273.120 5.420 274.320 ;
  RECT 4.280 272.340 5.140 272.620 ;
  RECT 2.000 274.320 5.420 275.520 ;
  RECT 2.000 276.800 5.420 278.000 ;
  RECT 4.280 276.020 5.140 276.300 ;
  RECT 2.000 278.000 5.420 279.200 ;
  RECT 2.000 280.480 5.420 281.680 ;
  RECT 4.280 279.700 5.140 279.980 ;
  RECT 2.000 281.680 5.420 282.880 ;
  RECT 2.000 284.160 5.420 285.360 ;
  RECT 4.280 283.380 5.140 283.660 ;
  RECT 2.000 285.360 5.420 286.560 ;
  RECT 2.000 287.840 5.420 289.040 ;
  RECT 4.280 287.060 5.140 287.340 ;
  RECT 2.000 289.040 5.420 290.240 ;
  RECT 2.000 291.520 5.420 292.720 ;
  RECT 4.280 290.740 5.140 291.020 ;
  RECT 2.000 292.720 5.420 293.920 ;
  RECT 2.000 295.200 5.420 296.400 ;
  RECT 4.280 294.420 5.140 294.700 ;
  RECT 2.000 296.400 5.420 297.600 ;
  RECT 2.000 298.880 5.420 300.080 ;
  RECT 4.280 298.100 5.140 298.380 ;
  RECT 2.000 300.080 5.420 301.280 ;
  RECT 2.000 302.560 5.420 303.760 ;
  RECT 4.280 301.780 5.140 302.060 ;
  RECT 2.000 303.760 5.420 304.960 ;
  RECT 2.000 306.240 5.420 307.440 ;
  RECT 4.280 305.460 5.140 305.740 ;
  RECT 2.000 307.440 5.420 308.640 ;
  RECT 2.000 309.920 5.420 311.120 ;
  RECT 4.280 309.140 5.140 309.420 ;
  RECT 2.000 311.120 5.420 312.320 ;
  RECT 2.000 313.600 5.420 314.800 ;
  RECT 4.280 312.820 5.140 313.100 ;
  RECT 2.000 314.800 5.420 316.000 ;
  RECT 2.000 317.280 5.420 318.480 ;
  RECT 4.280 316.500 5.140 316.780 ;
  RECT 2.000 318.480 5.420 319.680 ;
  RECT 2.000 320.960 5.420 322.160 ;
  RECT 4.280 320.180 5.140 320.460 ;
  RECT 2.000 322.160 5.420 323.360 ;
  RECT 2.000 324.640 5.420 325.840 ;
  RECT 4.280 323.860 5.140 324.140 ;
  RECT 2.000 325.840 5.420 327.040 ;
  RECT 2.000 328.320 5.420 329.520 ;
  RECT 4.280 327.540 5.140 327.820 ;
  RECT 2.000 329.520 5.420 330.720 ;
  RECT 2.000 332.000 5.420 333.200 ;
  RECT 4.280 331.220 5.140 331.500 ;
  RECT 2.000 333.200 5.420 334.400 ;
  RECT 2.000 335.680 5.420 336.880 ;
  RECT 4.280 334.900 5.140 335.180 ;
  RECT 2.000 336.880 5.420 338.080 ;
  RECT 2.000 339.360 5.420 340.560 ;
  RECT 4.280 338.580 5.140 338.860 ;
  RECT 2.000 340.560 5.420 341.760 ;
  RECT 2.000 343.040 5.420 344.240 ;
  RECT 4.280 342.260 5.140 342.540 ;
  RECT 2.000 344.240 5.420 345.440 ;
  RECT 2.000 346.720 5.420 347.920 ;
  RECT 4.280 345.940 5.140 346.220 ;
  RECT 2.000 347.920 5.420 349.120 ;
  RECT 2.000 350.400 5.420 351.600 ;
  RECT 4.280 349.620 5.140 349.900 ;
  RECT 2.000 351.600 5.420 352.800 ;
  RECT 2.000 354.080 5.420 355.280 ;
  RECT 4.280 353.300 5.140 353.580 ;
  RECT 2.000 355.280 5.420 356.480 ;
  RECT 2.000 357.760 5.420 358.960 ;
  RECT 4.280 356.980 5.140 357.260 ;
  RECT 2.000 358.960 5.420 360.160 ;
  RECT 2.000 361.440 5.420 362.640 ;
  RECT 4.280 360.660 5.140 360.940 ;
  RECT 2.000 362.640 5.420 363.840 ;
  RECT 2.000 365.120 5.420 366.320 ;
  RECT 4.280 364.340 5.140 364.620 ;
  RECT 2.000 366.320 5.420 367.520 ;
  RECT 2.000 368.800 5.420 370.000 ;
  RECT 4.280 368.020 5.140 368.300 ;
  RECT 2.000 370.000 5.420 371.200 ;
  RECT 2.000 372.480 5.420 373.680 ;
  RECT 4.280 371.700 5.140 371.980 ;
  RECT 2.000 373.680 5.420 374.880 ;
  RECT 2.000 376.160 5.420 377.360 ;
  RECT 4.280 375.380 5.140 375.660 ;
  RECT 2.000 377.360 5.420 378.560 ;
  RECT 2.000 379.840 5.420 381.040 ;
  RECT 4.280 379.060 5.140 379.340 ;
  RECT 2.000 381.040 5.420 382.240 ;
  RECT 2.000 383.520 5.420 384.720 ;
  RECT 4.280 382.740 5.140 383.020 ;
  RECT 2.000 384.720 5.420 385.920 ;
  RECT 2.000 387.200 5.420 388.400 ;
  RECT 4.280 386.420 5.140 386.700 ;
  RECT 2.000 388.400 5.420 389.600 ;
  RECT 2.000 390.880 5.420 392.080 ;
  RECT 4.280 390.100 5.140 390.380 ;
  RECT 2.000 392.080 5.420 393.280 ;
  RECT 2.000 394.560 5.420 395.760 ;
  RECT 4.280 393.780 5.140 394.060 ;
  RECT 2.000 395.760 5.420 396.960 ;
  RECT 2.000 398.240 5.420 399.440 ;
  RECT 4.280 397.460 5.140 397.740 ;
  RECT 2.000 399.440 5.420 400.640 ;
  RECT 2.000 401.920 5.420 403.120 ;
  RECT 4.280 401.140 5.140 401.420 ;
  RECT 2.000 403.120 5.420 404.320 ;
  RECT 2.000 405.600 5.420 406.800 ;
  RECT 4.280 404.820 5.140 405.100 ;
  RECT 2.000 406.800 5.420 408.000 ;
  RECT 2.000 409.280 5.420 410.480 ;
  RECT 4.280 408.500 5.140 408.780 ;
  RECT 2.000 410.480 5.420 411.680 ;
  RECT 2.000 412.960 5.420 414.160 ;
  RECT 4.280 412.180 5.140 412.460 ;
  RECT 2.000 414.160 5.420 415.360 ;
  RECT 2.000 416.640 5.420 417.840 ;
  RECT 4.280 415.860 5.140 416.140 ;
  RECT 2.000 417.840 5.420 419.040 ;
  RECT 2.000 420.320 5.420 421.520 ;
  RECT 4.280 419.540 5.140 419.820 ;
  RECT 2.000 421.520 5.420 422.720 ;
  RECT 2.000 424.000 5.420 425.200 ;
  RECT 4.280 423.220 5.140 423.500 ;
  RECT 2.000 425.200 5.420 426.400 ;
  RECT 2.000 427.680 5.420 428.880 ;
  RECT 4.280 426.900 5.140 427.180 ;
  RECT 2.000 428.880 5.420 430.080 ;
  RECT 2.000 431.360 5.420 432.560 ;
  RECT 4.280 430.580 5.140 430.860 ;
  RECT 2.000 432.560 5.420 433.760 ;
  RECT 2.000 435.040 5.420 436.240 ;
  RECT 4.280 434.260 5.140 434.540 ;
  RECT 2.000 436.240 5.420 437.440 ;
  RECT 2.000 438.720 5.420 439.920 ;
  RECT 4.280 437.940 5.140 438.220 ;
  RECT 2.000 439.920 5.420 441.120 ;
  RECT 2.000 442.400 5.420 443.600 ;
  RECT 4.280 441.620 5.140 441.900 ;
  RECT 2.000 443.600 5.420 444.800 ;
  RECT 2.000 446.080 5.420 447.280 ;
  RECT 4.280 445.300 5.140 445.580 ;
  RECT 2.000 447.280 5.420 448.480 ;
  RECT 2.000 449.760 5.420 450.960 ;
  RECT 4.280 448.980 5.140 449.260 ;
  RECT 2.000 450.960 5.420 452.160 ;
  RECT 2.000 453.440 5.420 454.640 ;
  RECT 4.280 452.660 5.140 452.940 ;
  RECT 2.000 454.640 5.420 455.840 ;
  RECT 2.000 457.120 5.420 458.320 ;
  RECT 4.280 456.340 5.140 456.620 ;
  RECT 2.000 458.320 5.420 459.520 ;
  RECT 2.000 460.800 5.420 462.000 ;
  RECT 4.280 460.020 5.140 460.300 ;
  RECT 2.000 462.000 5.420 463.200 ;
  RECT 2.000 464.480 5.420 465.680 ;
  RECT 4.280 463.700 5.140 463.980 ;
  RECT 2.000 465.680 5.420 466.880 ;
  RECT 2.000 468.160 5.420 469.360 ;
  RECT 4.280 467.380 5.140 467.660 ;
  RECT 2.000 469.360 5.420 470.560 ;
  RECT 2.000 471.840 5.420 473.040 ;
  RECT 4.280 471.060 5.140 471.340 ;
  RECT 2.000 473.040 5.420 474.240 ;
  RECT 2.000 475.520 5.420 476.720 ;
  RECT 4.280 474.740 5.140 475.020 ;
  RECT 2.000 476.720 5.420 477.920 ;
  RECT 2.000 479.200 5.420 480.400 ;
  RECT 4.280 478.420 5.140 478.700 ;
  RECT 2.000 480.400 5.420 481.600 ;
  RECT 2.000 482.880 5.420 484.080 ;
  RECT 4.280 482.100 5.140 482.380 ;
  RECT 2.000 484.080 5.420 485.280 ;
  RECT 2.000 486.560 5.420 487.760 ;
  RECT 4.280 485.780 5.140 486.060 ;
  RECT 2.000 487.760 5.420 488.960 ;
  RECT 2.000 490.240 5.420 491.440 ;
  RECT 4.280 489.460 5.140 489.740 ;
  RECT 2.000 491.440 5.420 492.640 ;
  RECT 2.000 493.920 5.420 495.120 ;
  RECT 4.280 493.140 5.140 493.420 ;
  RECT 2.000 495.120 5.420 496.320 ;
  RECT 2.000 497.600 5.420 498.800 ;
  RECT 4.280 496.820 5.140 497.100 ;
  RECT 2.000 498.800 5.420 500.000 ;
  RECT 2.000 501.280 5.420 502.480 ;
  RECT 4.280 500.500 5.140 500.780 ;
  RECT 2.000 502.480 5.420 503.680 ;
  RECT 2.000 504.960 5.420 506.160 ;
  RECT 4.280 504.180 5.140 504.460 ;
  RECT 2.000 506.160 5.420 507.360 ;
  RECT 2.000 508.640 5.420 509.840 ;
  RECT 4.280 507.860 5.140 508.140 ;
  RECT 2.000 509.840 5.420 511.040 ;
  RECT 2.000 512.320 5.420 513.520 ;
  RECT 4.280 511.540 5.140 511.820 ;
  RECT 2.000 513.520 5.420 514.720 ;
  RECT 2.000 516.000 5.420 517.200 ;
  RECT 4.280 515.220 5.140 515.500 ;
  RECT 2.000 517.200 5.420 518.400 ;
  RECT 2.000 519.680 5.420 520.880 ;
  RECT 4.280 518.900 5.140 519.180 ;
  RECT 2.000 520.880 5.420 522.080 ;
  RECT 2.000 523.360 5.420 524.560 ;
  RECT 4.280 522.580 5.140 522.860 ;
  RECT 2.000 524.560 5.420 525.760 ;
  RECT 2.000 527.040 5.420 528.240 ;
  RECT 4.280 526.260 5.140 526.540 ;
  RECT 2.000 528.240 5.420 529.440 ;
  RECT 2.000 530.720 5.420 531.920 ;
  RECT 4.280 529.940 5.140 530.220 ;
  RECT 2.000 531.920 5.420 533.120 ;
  RECT 2.000 534.400 5.420 535.600 ;
  RECT 4.280 533.620 5.140 533.900 ;
  RECT 2.000 535.600 5.420 536.800 ;
  RECT 2.000 538.080 5.420 539.280 ;
  RECT 4.280 537.300 5.140 537.580 ;
  RECT 2.000 539.280 5.420 540.480 ;
  RECT 2.000 541.760 5.420 542.960 ;
  RECT 4.280 540.980 5.140 541.260 ;
  RECT 2.000 542.960 5.420 544.160 ;
  RECT 2.000 545.440 5.420 546.640 ;
  RECT 4.280 544.660 5.140 544.940 ;
  RECT 2.000 546.640 5.420 547.840 ;
  RECT 2.000 549.120 5.420 550.320 ;
  RECT 4.280 548.340 5.140 548.620 ;
  RECT 2.000 550.320 5.420 551.520 ;
  RECT 2.000 552.800 5.420 554.000 ;
  RECT 4.280 552.020 5.140 552.300 ;
  RECT 4.280 559.940 5.140 560.320 ;
  RECT 47.920 560.510 48.170 563.930 ;
  RECT 47.350 560.790 47.600 561.650 ;
  RECT 88.840 560.510 89.090 563.930 ;
  RECT 88.270 560.790 88.520 561.650 ;
  RECT 129.760 560.510 130.010 563.930 ;
  RECT 129.190 560.790 129.440 561.650 ;
  RECT 170.680 560.510 170.930 563.930 ;
  RECT 170.110 560.790 170.360 561.650 ;
  RECT 211.600 560.510 211.850 563.930 ;
  RECT 211.030 560.790 211.280 561.650 ;
  RECT 252.520 560.510 252.770 563.930 ;
  RECT 251.950 560.790 252.200 561.650 ;
  RECT 293.440 560.510 293.690 563.930 ;
  RECT 292.870 560.790 293.120 561.650 ;
  RECT 334.360 560.510 334.610 563.930 ;
  RECT 333.790 560.790 334.040 561.650 ;
  RECT 375.280 560.510 375.530 563.930 ;
  RECT 374.710 560.790 374.960 561.650 ;
  RECT 416.200 560.510 416.450 563.930 ;
  RECT 415.630 560.790 415.880 561.650 ;
  RECT 457.120 560.510 457.370 563.930 ;
  RECT 456.550 560.790 456.800 561.650 ;
  RECT 498.040 560.510 498.290 563.930 ;
  RECT 497.470 560.790 497.720 561.650 ;
  RECT 538.960 560.510 539.210 563.930 ;
  RECT 538.390 560.790 538.640 561.650 ;
  RECT 579.880 560.510 580.130 563.930 ;
  RECT 579.310 560.790 579.560 561.650 ;
  RECT 620.800 560.510 621.050 563.930 ;
  RECT 620.230 560.790 620.480 561.650 ;
  RECT 661.720 560.510 661.970 563.930 ;
  RECT 661.150 560.790 661.400 561.650 ;
  RECT 702.640 560.510 702.890 563.930 ;
  RECT 702.070 560.790 702.320 561.650 ;
  RECT 743.560 560.510 743.810 563.930 ;
  RECT 742.990 560.790 743.240 561.650 ;
  RECT 784.480 560.510 784.730 563.930 ;
  RECT 783.910 560.790 784.160 561.650 ;
  RECT 825.400 560.510 825.650 563.930 ;
  RECT 824.830 560.790 825.080 561.650 ;
  RECT 866.320 560.510 866.570 563.930 ;
  RECT 865.750 560.790 866.000 561.650 ;
  RECT 907.240 560.510 907.490 563.930 ;
  RECT 906.670 560.790 906.920 561.650 ;
  RECT 948.160 560.510 948.410 563.930 ;
  RECT 947.590 560.790 947.840 561.650 ;
  RECT 989.080 560.510 989.330 563.930 ;
  RECT 988.510 560.790 988.760 561.650 ;
  RECT 1030.000 560.510 1030.250 563.930 ;
  RECT 1029.430 560.790 1029.680 561.650 ;
  RECT 1070.920 560.510 1071.170 563.930 ;
  RECT 1070.350 560.790 1070.600 561.650 ;
  RECT 1111.840 560.510 1112.090 563.930 ;
  RECT 1111.270 560.790 1111.520 561.650 ;
  RECT 1152.760 560.510 1153.010 563.930 ;
  RECT 1152.190 560.790 1152.440 561.650 ;
  RECT 1193.680 560.510 1193.930 563.930 ;
  RECT 1193.110 560.790 1193.360 561.650 ;
  RECT 1234.600 560.510 1234.850 563.930 ;
  RECT 1234.030 560.790 1234.280 561.650 ;
  RECT 1275.520 560.510 1275.770 563.930 ;
  RECT 1274.950 560.790 1275.200 561.650 ;
  RECT 0.000 563.930 2692.940 565.930 ;
  RECT 0.000 1.600 2692.940 3.600 ;
  RECT 2690.940 1.600 2692.940 565.930 ;
  RECT 0.000 1.600 2.000 565.930 ;
  LAYER ME2 ;
  RECT 5.420 7.020 2687.520 560.510 ;
  RECT 2691.080 3.460 2692.940 564.070 ;
  RECT 0.000 3.460 1.860 564.070 ;
  RECT 1.860 564.070 2691.080 565.930 ;
  RECT 2682.600 1.600 2691.080 3.460 ;
  RECT 2668.200 1.600 2680.280 3.460 ;
  RECT 2663.000 1.600 2665.650 3.460 ;
  RECT 2648.200 1.600 2660.440 3.460 ;
  RECT 2641.800 1.600 2645.810 3.460 ;
  RECT 2627.400 1.600 2639.360 3.460 ;
  RECT 2622.200 1.600 2624.730 3.460 ;
  RECT 2607.400 1.600 2619.520 3.460 ;
  RECT 2601.000 1.600 2604.890 3.460 ;
  RECT 2586.200 1.600 2598.440 3.460 ;
  RECT 2581.000 1.600 2583.810 3.460 ;
  RECT 2566.600 1.600 2578.600 3.460 ;
  RECT 2560.200 1.600 2563.970 3.460 ;
  RECT 2545.400 1.600 2557.520 3.460 ;
  RECT 2540.200 1.600 2542.890 3.460 ;
  RECT 2527.400 1.600 2537.680 3.460 ;
  RECT 2519.000 1.600 2523.050 3.460 ;
  RECT 2504.600 1.600 2516.600 3.460 ;
  RECT 2499.400 1.600 2501.970 3.460 ;
  RECT 2484.600 1.600 2496.760 3.460 ;
  RECT 2478.200 1.600 2482.130 3.460 ;
  RECT 2463.400 1.600 2475.680 3.460 ;
  RECT 2458.200 1.600 2461.050 3.460 ;
  RECT 2443.800 1.600 2455.840 3.460 ;
  RECT 2437.400 1.600 2441.210 3.460 ;
  RECT 2422.600 1.600 2434.760 3.460 ;
  RECT 2417.400 1.600 2420.130 3.460 ;
  RECT 2402.600 1.600 2414.920 3.460 ;
  RECT 2396.200 1.600 2400.290 3.460 ;
  RECT 2381.800 1.600 2393.840 3.460 ;
  RECT 2376.600 1.600 2379.210 3.460 ;
  RECT 2363.400 1.600 2374.000 3.460 ;
  RECT 2355.400 1.600 2359.370 3.460 ;
  RECT 2340.600 1.600 2352.920 3.460 ;
  RECT 2335.400 1.600 2338.290 3.460 ;
  RECT 2321.000 1.600 2333.080 3.460 ;
  RECT 2314.600 1.600 2318.450 3.460 ;
  RECT 2299.800 1.600 2312.000 3.460 ;
  RECT 2294.600 1.600 2297.370 3.460 ;
  RECT 2280.200 1.600 2292.160 3.460 ;
  RECT 2273.400 1.600 2277.530 3.460 ;
  RECT 2259.000 1.600 2271.080 3.460 ;
  RECT 2253.800 1.600 2256.450 3.460 ;
  RECT 2239.000 1.600 2251.240 3.460 ;
  RECT 2232.600 1.600 2236.610 3.460 ;
  RECT 2218.200 1.600 2230.160 3.460 ;
  RECT 2213.000 1.600 2215.530 3.460 ;
  RECT 2199.800 1.600 2210.320 3.460 ;
  RECT 2191.800 1.600 2195.690 3.460 ;
  RECT 2177.000 1.600 2189.240 3.460 ;
  RECT 2171.800 1.600 2174.610 3.460 ;
  RECT 2157.400 1.600 2169.400 3.460 ;
  RECT 2151.000 1.600 2154.770 3.460 ;
  RECT 2136.200 1.600 2148.320 3.460 ;
  RECT 2131.000 1.600 2133.690 3.460 ;
  RECT 2116.200 1.600 2128.480 3.460 ;
  RECT 2109.800 1.600 2113.850 3.460 ;
  RECT 2095.400 1.600 2107.400 3.460 ;
  RECT 2090.200 1.600 2092.770 3.460 ;
  RECT 2075.400 1.600 2087.560 3.460 ;
  RECT 2069.000 1.600 2072.930 3.460 ;
  RECT 2054.200 1.600 2066.480 3.460 ;
  RECT 2049.000 1.600 2051.850 3.460 ;
  RECT 2036.200 1.600 2046.640 3.460 ;
  RECT 2028.200 1.600 2032.010 3.460 ;
  RECT 2013.400 1.600 2025.560 3.460 ;
  RECT 2008.200 1.600 2010.930 3.460 ;
  RECT 1993.400 1.600 2005.720 3.460 ;
  RECT 1987.000 1.600 1991.090 3.460 ;
  RECT 1972.600 1.600 1984.640 3.460 ;
  RECT 1967.400 1.600 1970.010 3.460 ;
  RECT 1952.600 1.600 1964.800 3.460 ;
  RECT 1946.200 1.600 1950.170 3.460 ;
  RECT 1931.400 1.600 1943.720 3.460 ;
  RECT 1926.200 1.600 1929.090 3.460 ;
  RECT 1911.800 1.600 1923.880 3.460 ;
  RECT 1905.400 1.600 1909.250 3.460 ;
  RECT 1890.600 1.600 1902.800 3.460 ;
  RECT 1885.400 1.600 1888.170 3.460 ;
  RECT 1872.600 1.600 1882.960 3.460 ;
  RECT 1864.200 1.600 1868.330 3.460 ;
  RECT 1849.800 1.600 1861.880 3.460 ;
  RECT 1844.600 1.600 1847.250 3.460 ;
  RECT 1829.800 1.600 1842.040 3.460 ;
  RECT 1823.400 1.600 1827.410 3.460 ;
  RECT 1809.000 1.600 1820.960 3.460 ;
  RECT 1803.800 1.600 1806.330 3.460 ;
  RECT 1789.000 1.600 1801.120 3.460 ;
  RECT 1782.600 1.600 1786.490 3.460 ;
  RECT 1767.800 1.600 1780.040 3.460 ;
  RECT 1762.600 1.600 1765.410 3.460 ;
  RECT 1748.200 1.600 1760.200 3.460 ;
  RECT 1741.800 1.600 1745.570 3.460 ;
  RECT 1727.000 1.600 1739.120 3.460 ;
  RECT 1721.800 1.600 1724.490 3.460 ;
  RECT 1709.000 1.600 1719.280 3.460 ;
  RECT 1700.600 1.600 1704.650 3.460 ;
  RECT 1686.200 1.600 1698.200 3.460 ;
  RECT 1681.000 1.600 1683.570 3.460 ;
  RECT 1666.200 1.600 1678.360 3.460 ;
  RECT 1659.800 1.600 1663.730 3.460 ;
  RECT 1645.000 1.600 1657.280 3.460 ;
  RECT 1639.800 1.600 1642.650 3.460 ;
  RECT 1625.400 1.600 1637.440 3.460 ;
  RECT 1619.000 1.600 1622.810 3.460 ;
  RECT 1604.200 1.600 1616.360 3.460 ;
  RECT 1599.000 1.600 1601.730 3.460 ;
  RECT 1584.200 1.600 1596.520 3.460 ;
  RECT 1577.800 1.600 1581.890 3.460 ;
  RECT 1563.400 1.600 1575.440 3.460 ;
  RECT 1558.200 1.600 1560.810 3.460 ;
  RECT 1545.000 1.600 1555.600 3.460 ;
  RECT 1537.000 1.600 1540.970 3.460 ;
  RECT 1522.200 1.600 1534.520 3.460 ;
  RECT 1517.000 1.600 1519.890 3.460 ;
  RECT 1502.600 1.600 1514.680 3.460 ;
  RECT 1496.200 1.600 1500.050 3.460 ;
  RECT 1481.400 1.600 1493.600 3.460 ;
  RECT 1476.200 1.600 1478.970 3.460 ;
  RECT 1461.800 1.600 1473.760 3.460 ;
  RECT 1455.000 1.600 1459.130 3.460 ;
  RECT 1440.600 1.600 1452.680 3.460 ;
  RECT 1435.400 1.600 1438.050 3.460 ;
  RECT 1420.600 1.600 1432.840 3.460 ;
  RECT 1414.200 1.600 1418.210 3.460 ;
  RECT 1399.800 1.600 1411.760 3.460 ;
  RECT 1394.600 1.600 1397.130 3.460 ;
  RECT 1381.400 1.600 1391.920 3.460 ;
  RECT 1359.000 1.600 1377.290 3.460 ;
  RECT 1347.000 1.600 1350.450 3.460 ;
  RECT 1339.800 1.600 1344.480 3.460 ;
  RECT 1313.000 1.600 1319.840 3.460 ;
  RECT 1298.200 1.600 1310.460 3.460 ;
  RECT 1293.000 1.600 1295.830 3.460 ;
  RECT 1278.600 1.600 1290.620 3.460 ;
  RECT 1272.200 1.600 1275.990 3.460 ;
  RECT 1257.400 1.600 1269.540 3.460 ;
  RECT 1252.200 1.600 1254.910 3.460 ;
  RECT 1237.400 1.600 1249.700 3.460 ;
  RECT 1231.000 1.600 1235.070 3.460 ;
  RECT 1216.600 1.600 1228.620 3.460 ;
  RECT 1211.400 1.600 1213.990 3.460 ;
  RECT 1196.600 1.600 1208.780 3.460 ;
  RECT 1190.200 1.600 1194.150 3.460 ;
  RECT 1175.400 1.600 1187.700 3.460 ;
  RECT 1170.200 1.600 1173.070 3.460 ;
  RECT 1157.400 1.600 1167.860 3.460 ;
  RECT 1149.400 1.600 1153.230 3.460 ;
  RECT 1134.600 1.600 1146.780 3.460 ;
  RECT 1129.400 1.600 1132.150 3.460 ;
  RECT 1115.000 1.600 1126.940 3.460 ;
  RECT 1108.200 1.600 1112.310 3.460 ;
  RECT 1093.800 1.600 1105.860 3.460 ;
  RECT 1088.600 1.600 1091.230 3.460 ;
  RECT 1073.800 1.600 1086.020 3.460 ;
  RECT 1067.400 1.600 1071.390 3.460 ;
  RECT 1053.000 1.600 1064.940 3.460 ;
  RECT 1047.400 1.600 1050.310 3.460 ;
  RECT 1033.000 1.600 1045.100 3.460 ;
  RECT 1026.600 1.600 1030.470 3.460 ;
  RECT 1011.800 1.600 1024.020 3.460 ;
  RECT 1006.600 1.600 1009.390 3.460 ;
  RECT 993.800 1.600 1004.180 3.460 ;
  RECT 985.400 1.600 989.550 3.460 ;
  RECT 971.000 1.600 983.100 3.460 ;
  RECT 965.800 1.600 968.470 3.460 ;
  RECT 951.000 1.600 963.260 3.460 ;
  RECT 944.600 1.600 948.630 3.460 ;
  RECT 930.200 1.600 942.180 3.460 ;
  RECT 925.000 1.600 927.550 3.460 ;
  RECT 910.200 1.600 922.340 3.460 ;
  RECT 903.800 1.600 907.710 3.460 ;
  RECT 889.000 1.600 901.260 3.460 ;
  RECT 883.800 1.600 886.630 3.460 ;
  RECT 869.400 1.600 881.420 3.460 ;
  RECT 863.000 1.600 866.790 3.460 ;
  RECT 848.200 1.600 860.340 3.460 ;
  RECT 843.000 1.600 845.710 3.460 ;
  RECT 830.200 1.600 840.500 3.460 ;
  RECT 821.800 1.600 825.870 3.460 ;
  RECT 807.400 1.600 819.420 3.460 ;
  RECT 802.200 1.600 804.790 3.460 ;
  RECT 787.400 1.600 799.580 3.460 ;
  RECT 781.000 1.600 784.950 3.460 ;
  RECT 766.200 1.600 778.500 3.460 ;
  RECT 761.000 1.600 763.870 3.460 ;
  RECT 746.600 1.600 758.660 3.460 ;
  RECT 740.200 1.600 744.030 3.460 ;
  RECT 725.400 1.600 737.580 3.460 ;
  RECT 720.200 1.600 722.950 3.460 ;
  RECT 705.800 1.600 717.740 3.460 ;
  RECT 699.000 1.600 703.110 3.460 ;
  RECT 684.600 1.600 696.660 3.460 ;
  RECT 679.400 1.600 682.030 3.460 ;
  RECT 666.600 1.600 676.820 3.460 ;
  RECT 658.200 1.600 662.190 3.460 ;
  RECT 643.800 1.600 655.740 3.460 ;
  RECT 638.200 1.600 641.110 3.460 ;
  RECT 623.800 1.600 635.900 3.460 ;
  RECT 617.400 1.600 621.270 3.460 ;
  RECT 602.600 1.600 614.820 3.460 ;
  RECT 597.400 1.600 600.190 3.460 ;
  RECT 583.000 1.600 594.980 3.460 ;
  RECT 576.200 1.600 580.350 3.460 ;
  RECT 561.800 1.600 573.900 3.460 ;
  RECT 556.600 1.600 559.270 3.460 ;
  RECT 541.800 1.600 554.060 3.460 ;
  RECT 535.400 1.600 539.430 3.460 ;
  RECT 521.000 1.600 532.980 3.460 ;
  RECT 515.800 1.600 518.350 3.460 ;
  RECT 502.600 1.600 513.140 3.460 ;
  RECT 494.600 1.600 498.510 3.460 ;
  RECT 479.800 1.600 492.060 3.460 ;
  RECT 474.600 1.600 477.430 3.460 ;
  RECT 460.200 1.600 472.220 3.460 ;
  RECT 453.800 1.600 457.590 3.460 ;
  RECT 439.000 1.600 451.140 3.460 ;
  RECT 433.800 1.600 436.510 3.460 ;
  RECT 419.000 1.600 431.300 3.460 ;
  RECT 412.600 1.600 416.670 3.460 ;
  RECT 398.200 1.600 410.220 3.460 ;
  RECT 393.000 1.600 395.590 3.460 ;
  RECT 378.200 1.600 390.380 3.460 ;
  RECT 371.800 1.600 375.750 3.460 ;
  RECT 357.000 1.600 369.300 3.460 ;
  RECT 351.800 1.600 354.670 3.460 ;
  RECT 339.000 1.600 349.460 3.460 ;
  RECT 331.000 1.600 334.830 3.460 ;
  RECT 316.200 1.600 328.380 3.460 ;
  RECT 311.000 1.600 313.750 3.460 ;
  RECT 296.600 1.600 308.540 3.460 ;
  RECT 289.800 1.600 293.910 3.460 ;
  RECT 275.400 1.600 287.460 3.460 ;
  RECT 270.200 1.600 272.830 3.460 ;
  RECT 255.400 1.600 267.620 3.460 ;
  RECT 249.000 1.600 252.990 3.460 ;
  RECT 234.600 1.600 246.540 3.460 ;
  RECT 229.000 1.600 231.910 3.460 ;
  RECT 214.600 1.600 226.700 3.460 ;
  RECT 208.200 1.600 212.070 3.460 ;
  RECT 193.400 1.600 205.620 3.460 ;
  RECT 188.200 1.600 190.990 3.460 ;
  RECT 175.400 1.600 185.780 3.460 ;
  RECT 167.000 1.600 171.150 3.460 ;
  RECT 152.600 1.600 164.700 3.460 ;
  RECT 147.400 1.600 150.070 3.460 ;
  RECT 132.600 1.600 144.860 3.460 ;
  RECT 126.200 1.600 130.230 3.460 ;
  RECT 111.800 1.600 123.780 3.460 ;
  RECT 106.600 1.600 109.150 3.460 ;
  RECT 91.800 1.600 103.940 3.460 ;
  RECT 85.400 1.600 89.310 3.460 ;
  RECT 70.600 1.600 82.860 3.460 ;
  RECT 65.400 1.600 68.230 3.460 ;
  RECT 51.000 1.600 63.020 3.460 ;
  RECT 44.600 1.600 48.390 3.460 ;
  RECT 29.800 1.600 41.940 3.460 ;
  RECT 24.600 1.600 27.310 3.460 ;
  RECT 11.800 1.600 22.100 3.460 ;
  RECT 1.860 1.600 7.470 3.460 ;
  RECT 2688.940 5.600 2690.800 561.930 ;
  RECT 2.140 5.600 4.000 561.930 ;
  RECT 4.000 561.930 2688.940 563.790 ;
  RECT 2682.600 3.740 2688.940 5.600 ;
  RECT 2668.200 3.740 2680.280 5.600 ;
  RECT 2663.000 3.740 2665.650 5.600 ;
  RECT 2648.200 3.740 2660.440 5.600 ;
  RECT 2641.800 3.740 2645.810 5.600 ;
  RECT 2627.400 3.740 2639.360 5.600 ;
  RECT 2622.200 3.740 2624.730 5.600 ;
  RECT 2607.400 3.740 2619.520 5.600 ;
  RECT 2601.000 3.740 2604.890 5.600 ;
  RECT 2586.200 3.740 2598.440 5.600 ;
  RECT 2581.000 3.740 2583.810 5.600 ;
  RECT 2566.600 3.740 2578.600 5.600 ;
  RECT 2560.200 3.740 2563.970 5.600 ;
  RECT 2545.400 3.740 2557.520 5.600 ;
  RECT 2540.200 3.740 2542.890 5.600 ;
  RECT 2527.400 3.740 2537.680 5.600 ;
  RECT 2519.000 3.740 2523.050 5.600 ;
  RECT 2504.600 3.740 2516.600 5.600 ;
  RECT 2499.400 3.740 2501.970 5.600 ;
  RECT 2484.600 3.740 2496.760 5.600 ;
  RECT 2478.200 3.740 2482.130 5.600 ;
  RECT 2463.400 3.740 2475.680 5.600 ;
  RECT 2458.200 3.740 2461.050 5.600 ;
  RECT 2443.800 3.740 2455.840 5.600 ;
  RECT 2437.400 3.740 2441.210 5.600 ;
  RECT 2422.600 3.740 2434.760 5.600 ;
  RECT 2417.400 3.740 2420.130 5.600 ;
  RECT 2402.600 3.740 2414.920 5.600 ;
  RECT 2396.200 3.740 2400.290 5.600 ;
  RECT 2381.800 3.740 2393.840 5.600 ;
  RECT 2376.600 3.740 2379.210 5.600 ;
  RECT 2363.400 3.740 2374.000 5.600 ;
  RECT 2355.400 3.740 2359.370 5.600 ;
  RECT 2340.600 3.740 2352.920 5.600 ;
  RECT 2335.400 3.740 2338.290 5.600 ;
  RECT 2321.000 3.740 2333.080 5.600 ;
  RECT 2314.600 3.740 2318.450 5.600 ;
  RECT 2299.800 3.740 2312.000 5.600 ;
  RECT 2294.600 3.740 2297.370 5.600 ;
  RECT 2280.200 3.740 2292.160 5.600 ;
  RECT 2273.400 3.740 2277.530 5.600 ;
  RECT 2259.000 3.740 2271.080 5.600 ;
  RECT 2253.800 3.740 2256.450 5.600 ;
  RECT 2239.000 3.740 2251.240 5.600 ;
  RECT 2232.600 3.740 2236.610 5.600 ;
  RECT 2218.200 3.740 2230.160 5.600 ;
  RECT 2213.000 3.740 2215.530 5.600 ;
  RECT 2199.800 3.740 2210.320 5.600 ;
  RECT 2191.800 3.740 2195.690 5.600 ;
  RECT 2177.000 3.740 2189.240 5.600 ;
  RECT 2171.800 3.740 2174.610 5.600 ;
  RECT 2157.400 3.740 2169.400 5.600 ;
  RECT 2151.000 3.740 2154.770 5.600 ;
  RECT 2136.200 3.740 2148.320 5.600 ;
  RECT 2131.000 3.740 2133.690 5.600 ;
  RECT 2116.200 3.740 2128.480 5.600 ;
  RECT 2109.800 3.740 2113.850 5.600 ;
  RECT 2095.400 3.740 2107.400 5.600 ;
  RECT 2090.200 3.740 2092.770 5.600 ;
  RECT 2075.400 3.740 2087.560 5.600 ;
  RECT 2069.000 3.740 2072.930 5.600 ;
  RECT 2054.200 3.740 2066.480 5.600 ;
  RECT 2049.000 3.740 2051.850 5.600 ;
  RECT 2036.200 3.740 2046.640 5.600 ;
  RECT 2028.200 3.740 2032.010 5.600 ;
  RECT 2013.400 3.740 2025.560 5.600 ;
  RECT 2008.200 3.740 2010.930 5.600 ;
  RECT 1993.400 3.740 2005.720 5.600 ;
  RECT 1987.000 3.740 1991.090 5.600 ;
  RECT 1972.600 3.740 1984.640 5.600 ;
  RECT 1967.400 3.740 1970.010 5.600 ;
  RECT 1952.600 3.740 1964.800 5.600 ;
  RECT 1946.200 3.740 1950.170 5.600 ;
  RECT 1931.400 3.740 1943.720 5.600 ;
  RECT 1926.200 3.740 1929.090 5.600 ;
  RECT 1911.800 3.740 1923.880 5.600 ;
  RECT 1905.400 3.740 1909.250 5.600 ;
  RECT 1890.600 3.740 1902.800 5.600 ;
  RECT 1885.400 3.740 1888.170 5.600 ;
  RECT 1872.600 3.740 1882.960 5.600 ;
  RECT 1864.200 3.740 1868.330 5.600 ;
  RECT 1849.800 3.740 1861.880 5.600 ;
  RECT 1844.600 3.740 1847.250 5.600 ;
  RECT 1829.800 3.740 1842.040 5.600 ;
  RECT 1823.400 3.740 1827.410 5.600 ;
  RECT 1809.000 3.740 1820.960 5.600 ;
  RECT 1803.800 3.740 1806.330 5.600 ;
  RECT 1789.000 3.740 1801.120 5.600 ;
  RECT 1782.600 3.740 1786.490 5.600 ;
  RECT 1767.800 3.740 1780.040 5.600 ;
  RECT 1762.600 3.740 1765.410 5.600 ;
  RECT 1748.200 3.740 1760.200 5.600 ;
  RECT 1741.800 3.740 1745.570 5.600 ;
  RECT 1727.000 3.740 1739.120 5.600 ;
  RECT 1721.800 3.740 1724.490 5.600 ;
  RECT 1709.000 3.740 1719.280 5.600 ;
  RECT 1700.600 3.740 1704.650 5.600 ;
  RECT 1686.200 3.740 1698.200 5.600 ;
  RECT 1681.000 3.740 1683.570 5.600 ;
  RECT 1666.200 3.740 1678.360 5.600 ;
  RECT 1659.800 3.740 1663.730 5.600 ;
  RECT 1645.000 3.740 1657.280 5.600 ;
  RECT 1639.800 3.740 1642.650 5.600 ;
  RECT 1625.400 3.740 1637.440 5.600 ;
  RECT 1619.000 3.740 1622.810 5.600 ;
  RECT 1604.200 3.740 1616.360 5.600 ;
  RECT 1599.000 3.740 1601.730 5.600 ;
  RECT 1584.200 3.740 1596.520 5.600 ;
  RECT 1577.800 3.740 1581.890 5.600 ;
  RECT 1563.400 3.740 1575.440 5.600 ;
  RECT 1558.200 3.740 1560.810 5.600 ;
  RECT 1545.000 3.740 1555.600 5.600 ;
  RECT 1537.000 3.740 1540.970 5.600 ;
  RECT 1522.200 3.740 1534.520 5.600 ;
  RECT 1517.000 3.740 1519.890 5.600 ;
  RECT 1502.600 3.740 1514.680 5.600 ;
  RECT 1496.200 3.740 1500.050 5.600 ;
  RECT 1481.400 3.740 1493.600 5.600 ;
  RECT 1476.200 3.740 1478.970 5.600 ;
  RECT 1461.800 3.740 1473.760 5.600 ;
  RECT 1455.000 3.740 1459.130 5.600 ;
  RECT 1440.600 3.740 1452.680 5.600 ;
  RECT 1435.400 3.740 1438.050 5.600 ;
  RECT 1420.600 3.740 1432.840 5.600 ;
  RECT 1414.200 3.740 1418.210 5.600 ;
  RECT 1399.800 3.740 1411.760 5.600 ;
  RECT 1394.600 3.740 1397.130 5.600 ;
  RECT 1381.400 3.740 1391.920 5.600 ;
  RECT 1359.000 3.740 1377.290 5.600 ;
  RECT 1347.000 3.740 1350.450 5.600 ;
  RECT 1339.800 3.740 1344.480 5.600 ;
  RECT 1313.000 3.740 1319.840 5.600 ;
  RECT 1298.200 3.740 1310.460 5.600 ;
  RECT 1293.000 3.740 1295.830 5.600 ;
  RECT 1278.600 3.740 1290.620 5.600 ;
  RECT 1272.200 3.740 1275.990 5.600 ;
  RECT 1257.400 3.740 1269.540 5.600 ;
  RECT 1252.200 3.740 1254.910 5.600 ;
  RECT 1237.400 3.740 1249.700 5.600 ;
  RECT 1231.000 3.740 1235.070 5.600 ;
  RECT 1216.600 3.740 1228.620 5.600 ;
  RECT 1211.400 3.740 1213.990 5.600 ;
  RECT 1196.600 3.740 1208.780 5.600 ;
  RECT 1190.200 3.740 1194.150 5.600 ;
  RECT 1175.400 3.740 1187.700 5.600 ;
  RECT 1170.200 3.740 1173.070 5.600 ;
  RECT 1157.400 3.740 1167.860 5.600 ;
  RECT 1149.400 3.740 1153.230 5.600 ;
  RECT 1134.600 3.740 1146.780 5.600 ;
  RECT 1129.400 3.740 1132.150 5.600 ;
  RECT 1115.000 3.740 1126.940 5.600 ;
  RECT 1108.200 3.740 1112.310 5.600 ;
  RECT 1093.800 3.740 1105.860 5.600 ;
  RECT 1088.600 3.740 1091.230 5.600 ;
  RECT 1073.800 3.740 1086.020 5.600 ;
  RECT 1067.400 3.740 1071.390 5.600 ;
  RECT 1053.000 3.740 1064.940 5.600 ;
  RECT 1047.400 3.740 1050.310 5.600 ;
  RECT 1033.000 3.740 1045.100 5.600 ;
  RECT 1026.600 3.740 1030.470 5.600 ;
  RECT 1011.800 3.740 1024.020 5.600 ;
  RECT 1006.600 3.740 1009.390 5.600 ;
  RECT 993.800 3.740 1004.180 5.600 ;
  RECT 985.400 3.740 989.550 5.600 ;
  RECT 971.000 3.740 983.100 5.600 ;
  RECT 965.800 3.740 968.470 5.600 ;
  RECT 951.000 3.740 963.260 5.600 ;
  RECT 944.600 3.740 948.630 5.600 ;
  RECT 930.200 3.740 942.180 5.600 ;
  RECT 925.000 3.740 927.550 5.600 ;
  RECT 910.200 3.740 922.340 5.600 ;
  RECT 903.800 3.740 907.710 5.600 ;
  RECT 889.000 3.740 901.260 5.600 ;
  RECT 883.800 3.740 886.630 5.600 ;
  RECT 869.400 3.740 881.420 5.600 ;
  RECT 863.000 3.740 866.790 5.600 ;
  RECT 848.200 3.740 860.340 5.600 ;
  RECT 843.000 3.740 845.710 5.600 ;
  RECT 830.200 3.740 840.500 5.600 ;
  RECT 821.800 3.740 825.870 5.600 ;
  RECT 807.400 3.740 819.420 5.600 ;
  RECT 802.200 3.740 804.790 5.600 ;
  RECT 787.400 3.740 799.580 5.600 ;
  RECT 781.000 3.740 784.950 5.600 ;
  RECT 766.200 3.740 778.500 5.600 ;
  RECT 761.000 3.740 763.870 5.600 ;
  RECT 746.600 3.740 758.660 5.600 ;
  RECT 740.200 3.740 744.030 5.600 ;
  RECT 725.400 3.740 737.580 5.600 ;
  RECT 720.200 3.740 722.950 5.600 ;
  RECT 705.800 3.740 717.740 5.600 ;
  RECT 699.000 3.740 703.110 5.600 ;
  RECT 684.600 3.740 696.660 5.600 ;
  RECT 679.400 3.740 682.030 5.600 ;
  RECT 666.600 3.740 676.820 5.600 ;
  RECT 658.200 3.740 662.190 5.600 ;
  RECT 643.800 3.740 655.740 5.600 ;
  RECT 638.200 3.740 641.110 5.600 ;
  RECT 623.800 3.740 635.900 5.600 ;
  RECT 617.400 3.740 621.270 5.600 ;
  RECT 602.600 3.740 614.820 5.600 ;
  RECT 597.400 3.740 600.190 5.600 ;
  RECT 583.000 3.740 594.980 5.600 ;
  RECT 576.200 3.740 580.350 5.600 ;
  RECT 561.800 3.740 573.900 5.600 ;
  RECT 556.600 3.740 559.270 5.600 ;
  RECT 541.800 3.740 554.060 5.600 ;
  RECT 535.400 3.740 539.430 5.600 ;
  RECT 521.000 3.740 532.980 5.600 ;
  RECT 515.800 3.740 518.350 5.600 ;
  RECT 502.600 3.740 513.140 5.600 ;
  RECT 494.600 3.740 498.510 5.600 ;
  RECT 479.800 3.740 492.060 5.600 ;
  RECT 474.600 3.740 477.430 5.600 ;
  RECT 460.200 3.740 472.220 5.600 ;
  RECT 453.800 3.740 457.590 5.600 ;
  RECT 439.000 3.740 451.140 5.600 ;
  RECT 433.800 3.740 436.510 5.600 ;
  RECT 419.000 3.740 431.300 5.600 ;
  RECT 412.600 3.740 416.670 5.600 ;
  RECT 398.200 3.740 410.220 5.600 ;
  RECT 393.000 3.740 395.590 5.600 ;
  RECT 378.200 3.740 390.380 5.600 ;
  RECT 371.800 3.740 375.750 5.600 ;
  RECT 357.000 3.740 369.300 5.600 ;
  RECT 351.800 3.740 354.670 5.600 ;
  RECT 339.000 3.740 349.460 5.600 ;
  RECT 331.000 3.740 334.830 5.600 ;
  RECT 316.200 3.740 328.380 5.600 ;
  RECT 311.000 3.740 313.750 5.600 ;
  RECT 296.600 3.740 308.540 5.600 ;
  RECT 289.800 3.740 293.910 5.600 ;
  RECT 275.400 3.740 287.460 5.600 ;
  RECT 270.200 3.740 272.830 5.600 ;
  RECT 255.400 3.740 267.620 5.600 ;
  RECT 249.000 3.740 252.990 5.600 ;
  RECT 234.600 3.740 246.540 5.600 ;
  RECT 229.000 3.740 231.910 5.600 ;
  RECT 214.600 3.740 226.700 5.600 ;
  RECT 208.200 3.740 212.070 5.600 ;
  RECT 193.400 3.740 205.620 5.600 ;
  RECT 188.200 3.740 190.990 5.600 ;
  RECT 175.400 3.740 185.780 5.600 ;
  RECT 167.000 3.740 171.150 5.600 ;
  RECT 152.600 3.740 164.700 5.600 ;
  RECT 147.400 3.740 150.070 5.600 ;
  RECT 132.600 3.740 144.860 5.600 ;
  RECT 126.200 3.740 130.230 5.600 ;
  RECT 111.800 3.740 123.780 5.600 ;
  RECT 106.600 3.740 109.150 5.600 ;
  RECT 91.800 3.740 103.940 5.600 ;
  RECT 85.400 3.740 89.310 5.600 ;
  RECT 70.600 3.740 82.860 5.600 ;
  RECT 65.400 3.740 68.230 5.600 ;
  RECT 51.000 3.740 63.020 5.600 ;
  RECT 44.600 3.740 48.390 5.600 ;
  RECT 29.800 3.740 41.940 5.600 ;
  RECT 24.600 3.740 27.310 5.600 ;
  RECT 11.800 3.740 22.100 5.600 ;
  RECT 4.000 3.740 7.470 5.600 ;
  RECT 2.140 561.930 4.000 563.790 ;
  RECT 0.000 564.070 1.860 565.930 ;
  RECT 2688.940 3.740 2690.800 5.600 ;
  RECT 2691.080 1.600 2692.940 3.460 ;
  RECT 2688.940 561.930 2690.800 563.790 ;
  RECT 2691.080 564.070 2692.940 565.930 ;
  RECT 2.140 3.740 4.000 5.600 ;
  RECT 0.000 1.600 1.860 3.460 ;
  RECT 2680.800 0.000 2681.600 1.000 ;
  RECT 2681.100 1.000 2681.300 5.200 ;
  RECT 2681.100 5.200 2681.480 5.400 ;
  RECT 2681.280 5.400 2681.480 7.020 ;
  RECT 2666.400 0.000 2667.200 1.000 ;
  RECT 2666.700 1.000 2666.900 5.200 ;
  RECT 2666.650 5.200 2666.900 5.400 ;
  RECT 2666.650 5.400 2666.850 7.020 ;
  RECT 2661.200 0.000 2662.000 1.000 ;
  RECT 2661.500 1.000 2661.700 5.200 ;
  RECT 2661.440 5.200 2661.700 5.400 ;
  RECT 2661.440 5.400 2661.640 7.020 ;
  RECT 2646.400 0.000 2647.200 1.000 ;
  RECT 2646.700 1.000 2646.900 5.200 ;
  RECT 2646.700 5.200 2647.010 5.400 ;
  RECT 2646.810 5.400 2647.010 7.020 ;
  RECT 2640.000 0.000 2640.800 1.000 ;
  RECT 2640.300 1.000 2640.500 5.200 ;
  RECT 2640.300 5.200 2640.560 5.400 ;
  RECT 2640.360 5.400 2640.560 7.020 ;
  RECT 2625.600 0.000 2626.400 1.000 ;
  RECT 2625.900 1.000 2626.100 5.200 ;
  RECT 2625.730 5.200 2626.100 5.400 ;
  RECT 2625.730 5.400 2625.930 7.020 ;
  RECT 2620.400 0.000 2621.200 1.000 ;
  RECT 2620.700 1.000 2620.900 5.200 ;
  RECT 2620.520 5.200 2620.900 5.400 ;
  RECT 2620.520 5.400 2620.720 7.020 ;
  RECT 2605.600 0.000 2606.400 1.000 ;
  RECT 2605.900 1.000 2606.100 5.200 ;
  RECT 2605.890 5.200 2606.100 5.400 ;
  RECT 2605.890 5.400 2606.090 7.020 ;
  RECT 2599.200 0.000 2600.000 1.000 ;
  RECT 2599.500 1.000 2599.700 5.200 ;
  RECT 2599.440 5.200 2599.700 5.400 ;
  RECT 2599.440 5.400 2599.640 7.020 ;
  RECT 2584.400 0.000 2585.200 1.000 ;
  RECT 2584.700 1.000 2584.900 5.200 ;
  RECT 2584.700 5.200 2585.010 5.400 ;
  RECT 2584.810 5.400 2585.010 7.020 ;
  RECT 2579.200 0.000 2580.000 1.000 ;
  RECT 2579.500 1.000 2579.700 5.200 ;
  RECT 2579.500 5.200 2579.800 5.400 ;
  RECT 2579.600 5.400 2579.800 7.020 ;
  RECT 2564.800 0.000 2565.600 1.000 ;
  RECT 2565.100 1.000 2565.300 5.200 ;
  RECT 2564.970 5.200 2565.300 5.400 ;
  RECT 2564.970 5.400 2565.170 7.020 ;
  RECT 2558.400 0.000 2559.200 1.000 ;
  RECT 2558.700 1.000 2558.900 5.200 ;
  RECT 2558.520 5.200 2558.900 5.400 ;
  RECT 2558.520 5.400 2558.720 7.020 ;
  RECT 2543.600 0.000 2544.400 1.000 ;
  RECT 2543.900 1.000 2544.100 5.200 ;
  RECT 2543.890 5.200 2544.100 5.400 ;
  RECT 2543.890 5.400 2544.090 7.020 ;
  RECT 2538.400 0.000 2539.200 1.000 ;
  RECT 2538.700 1.000 2538.900 5.200 ;
  RECT 2538.680 5.200 2538.900 5.400 ;
  RECT 2538.680 5.400 2538.880 7.020 ;
  RECT 2525.600 0.000 2526.400 1.000 ;
  RECT 2525.900 1.000 2526.100 5.200 ;
  RECT 2525.770 5.200 2526.100 5.400 ;
  RECT 2525.770 5.400 2525.970 7.020 ;
  RECT 2523.600 0.000 2524.400 1.000 ;
  RECT 2523.900 1.000 2524.100 5.200 ;
  RECT 2523.900 5.200 2524.250 5.400 ;
  RECT 2524.050 5.400 2524.250 7.020 ;
  RECT 2517.200 0.000 2518.000 1.000 ;
  RECT 2517.500 1.000 2517.700 5.200 ;
  RECT 2517.500 5.200 2517.800 5.400 ;
  RECT 2517.600 5.400 2517.800 7.020 ;
  RECT 2502.800 0.000 2503.600 1.000 ;
  RECT 2503.100 1.000 2503.300 5.200 ;
  RECT 2502.970 5.200 2503.300 5.400 ;
  RECT 2502.970 5.400 2503.170 7.020 ;
  RECT 2497.600 0.000 2498.400 1.000 ;
  RECT 2497.900 1.000 2498.100 5.200 ;
  RECT 2497.760 5.200 2498.100 5.400 ;
  RECT 2497.760 5.400 2497.960 7.020 ;
  RECT 2482.800 0.000 2483.600 1.000 ;
  RECT 2483.100 1.000 2483.300 5.200 ;
  RECT 2483.100 5.200 2483.330 5.400 ;
  RECT 2483.130 5.400 2483.330 7.020 ;
  RECT 2476.400 0.000 2477.200 1.000 ;
  RECT 2476.700 1.000 2476.900 5.200 ;
  RECT 2476.680 5.200 2476.900 5.400 ;
  RECT 2476.680 5.400 2476.880 7.020 ;
  RECT 2461.600 0.000 2462.400 1.000 ;
  RECT 2461.900 1.000 2462.100 5.200 ;
  RECT 2461.900 5.200 2462.250 5.400 ;
  RECT 2462.050 5.400 2462.250 7.020 ;
  RECT 2456.400 0.000 2457.200 1.000 ;
  RECT 2456.700 1.000 2456.900 5.200 ;
  RECT 2456.700 5.200 2457.040 5.400 ;
  RECT 2456.840 5.400 2457.040 7.020 ;
  RECT 2442.000 0.000 2442.800 1.000 ;
  RECT 2442.300 1.000 2442.500 5.200 ;
  RECT 2442.210 5.200 2442.500 5.400 ;
  RECT 2442.210 5.400 2442.410 7.020 ;
  RECT 2435.600 0.000 2436.400 1.000 ;
  RECT 2435.900 1.000 2436.100 5.200 ;
  RECT 2435.760 5.200 2436.100 5.400 ;
  RECT 2435.760 5.400 2435.960 7.020 ;
  RECT 2420.800 0.000 2421.600 1.000 ;
  RECT 2421.100 1.000 2421.300 5.200 ;
  RECT 2421.100 5.200 2421.330 5.400 ;
  RECT 2421.130 5.400 2421.330 7.020 ;
  RECT 2415.600 0.000 2416.400 1.000 ;
  RECT 2415.900 1.000 2416.100 5.200 ;
  RECT 2415.900 5.200 2416.120 5.400 ;
  RECT 2415.920 5.400 2416.120 7.020 ;
  RECT 2400.800 0.000 2401.600 1.000 ;
  RECT 2401.100 1.000 2401.300 5.200 ;
  RECT 2401.100 5.200 2401.490 5.400 ;
  RECT 2401.290 5.400 2401.490 7.020 ;
  RECT 2394.400 0.000 2395.200 1.000 ;
  RECT 2394.700 1.000 2394.900 5.200 ;
  RECT 2394.700 5.200 2395.040 5.400 ;
  RECT 2394.840 5.400 2395.040 7.020 ;
  RECT 2380.000 0.000 2380.800 1.000 ;
  RECT 2380.300 1.000 2380.500 5.200 ;
  RECT 2380.210 5.200 2380.500 5.400 ;
  RECT 2380.210 5.400 2380.410 7.020 ;
  RECT 2374.800 0.000 2375.600 1.000 ;
  RECT 2375.100 1.000 2375.300 5.200 ;
  RECT 2375.000 5.200 2375.300 5.400 ;
  RECT 2375.000 5.400 2375.200 7.020 ;
  RECT 2361.600 0.000 2362.400 1.000 ;
  RECT 2361.900 1.000 2362.100 5.200 ;
  RECT 2361.900 5.200 2362.290 5.400 ;
  RECT 2362.090 5.400 2362.290 7.020 ;
  RECT 2360.000 0.000 2360.800 1.000 ;
  RECT 2360.300 1.000 2360.500 5.200 ;
  RECT 2360.300 5.200 2360.570 5.400 ;
  RECT 2360.370 5.400 2360.570 7.020 ;
  RECT 2353.600 0.000 2354.400 1.000 ;
  RECT 2353.900 1.000 2354.100 5.200 ;
  RECT 2353.900 5.200 2354.120 5.400 ;
  RECT 2353.920 5.400 2354.120 7.020 ;
  RECT 2338.800 0.000 2339.600 1.000 ;
  RECT 2339.100 1.000 2339.300 5.200 ;
  RECT 2339.100 5.200 2339.490 5.400 ;
  RECT 2339.290 5.400 2339.490 7.020 ;
  RECT 2333.600 0.000 2334.400 1.000 ;
  RECT 2333.900 1.000 2334.100 5.200 ;
  RECT 2333.900 5.200 2334.280 5.400 ;
  RECT 2334.080 5.400 2334.280 7.020 ;
  RECT 2319.200 0.000 2320.000 1.000 ;
  RECT 2319.500 1.000 2319.700 5.200 ;
  RECT 2319.450 5.200 2319.700 5.400 ;
  RECT 2319.450 5.400 2319.650 7.020 ;
  RECT 2312.800 0.000 2313.600 1.000 ;
  RECT 2313.100 1.000 2313.300 5.200 ;
  RECT 2313.000 5.200 2313.300 5.400 ;
  RECT 2313.000 5.400 2313.200 7.020 ;
  RECT 2298.000 0.000 2298.800 1.000 ;
  RECT 2298.300 1.000 2298.500 5.200 ;
  RECT 2298.300 5.200 2298.570 5.400 ;
  RECT 2298.370 5.400 2298.570 7.020 ;
  RECT 2292.800 0.000 2293.600 1.000 ;
  RECT 2293.100 1.000 2293.300 5.200 ;
  RECT 2293.100 5.200 2293.360 5.400 ;
  RECT 2293.160 5.400 2293.360 7.020 ;
  RECT 2278.400 0.000 2279.200 1.000 ;
  RECT 2278.700 1.000 2278.900 5.200 ;
  RECT 2278.530 5.200 2278.900 5.400 ;
  RECT 2278.530 5.400 2278.730 7.020 ;
  RECT 2271.600 0.000 2272.400 1.000 ;
  RECT 2271.900 1.000 2272.100 5.200 ;
  RECT 2271.900 5.200 2272.280 5.400 ;
  RECT 2272.080 5.400 2272.280 7.020 ;
  RECT 2257.200 0.000 2258.000 1.000 ;
  RECT 2257.500 1.000 2257.700 5.200 ;
  RECT 2257.450 5.200 2257.700 5.400 ;
  RECT 2257.450 5.400 2257.650 7.020 ;
  RECT 2252.000 0.000 2252.800 1.000 ;
  RECT 2252.300 1.000 2252.500 5.200 ;
  RECT 2252.240 5.200 2252.500 5.400 ;
  RECT 2252.240 5.400 2252.440 7.020 ;
  RECT 2237.200 0.000 2238.000 1.000 ;
  RECT 2237.500 1.000 2237.700 5.200 ;
  RECT 2237.500 5.200 2237.810 5.400 ;
  RECT 2237.610 5.400 2237.810 7.020 ;
  RECT 2230.800 0.000 2231.600 1.000 ;
  RECT 2231.100 1.000 2231.300 5.200 ;
  RECT 2231.100 5.200 2231.360 5.400 ;
  RECT 2231.160 5.400 2231.360 7.020 ;
  RECT 2216.400 0.000 2217.200 1.000 ;
  RECT 2216.700 1.000 2216.900 5.200 ;
  RECT 2216.530 5.200 2216.900 5.400 ;
  RECT 2216.530 5.400 2216.730 7.020 ;
  RECT 2211.200 0.000 2212.000 1.000 ;
  RECT 2211.500 1.000 2211.700 5.200 ;
  RECT 2211.320 5.200 2211.700 5.400 ;
  RECT 2211.320 5.400 2211.520 7.020 ;
  RECT 2198.000 0.000 2198.800 1.000 ;
  RECT 2198.300 1.000 2198.500 5.200 ;
  RECT 2198.300 5.200 2198.610 5.400 ;
  RECT 2198.410 5.400 2198.610 7.020 ;
  RECT 2196.400 0.000 2197.200 1.000 ;
  RECT 2196.700 1.000 2196.900 5.200 ;
  RECT 2196.690 5.200 2196.900 5.400 ;
  RECT 2196.690 5.400 2196.890 7.020 ;
  RECT 2190.000 0.000 2190.800 1.000 ;
  RECT 2190.300 1.000 2190.500 5.200 ;
  RECT 2190.240 5.200 2190.500 5.400 ;
  RECT 2190.240 5.400 2190.440 7.020 ;
  RECT 2175.200 0.000 2176.000 1.000 ;
  RECT 2175.500 1.000 2175.700 5.200 ;
  RECT 2175.500 5.200 2175.810 5.400 ;
  RECT 2175.610 5.400 2175.810 7.020 ;
  RECT 2170.000 0.000 2170.800 1.000 ;
  RECT 2170.300 1.000 2170.500 5.200 ;
  RECT 2170.300 5.200 2170.600 5.400 ;
  RECT 2170.400 5.400 2170.600 7.020 ;
  RECT 2155.600 0.000 2156.400 1.000 ;
  RECT 2155.900 1.000 2156.100 5.200 ;
  RECT 2155.770 5.200 2156.100 5.400 ;
  RECT 2155.770 5.400 2155.970 7.020 ;
  RECT 2149.200 0.000 2150.000 1.000 ;
  RECT 2149.500 1.000 2149.700 5.200 ;
  RECT 2149.320 5.200 2149.700 5.400 ;
  RECT 2149.320 5.400 2149.520 7.020 ;
  RECT 2134.400 0.000 2135.200 1.000 ;
  RECT 2134.700 1.000 2134.900 5.200 ;
  RECT 2134.690 5.200 2134.900 5.400 ;
  RECT 2134.690 5.400 2134.890 7.020 ;
  RECT 2129.200 0.000 2130.000 1.000 ;
  RECT 2129.500 1.000 2129.700 5.200 ;
  RECT 2129.480 5.200 2129.700 5.400 ;
  RECT 2129.480 5.400 2129.680 7.020 ;
  RECT 2114.400 0.000 2115.200 1.000 ;
  RECT 2114.700 1.000 2114.900 5.200 ;
  RECT 2114.700 5.200 2115.050 5.400 ;
  RECT 2114.850 5.400 2115.050 7.020 ;
  RECT 2108.000 0.000 2108.800 1.000 ;
  RECT 2108.300 1.000 2108.500 5.200 ;
  RECT 2108.300 5.200 2108.600 5.400 ;
  RECT 2108.400 5.400 2108.600 7.020 ;
  RECT 2093.600 0.000 2094.400 1.000 ;
  RECT 2093.900 1.000 2094.100 5.200 ;
  RECT 2093.770 5.200 2094.100 5.400 ;
  RECT 2093.770 5.400 2093.970 7.020 ;
  RECT 2088.400 0.000 2089.200 1.000 ;
  RECT 2088.700 1.000 2088.900 5.200 ;
  RECT 2088.560 5.200 2088.900 5.400 ;
  RECT 2088.560 5.400 2088.760 7.020 ;
  RECT 2073.600 0.000 2074.400 1.000 ;
  RECT 2073.900 1.000 2074.100 5.200 ;
  RECT 2073.900 5.200 2074.130 5.400 ;
  RECT 2073.930 5.400 2074.130 7.020 ;
  RECT 2067.200 0.000 2068.000 1.000 ;
  RECT 2067.500 1.000 2067.700 5.200 ;
  RECT 2067.480 5.200 2067.700 5.400 ;
  RECT 2067.480 5.400 2067.680 7.020 ;
  RECT 2052.400 0.000 2053.200 1.000 ;
  RECT 2052.700 1.000 2052.900 5.200 ;
  RECT 2052.700 5.200 2053.050 5.400 ;
  RECT 2052.850 5.400 2053.050 7.020 ;
  RECT 2047.200 0.000 2048.000 1.000 ;
  RECT 2047.500 1.000 2047.700 5.200 ;
  RECT 2047.500 5.200 2047.840 5.400 ;
  RECT 2047.640 5.400 2047.840 7.020 ;
  RECT 2034.400 0.000 2035.200 1.000 ;
  RECT 2034.700 1.000 2034.900 5.200 ;
  RECT 2034.700 5.200 2034.930 5.400 ;
  RECT 2034.730 5.400 2034.930 7.020 ;
  RECT 2032.800 0.000 2033.600 1.000 ;
  RECT 2033.100 1.000 2033.300 5.200 ;
  RECT 2033.010 5.200 2033.300 5.400 ;
  RECT 2033.010 5.400 2033.210 7.020 ;
  RECT 2026.400 0.000 2027.200 1.000 ;
  RECT 2026.700 1.000 2026.900 5.200 ;
  RECT 2026.560 5.200 2026.900 5.400 ;
  RECT 2026.560 5.400 2026.760 7.020 ;
  RECT 2011.600 0.000 2012.400 1.000 ;
  RECT 2011.900 1.000 2012.100 5.200 ;
  RECT 2011.900 5.200 2012.130 5.400 ;
  RECT 2011.930 5.400 2012.130 7.020 ;
  RECT 2006.400 0.000 2007.200 1.000 ;
  RECT 2006.700 1.000 2006.900 5.200 ;
  RECT 2006.700 5.200 2006.920 5.400 ;
  RECT 2006.720 5.400 2006.920 7.020 ;
  RECT 1991.600 0.000 1992.400 1.000 ;
  RECT 1991.900 1.000 1992.100 5.200 ;
  RECT 1991.900 5.200 1992.290 5.400 ;
  RECT 1992.090 5.400 1992.290 7.020 ;
  RECT 1985.200 0.000 1986.000 1.000 ;
  RECT 1985.500 1.000 1985.700 5.200 ;
  RECT 1985.500 5.200 1985.840 5.400 ;
  RECT 1985.640 5.400 1985.840 7.020 ;
  RECT 1970.800 0.000 1971.600 1.000 ;
  RECT 1971.100 1.000 1971.300 5.200 ;
  RECT 1971.010 5.200 1971.300 5.400 ;
  RECT 1971.010 5.400 1971.210 7.020 ;
  RECT 1965.600 0.000 1966.400 1.000 ;
  RECT 1965.900 1.000 1966.100 5.200 ;
  RECT 1965.800 5.200 1966.100 5.400 ;
  RECT 1965.800 5.400 1966.000 7.020 ;
  RECT 1950.800 0.000 1951.600 1.000 ;
  RECT 1951.100 1.000 1951.300 5.200 ;
  RECT 1951.100 5.200 1951.370 5.400 ;
  RECT 1951.170 5.400 1951.370 7.020 ;
  RECT 1944.400 0.000 1945.200 1.000 ;
  RECT 1944.700 1.000 1944.900 5.200 ;
  RECT 1944.700 5.200 1944.920 5.400 ;
  RECT 1944.720 5.400 1944.920 7.020 ;
  RECT 1929.600 0.000 1930.400 1.000 ;
  RECT 1929.900 1.000 1930.100 5.200 ;
  RECT 1929.900 5.200 1930.290 5.400 ;
  RECT 1930.090 5.400 1930.290 7.020 ;
  RECT 1924.400 0.000 1925.200 1.000 ;
  RECT 1924.700 1.000 1924.900 5.200 ;
  RECT 1924.700 5.200 1925.080 5.400 ;
  RECT 1924.880 5.400 1925.080 7.020 ;
  RECT 1910.000 0.000 1910.800 1.000 ;
  RECT 1910.300 1.000 1910.500 5.200 ;
  RECT 1910.250 5.200 1910.500 5.400 ;
  RECT 1910.250 5.400 1910.450 7.020 ;
  RECT 1903.600 0.000 1904.400 1.000 ;
  RECT 1903.900 1.000 1904.100 5.200 ;
  RECT 1903.800 5.200 1904.100 5.400 ;
  RECT 1903.800 5.400 1904.000 7.020 ;
  RECT 1888.800 0.000 1889.600 1.000 ;
  RECT 1889.100 1.000 1889.300 5.200 ;
  RECT 1889.100 5.200 1889.370 5.400 ;
  RECT 1889.170 5.400 1889.370 7.020 ;
  RECT 1883.600 0.000 1884.400 1.000 ;
  RECT 1883.900 1.000 1884.100 5.200 ;
  RECT 1883.900 5.200 1884.160 5.400 ;
  RECT 1883.960 5.400 1884.160 7.020 ;
  RECT 1870.800 0.000 1871.600 1.000 ;
  RECT 1871.100 1.000 1871.300 5.200 ;
  RECT 1871.050 5.200 1871.300 5.400 ;
  RECT 1871.050 5.400 1871.250 7.020 ;
  RECT 1869.200 0.000 1870.000 1.000 ;
  RECT 1869.500 1.000 1869.700 5.200 ;
  RECT 1869.330 5.200 1869.700 5.400 ;
  RECT 1869.330 5.400 1869.530 7.020 ;
  RECT 1862.400 0.000 1863.200 1.000 ;
  RECT 1862.700 1.000 1862.900 5.200 ;
  RECT 1862.700 5.200 1863.080 5.400 ;
  RECT 1862.880 5.400 1863.080 7.020 ;
  RECT 1848.000 0.000 1848.800 1.000 ;
  RECT 1848.300 1.000 1848.500 5.200 ;
  RECT 1848.250 5.200 1848.500 5.400 ;
  RECT 1848.250 5.400 1848.450 7.020 ;
  RECT 1842.800 0.000 1843.600 1.000 ;
  RECT 1843.100 1.000 1843.300 5.200 ;
  RECT 1843.040 5.200 1843.300 5.400 ;
  RECT 1843.040 5.400 1843.240 7.020 ;
  RECT 1828.000 0.000 1828.800 1.000 ;
  RECT 1828.300 1.000 1828.500 5.200 ;
  RECT 1828.300 5.200 1828.610 5.400 ;
  RECT 1828.410 5.400 1828.610 7.020 ;
  RECT 1821.600 0.000 1822.400 1.000 ;
  RECT 1821.900 1.000 1822.100 5.200 ;
  RECT 1821.900 5.200 1822.160 5.400 ;
  RECT 1821.960 5.400 1822.160 7.020 ;
  RECT 1807.200 0.000 1808.000 1.000 ;
  RECT 1807.500 1.000 1807.700 5.200 ;
  RECT 1807.330 5.200 1807.700 5.400 ;
  RECT 1807.330 5.400 1807.530 7.020 ;
  RECT 1802.000 0.000 1802.800 1.000 ;
  RECT 1802.300 1.000 1802.500 5.200 ;
  RECT 1802.120 5.200 1802.500 5.400 ;
  RECT 1802.120 5.400 1802.320 7.020 ;
  RECT 1787.200 0.000 1788.000 1.000 ;
  RECT 1787.500 1.000 1787.700 5.200 ;
  RECT 1787.490 5.200 1787.700 5.400 ;
  RECT 1787.490 5.400 1787.690 7.020 ;
  RECT 1780.800 0.000 1781.600 1.000 ;
  RECT 1781.100 1.000 1781.300 5.200 ;
  RECT 1781.040 5.200 1781.300 5.400 ;
  RECT 1781.040 5.400 1781.240 7.020 ;
  RECT 1766.000 0.000 1766.800 1.000 ;
  RECT 1766.300 1.000 1766.500 5.200 ;
  RECT 1766.300 5.200 1766.610 5.400 ;
  RECT 1766.410 5.400 1766.610 7.020 ;
  RECT 1760.800 0.000 1761.600 1.000 ;
  RECT 1761.100 1.000 1761.300 5.200 ;
  RECT 1761.100 5.200 1761.400 5.400 ;
  RECT 1761.200 5.400 1761.400 7.020 ;
  RECT 1746.400 0.000 1747.200 1.000 ;
  RECT 1746.700 1.000 1746.900 5.200 ;
  RECT 1746.570 5.200 1746.900 5.400 ;
  RECT 1746.570 5.400 1746.770 7.020 ;
  RECT 1740.000 0.000 1740.800 1.000 ;
  RECT 1740.300 1.000 1740.500 5.200 ;
  RECT 1740.120 5.200 1740.500 5.400 ;
  RECT 1740.120 5.400 1740.320 7.020 ;
  RECT 1725.200 0.000 1726.000 1.000 ;
  RECT 1725.500 1.000 1725.700 5.200 ;
  RECT 1725.490 5.200 1725.700 5.400 ;
  RECT 1725.490 5.400 1725.690 7.020 ;
  RECT 1720.000 0.000 1720.800 1.000 ;
  RECT 1720.300 1.000 1720.500 5.200 ;
  RECT 1720.280 5.200 1720.500 5.400 ;
  RECT 1720.280 5.400 1720.480 7.020 ;
  RECT 1707.200 0.000 1708.000 1.000 ;
  RECT 1707.500 1.000 1707.700 5.200 ;
  RECT 1707.370 5.200 1707.700 5.400 ;
  RECT 1707.370 5.400 1707.570 7.020 ;
  RECT 1705.200 0.000 1706.000 1.000 ;
  RECT 1705.500 1.000 1705.700 5.200 ;
  RECT 1705.500 5.200 1705.850 5.400 ;
  RECT 1705.650 5.400 1705.850 7.020 ;
  RECT 1698.800 0.000 1699.600 1.000 ;
  RECT 1699.100 1.000 1699.300 5.200 ;
  RECT 1699.100 5.200 1699.400 5.400 ;
  RECT 1699.200 5.400 1699.400 7.020 ;
  RECT 1684.400 0.000 1685.200 1.000 ;
  RECT 1684.700 1.000 1684.900 5.200 ;
  RECT 1684.570 5.200 1684.900 5.400 ;
  RECT 1684.570 5.400 1684.770 7.020 ;
  RECT 1679.200 0.000 1680.000 1.000 ;
  RECT 1679.500 1.000 1679.700 5.200 ;
  RECT 1679.360 5.200 1679.700 5.400 ;
  RECT 1679.360 5.400 1679.560 7.020 ;
  RECT 1664.400 0.000 1665.200 1.000 ;
  RECT 1664.700 1.000 1664.900 5.200 ;
  RECT 1664.700 5.200 1664.930 5.400 ;
  RECT 1664.730 5.400 1664.930 7.020 ;
  RECT 1658.000 0.000 1658.800 1.000 ;
  RECT 1658.300 1.000 1658.500 5.200 ;
  RECT 1658.280 5.200 1658.500 5.400 ;
  RECT 1658.280 5.400 1658.480 7.020 ;
  RECT 1643.200 0.000 1644.000 1.000 ;
  RECT 1643.500 1.000 1643.700 5.200 ;
  RECT 1643.500 5.200 1643.850 5.400 ;
  RECT 1643.650 5.400 1643.850 7.020 ;
  RECT 1638.000 0.000 1638.800 1.000 ;
  RECT 1638.300 1.000 1638.500 5.200 ;
  RECT 1638.300 5.200 1638.640 5.400 ;
  RECT 1638.440 5.400 1638.640 7.020 ;
  RECT 1623.600 0.000 1624.400 1.000 ;
  RECT 1623.900 1.000 1624.100 5.200 ;
  RECT 1623.810 5.200 1624.100 5.400 ;
  RECT 1623.810 5.400 1624.010 7.020 ;
  RECT 1617.200 0.000 1618.000 1.000 ;
  RECT 1617.500 1.000 1617.700 5.200 ;
  RECT 1617.360 5.200 1617.700 5.400 ;
  RECT 1617.360 5.400 1617.560 7.020 ;
  RECT 1602.400 0.000 1603.200 1.000 ;
  RECT 1602.700 1.000 1602.900 5.200 ;
  RECT 1602.700 5.200 1602.930 5.400 ;
  RECT 1602.730 5.400 1602.930 7.020 ;
  RECT 1597.200 0.000 1598.000 1.000 ;
  RECT 1597.500 1.000 1597.700 5.200 ;
  RECT 1597.500 5.200 1597.720 5.400 ;
  RECT 1597.520 5.400 1597.720 7.020 ;
  RECT 1582.400 0.000 1583.200 1.000 ;
  RECT 1582.700 1.000 1582.900 5.200 ;
  RECT 1582.700 5.200 1583.090 5.400 ;
  RECT 1582.890 5.400 1583.090 7.020 ;
  RECT 1576.000 0.000 1576.800 1.000 ;
  RECT 1576.300 1.000 1576.500 5.200 ;
  RECT 1576.300 5.200 1576.640 5.400 ;
  RECT 1576.440 5.400 1576.640 7.020 ;
  RECT 1561.600 0.000 1562.400 1.000 ;
  RECT 1561.900 1.000 1562.100 5.200 ;
  RECT 1561.810 5.200 1562.100 5.400 ;
  RECT 1561.810 5.400 1562.010 7.020 ;
  RECT 1556.400 0.000 1557.200 1.000 ;
  RECT 1556.700 1.000 1556.900 5.200 ;
  RECT 1556.600 5.200 1556.900 5.400 ;
  RECT 1556.600 5.400 1556.800 7.020 ;
  RECT 1543.200 0.000 1544.000 1.000 ;
  RECT 1543.500 1.000 1543.700 5.200 ;
  RECT 1543.500 5.200 1543.890 5.400 ;
  RECT 1543.690 5.400 1543.890 7.020 ;
  RECT 1541.600 0.000 1542.400 1.000 ;
  RECT 1541.900 1.000 1542.100 5.200 ;
  RECT 1541.900 5.200 1542.170 5.400 ;
  RECT 1541.970 5.400 1542.170 7.020 ;
  RECT 1535.200 0.000 1536.000 1.000 ;
  RECT 1535.500 1.000 1535.700 5.200 ;
  RECT 1535.500 5.200 1535.720 5.400 ;
  RECT 1535.520 5.400 1535.720 7.020 ;
  RECT 1520.400 0.000 1521.200 1.000 ;
  RECT 1520.700 1.000 1520.900 5.200 ;
  RECT 1520.700 5.200 1521.090 5.400 ;
  RECT 1520.890 5.400 1521.090 7.020 ;
  RECT 1515.200 0.000 1516.000 1.000 ;
  RECT 1515.500 1.000 1515.700 5.200 ;
  RECT 1515.500 5.200 1515.880 5.400 ;
  RECT 1515.680 5.400 1515.880 7.020 ;
  RECT 1500.800 0.000 1501.600 1.000 ;
  RECT 1501.100 1.000 1501.300 5.200 ;
  RECT 1501.050 5.200 1501.300 5.400 ;
  RECT 1501.050 5.400 1501.250 7.020 ;
  RECT 1494.400 0.000 1495.200 1.000 ;
  RECT 1494.700 1.000 1494.900 5.200 ;
  RECT 1494.600 5.200 1494.900 5.400 ;
  RECT 1494.600 5.400 1494.800 7.020 ;
  RECT 1479.600 0.000 1480.400 1.000 ;
  RECT 1479.900 1.000 1480.100 5.200 ;
  RECT 1479.900 5.200 1480.170 5.400 ;
  RECT 1479.970 5.400 1480.170 7.020 ;
  RECT 1474.400 0.000 1475.200 1.000 ;
  RECT 1474.700 1.000 1474.900 5.200 ;
  RECT 1474.700 5.200 1474.960 5.400 ;
  RECT 1474.760 5.400 1474.960 7.020 ;
  RECT 1460.000 0.000 1460.800 1.000 ;
  RECT 1460.300 1.000 1460.500 5.200 ;
  RECT 1460.130 5.200 1460.500 5.400 ;
  RECT 1460.130 5.400 1460.330 7.020 ;
  RECT 1453.200 0.000 1454.000 1.000 ;
  RECT 1453.500 1.000 1453.700 5.200 ;
  RECT 1453.500 5.200 1453.880 5.400 ;
  RECT 1453.680 5.400 1453.880 7.020 ;
  RECT 1438.800 0.000 1439.600 1.000 ;
  RECT 1439.100 1.000 1439.300 5.200 ;
  RECT 1439.050 5.200 1439.300 5.400 ;
  RECT 1439.050 5.400 1439.250 7.020 ;
  RECT 1433.600 0.000 1434.400 1.000 ;
  RECT 1433.900 1.000 1434.100 5.200 ;
  RECT 1433.840 5.200 1434.100 5.400 ;
  RECT 1433.840 5.400 1434.040 7.020 ;
  RECT 1418.800 0.000 1419.600 1.000 ;
  RECT 1419.100 1.000 1419.300 5.200 ;
  RECT 1419.100 5.200 1419.410 5.400 ;
  RECT 1419.210 5.400 1419.410 7.020 ;
  RECT 1412.400 0.000 1413.200 1.000 ;
  RECT 1412.700 1.000 1412.900 5.200 ;
  RECT 1412.700 5.200 1412.960 5.400 ;
  RECT 1412.760 5.400 1412.960 7.020 ;
  RECT 1398.000 0.000 1398.800 1.000 ;
  RECT 1398.300 1.000 1398.500 5.200 ;
  RECT 1398.130 5.200 1398.500 5.400 ;
  RECT 1398.130 5.400 1398.330 7.020 ;
  RECT 1392.800 0.000 1393.600 1.000 ;
  RECT 1393.100 1.000 1393.300 5.200 ;
  RECT 1392.920 5.200 1393.300 5.400 ;
  RECT 1392.920 5.400 1393.120 7.020 ;
  RECT 1379.600 0.000 1380.400 1.000 ;
  RECT 1379.900 1.000 1380.100 5.200 ;
  RECT 1379.900 5.200 1380.210 5.400 ;
  RECT 1380.010 5.400 1380.210 7.020 ;
  RECT 1378.000 0.000 1378.800 1.000 ;
  RECT 1378.300 1.000 1378.500 5.200 ;
  RECT 1378.290 5.200 1378.500 5.400 ;
  RECT 1378.290 5.400 1378.490 7.020 ;
  RECT 1357.200 0.000 1358.000 1.000 ;
  RECT 1357.500 1.000 1357.700 5.200 ;
  RECT 1357.500 5.200 1357.720 5.400 ;
  RECT 1357.520 5.400 1357.720 7.020 ;
  RECT 1356.000 0.000 1356.800 1.000 ;
  RECT 1356.300 1.000 1356.500 5.200 ;
  RECT 1356.300 5.200 1356.570 5.400 ;
  RECT 1356.370 5.400 1356.570 7.020 ;
  RECT 1354.800 0.000 1355.600 1.000 ;
  RECT 1355.100 1.000 1355.300 5.200 ;
  RECT 1355.100 5.200 1355.400 5.400 ;
  RECT 1355.200 5.400 1355.400 7.020 ;
  RECT 1353.600 0.000 1354.400 1.000 ;
  RECT 1353.900 1.000 1354.100 5.200 ;
  RECT 1353.900 5.200 1354.150 5.400 ;
  RECT 1353.950 5.400 1354.150 7.020 ;
  RECT 1352.400 0.000 1353.200 1.000 ;
  RECT 1352.700 1.000 1352.900 5.200 ;
  RECT 1352.700 5.200 1352.900 5.400 ;
  RECT 1352.700 5.400 1352.900 7.020 ;
  RECT 1351.200 0.000 1352.000 1.000 ;
  RECT 1351.500 1.000 1351.700 5.200 ;
  RECT 1351.450 5.200 1351.700 5.400 ;
  RECT 1351.450 5.400 1351.650 7.020 ;
  RECT 1345.200 0.000 1346.000 1.000 ;
  RECT 1345.500 1.000 1345.700 5.200 ;
  RECT 1345.480 5.200 1345.700 5.400 ;
  RECT 1345.480 5.400 1345.680 7.020 ;
  RECT 1338.000 0.000 1338.800 1.000 ;
  RECT 1338.300 1.000 1338.500 5.200 ;
  RECT 1338.180 5.200 1338.500 5.400 ;
  RECT 1338.180 5.400 1338.380 7.020 ;
  RECT 1335.200 0.000 1336.000 1.000 ;
  RECT 1335.500 1.000 1335.700 5.200 ;
  RECT 1335.500 5.200 1335.900 5.400 ;
  RECT 1335.700 5.400 1335.900 7.020 ;
  RECT 1332.400 0.000 1333.200 1.000 ;
  RECT 1332.700 1.000 1332.900 5.200 ;
  RECT 1332.700 5.200 1333.040 5.400 ;
  RECT 1332.840 5.400 1333.040 7.020 ;
  RECT 1330.000 0.000 1330.800 1.000 ;
  RECT 1330.300 1.000 1330.500 5.200 ;
  RECT 1330.300 5.200 1330.560 5.400 ;
  RECT 1330.360 5.400 1330.560 7.020 ;
  RECT 1328.400 0.000 1329.200 1.000 ;
  RECT 1328.700 1.000 1328.900 5.200 ;
  RECT 1328.700 5.200 1329.040 5.400 ;
  RECT 1328.840 5.400 1329.040 7.020 ;
  RECT 1326.000 0.000 1326.800 1.000 ;
  RECT 1326.300 1.000 1326.500 5.200 ;
  RECT 1326.300 5.200 1326.560 5.400 ;
  RECT 1326.360 5.400 1326.560 7.020 ;
  RECT 1324.400 0.000 1325.200 1.000 ;
  RECT 1324.700 1.000 1324.900 5.200 ;
  RECT 1324.700 5.200 1325.040 5.400 ;
  RECT 1324.840 5.400 1325.040 7.020 ;
  RECT 1322.000 0.000 1322.800 1.000 ;
  RECT 1322.300 1.000 1322.500 5.200 ;
  RECT 1322.300 5.200 1322.560 5.400 ;
  RECT 1322.360 5.400 1322.560 7.020 ;
  RECT 1320.400 0.000 1321.200 1.000 ;
  RECT 1320.700 1.000 1320.900 5.200 ;
  RECT 1320.700 5.200 1321.040 5.400 ;
  RECT 1320.840 5.400 1321.040 7.020 ;
  RECT 1311.200 0.000 1312.000 1.000 ;
  RECT 1311.500 1.000 1311.700 5.200 ;
  RECT 1311.460 5.200 1311.700 5.400 ;
  RECT 1311.460 5.400 1311.660 7.020 ;
  RECT 1296.400 0.000 1297.200 1.000 ;
  RECT 1296.700 1.000 1296.900 5.200 ;
  RECT 1296.700 5.200 1297.030 5.400 ;
  RECT 1296.830 5.400 1297.030 7.020 ;
  RECT 1291.200 0.000 1292.000 1.000 ;
  RECT 1291.500 1.000 1291.700 5.200 ;
  RECT 1291.500 5.200 1291.820 5.400 ;
  RECT 1291.620 5.400 1291.820 7.020 ;
  RECT 1276.800 0.000 1277.600 1.000 ;
  RECT 1277.100 1.000 1277.300 5.200 ;
  RECT 1276.990 5.200 1277.300 5.400 ;
  RECT 1276.990 5.400 1277.190 7.020 ;
  RECT 1270.400 0.000 1271.200 1.000 ;
  RECT 1270.700 1.000 1270.900 5.200 ;
  RECT 1270.540 5.200 1270.900 5.400 ;
  RECT 1270.540 5.400 1270.740 7.020 ;
  RECT 1255.600 0.000 1256.400 1.000 ;
  RECT 1255.900 1.000 1256.100 5.200 ;
  RECT 1255.900 5.200 1256.110 5.400 ;
  RECT 1255.910 5.400 1256.110 7.020 ;
  RECT 1250.400 0.000 1251.200 1.000 ;
  RECT 1250.700 1.000 1250.900 5.200 ;
  RECT 1250.700 5.200 1250.900 5.400 ;
  RECT 1250.700 5.400 1250.900 7.020 ;
  RECT 1235.600 0.000 1236.400 1.000 ;
  RECT 1235.900 1.000 1236.100 5.200 ;
  RECT 1235.900 5.200 1236.270 5.400 ;
  RECT 1236.070 5.400 1236.270 7.020 ;
  RECT 1229.200 0.000 1230.000 1.000 ;
  RECT 1229.500 1.000 1229.700 5.200 ;
  RECT 1229.500 5.200 1229.820 5.400 ;
  RECT 1229.620 5.400 1229.820 7.020 ;
  RECT 1214.800 0.000 1215.600 1.000 ;
  RECT 1215.100 1.000 1215.300 5.200 ;
  RECT 1214.990 5.200 1215.300 5.400 ;
  RECT 1214.990 5.400 1215.190 7.020 ;
  RECT 1209.600 0.000 1210.400 1.000 ;
  RECT 1209.900 1.000 1210.100 5.200 ;
  RECT 1209.780 5.200 1210.100 5.400 ;
  RECT 1209.780 5.400 1209.980 7.020 ;
  RECT 1194.800 0.000 1195.600 1.000 ;
  RECT 1195.100 1.000 1195.300 5.200 ;
  RECT 1195.100 5.200 1195.350 5.400 ;
  RECT 1195.150 5.400 1195.350 7.020 ;
  RECT 1188.400 0.000 1189.200 1.000 ;
  RECT 1188.700 1.000 1188.900 5.200 ;
  RECT 1188.700 5.200 1188.900 5.400 ;
  RECT 1188.700 5.400 1188.900 7.020 ;
  RECT 1173.600 0.000 1174.400 1.000 ;
  RECT 1173.900 1.000 1174.100 5.200 ;
  RECT 1173.900 5.200 1174.270 5.400 ;
  RECT 1174.070 5.400 1174.270 7.020 ;
  RECT 1168.400 0.000 1169.200 1.000 ;
  RECT 1168.700 1.000 1168.900 5.200 ;
  RECT 1168.700 5.200 1169.060 5.400 ;
  RECT 1168.860 5.400 1169.060 7.020 ;
  RECT 1155.600 0.000 1156.400 1.000 ;
  RECT 1155.900 1.000 1156.100 5.200 ;
  RECT 1155.900 5.200 1156.150 5.400 ;
  RECT 1155.950 5.400 1156.150 7.020 ;
  RECT 1154.000 0.000 1154.800 1.000 ;
  RECT 1154.300 1.000 1154.500 5.200 ;
  RECT 1154.230 5.200 1154.500 5.400 ;
  RECT 1154.230 5.400 1154.430 7.020 ;
  RECT 1147.600 0.000 1148.400 1.000 ;
  RECT 1147.900 1.000 1148.100 5.200 ;
  RECT 1147.780 5.200 1148.100 5.400 ;
  RECT 1147.780 5.400 1147.980 7.020 ;
  RECT 1132.800 0.000 1133.600 1.000 ;
  RECT 1133.100 1.000 1133.300 5.200 ;
  RECT 1133.100 5.200 1133.350 5.400 ;
  RECT 1133.150 5.400 1133.350 7.020 ;
  RECT 1127.600 0.000 1128.400 1.000 ;
  RECT 1127.900 1.000 1128.100 5.200 ;
  RECT 1127.900 5.200 1128.140 5.400 ;
  RECT 1127.940 5.400 1128.140 7.020 ;
  RECT 1113.200 0.000 1114.000 1.000 ;
  RECT 1113.500 1.000 1113.700 5.200 ;
  RECT 1113.310 5.200 1113.700 5.400 ;
  RECT 1113.310 5.400 1113.510 7.020 ;
  RECT 1106.400 0.000 1107.200 1.000 ;
  RECT 1106.700 1.000 1106.900 5.200 ;
  RECT 1106.700 5.200 1107.060 5.400 ;
  RECT 1106.860 5.400 1107.060 7.020 ;
  RECT 1092.000 0.000 1092.800 1.000 ;
  RECT 1092.300 1.000 1092.500 5.200 ;
  RECT 1092.230 5.200 1092.500 5.400 ;
  RECT 1092.230 5.400 1092.430 7.020 ;
  RECT 1086.800 0.000 1087.600 1.000 ;
  RECT 1087.100 1.000 1087.300 5.200 ;
  RECT 1087.020 5.200 1087.300 5.400 ;
  RECT 1087.020 5.400 1087.220 7.020 ;
  RECT 1072.000 0.000 1072.800 1.000 ;
  RECT 1072.300 1.000 1072.500 5.200 ;
  RECT 1072.300 5.200 1072.590 5.400 ;
  RECT 1072.390 5.400 1072.590 7.020 ;
  RECT 1065.600 0.000 1066.400 1.000 ;
  RECT 1065.900 1.000 1066.100 5.200 ;
  RECT 1065.900 5.200 1066.140 5.400 ;
  RECT 1065.940 5.400 1066.140 7.020 ;
  RECT 1051.200 0.000 1052.000 1.000 ;
  RECT 1051.500 1.000 1051.700 5.200 ;
  RECT 1051.310 5.200 1051.700 5.400 ;
  RECT 1051.310 5.400 1051.510 7.020 ;
  RECT 1045.600 0.000 1046.400 1.000 ;
  RECT 1045.900 1.000 1046.100 5.200 ;
  RECT 1045.900 5.200 1046.300 5.400 ;
  RECT 1046.100 5.400 1046.300 7.020 ;
  RECT 1031.200 0.000 1032.000 1.000 ;
  RECT 1031.500 1.000 1031.700 5.200 ;
  RECT 1031.470 5.200 1031.700 5.400 ;
  RECT 1031.470 5.400 1031.670 7.020 ;
  RECT 1024.800 0.000 1025.600 1.000 ;
  RECT 1025.100 1.000 1025.300 5.200 ;
  RECT 1025.020 5.200 1025.300 5.400 ;
  RECT 1025.020 5.400 1025.220 7.020 ;
  RECT 1010.000 0.000 1010.800 1.000 ;
  RECT 1010.300 1.000 1010.500 5.200 ;
  RECT 1010.300 5.200 1010.590 5.400 ;
  RECT 1010.390 5.400 1010.590 7.020 ;
  RECT 1004.800 0.000 1005.600 1.000 ;
  RECT 1005.100 1.000 1005.300 5.200 ;
  RECT 1005.100 5.200 1005.380 5.400 ;
  RECT 1005.180 5.400 1005.380 7.020 ;
  RECT 992.000 0.000 992.800 1.000 ;
  RECT 992.300 1.000 992.500 5.200 ;
  RECT 992.270 5.200 992.500 5.400 ;
  RECT 992.270 5.400 992.470 7.020 ;
  RECT 990.400 0.000 991.200 1.000 ;
  RECT 990.700 1.000 990.900 5.200 ;
  RECT 990.550 5.200 990.900 5.400 ;
  RECT 990.550 5.400 990.750 7.020 ;
  RECT 983.600 0.000 984.400 1.000 ;
  RECT 983.900 1.000 984.100 5.200 ;
  RECT 983.900 5.200 984.300 5.400 ;
  RECT 984.100 5.400 984.300 7.020 ;
  RECT 969.200 0.000 970.000 1.000 ;
  RECT 969.500 1.000 969.700 5.200 ;
  RECT 969.470 5.200 969.700 5.400 ;
  RECT 969.470 5.400 969.670 7.020 ;
  RECT 964.000 0.000 964.800 1.000 ;
  RECT 964.300 1.000 964.500 5.200 ;
  RECT 964.260 5.200 964.500 5.400 ;
  RECT 964.260 5.400 964.460 7.020 ;
  RECT 949.200 0.000 950.000 1.000 ;
  RECT 949.500 1.000 949.700 5.200 ;
  RECT 949.500 5.200 949.830 5.400 ;
  RECT 949.630 5.400 949.830 7.020 ;
  RECT 942.800 0.000 943.600 1.000 ;
  RECT 943.100 1.000 943.300 5.200 ;
  RECT 943.100 5.200 943.380 5.400 ;
  RECT 943.180 5.400 943.380 7.020 ;
  RECT 928.400 0.000 929.200 1.000 ;
  RECT 928.700 1.000 928.900 5.200 ;
  RECT 928.550 5.200 928.900 5.400 ;
  RECT 928.550 5.400 928.750 7.020 ;
  RECT 923.200 0.000 924.000 1.000 ;
  RECT 923.500 1.000 923.700 5.200 ;
  RECT 923.340 5.200 923.700 5.400 ;
  RECT 923.340 5.400 923.540 7.020 ;
  RECT 908.400 0.000 909.200 1.000 ;
  RECT 908.700 1.000 908.900 5.200 ;
  RECT 908.700 5.200 908.910 5.400 ;
  RECT 908.710 5.400 908.910 7.020 ;
  RECT 902.000 0.000 902.800 1.000 ;
  RECT 902.300 1.000 902.500 5.200 ;
  RECT 902.260 5.200 902.500 5.400 ;
  RECT 902.260 5.400 902.460 7.020 ;
  RECT 887.200 0.000 888.000 1.000 ;
  RECT 887.500 1.000 887.700 5.200 ;
  RECT 887.500 5.200 887.830 5.400 ;
  RECT 887.630 5.400 887.830 7.020 ;
  RECT 882.000 0.000 882.800 1.000 ;
  RECT 882.300 1.000 882.500 5.200 ;
  RECT 882.300 5.200 882.620 5.400 ;
  RECT 882.420 5.400 882.620 7.020 ;
  RECT 867.600 0.000 868.400 1.000 ;
  RECT 867.900 1.000 868.100 5.200 ;
  RECT 867.790 5.200 868.100 5.400 ;
  RECT 867.790 5.400 867.990 7.020 ;
  RECT 861.200 0.000 862.000 1.000 ;
  RECT 861.500 1.000 861.700 5.200 ;
  RECT 861.340 5.200 861.700 5.400 ;
  RECT 861.340 5.400 861.540 7.020 ;
  RECT 846.400 0.000 847.200 1.000 ;
  RECT 846.700 1.000 846.900 5.200 ;
  RECT 846.700 5.200 846.910 5.400 ;
  RECT 846.710 5.400 846.910 7.020 ;
  RECT 841.200 0.000 842.000 1.000 ;
  RECT 841.500 1.000 841.700 5.200 ;
  RECT 841.500 5.200 841.700 5.400 ;
  RECT 841.500 5.400 841.700 7.020 ;
  RECT 828.400 0.000 829.200 1.000 ;
  RECT 828.700 1.000 828.900 5.200 ;
  RECT 828.590 5.200 828.900 5.400 ;
  RECT 828.590 5.400 828.790 7.020 ;
  RECT 826.400 0.000 827.200 1.000 ;
  RECT 826.700 1.000 826.900 5.200 ;
  RECT 826.700 5.200 827.070 5.400 ;
  RECT 826.870 5.400 827.070 7.020 ;
  RECT 820.000 0.000 820.800 1.000 ;
  RECT 820.300 1.000 820.500 5.200 ;
  RECT 820.300 5.200 820.620 5.400 ;
  RECT 820.420 5.400 820.620 7.020 ;
  RECT 805.600 0.000 806.400 1.000 ;
  RECT 805.900 1.000 806.100 5.200 ;
  RECT 805.790 5.200 806.100 5.400 ;
  RECT 805.790 5.400 805.990 7.020 ;
  RECT 800.400 0.000 801.200 1.000 ;
  RECT 800.700 1.000 800.900 5.200 ;
  RECT 800.580 5.200 800.900 5.400 ;
  RECT 800.580 5.400 800.780 7.020 ;
  RECT 785.600 0.000 786.400 1.000 ;
  RECT 785.900 1.000 786.100 5.200 ;
  RECT 785.900 5.200 786.150 5.400 ;
  RECT 785.950 5.400 786.150 7.020 ;
  RECT 779.200 0.000 780.000 1.000 ;
  RECT 779.500 1.000 779.700 5.200 ;
  RECT 779.500 5.200 779.700 5.400 ;
  RECT 779.500 5.400 779.700 7.020 ;
  RECT 764.400 0.000 765.200 1.000 ;
  RECT 764.700 1.000 764.900 5.200 ;
  RECT 764.700 5.200 765.070 5.400 ;
  RECT 764.870 5.400 765.070 7.020 ;
  RECT 759.200 0.000 760.000 1.000 ;
  RECT 759.500 1.000 759.700 5.200 ;
  RECT 759.500 5.200 759.860 5.400 ;
  RECT 759.660 5.400 759.860 7.020 ;
  RECT 744.800 0.000 745.600 1.000 ;
  RECT 745.100 1.000 745.300 5.200 ;
  RECT 745.030 5.200 745.300 5.400 ;
  RECT 745.030 5.400 745.230 7.020 ;
  RECT 738.400 0.000 739.200 1.000 ;
  RECT 738.700 1.000 738.900 5.200 ;
  RECT 738.580 5.200 738.900 5.400 ;
  RECT 738.580 5.400 738.780 7.020 ;
  RECT 723.600 0.000 724.400 1.000 ;
  RECT 723.900 1.000 724.100 5.200 ;
  RECT 723.900 5.200 724.150 5.400 ;
  RECT 723.950 5.400 724.150 7.020 ;
  RECT 718.400 0.000 719.200 1.000 ;
  RECT 718.700 1.000 718.900 5.200 ;
  RECT 718.700 5.200 718.940 5.400 ;
  RECT 718.740 5.400 718.940 7.020 ;
  RECT 704.000 0.000 704.800 1.000 ;
  RECT 704.300 1.000 704.500 5.200 ;
  RECT 704.110 5.200 704.500 5.400 ;
  RECT 704.110 5.400 704.310 7.020 ;
  RECT 697.200 0.000 698.000 1.000 ;
  RECT 697.500 1.000 697.700 5.200 ;
  RECT 697.500 5.200 697.860 5.400 ;
  RECT 697.660 5.400 697.860 7.020 ;
  RECT 682.800 0.000 683.600 1.000 ;
  RECT 683.100 1.000 683.300 5.200 ;
  RECT 683.030 5.200 683.300 5.400 ;
  RECT 683.030 5.400 683.230 7.020 ;
  RECT 677.600 0.000 678.400 1.000 ;
  RECT 677.900 1.000 678.100 5.200 ;
  RECT 677.820 5.200 678.100 5.400 ;
  RECT 677.820 5.400 678.020 7.020 ;
  RECT 664.800 0.000 665.600 1.000 ;
  RECT 665.100 1.000 665.300 5.200 ;
  RECT 664.910 5.200 665.300 5.400 ;
  RECT 664.910 5.400 665.110 7.020 ;
  RECT 662.800 0.000 663.600 1.000 ;
  RECT 663.100 1.000 663.300 5.200 ;
  RECT 663.100 5.200 663.390 5.400 ;
  RECT 663.190 5.400 663.390 7.020 ;
  RECT 656.400 0.000 657.200 1.000 ;
  RECT 656.700 1.000 656.900 5.200 ;
  RECT 656.700 5.200 656.940 5.400 ;
  RECT 656.740 5.400 656.940 7.020 ;
  RECT 642.000 0.000 642.800 1.000 ;
  RECT 642.300 1.000 642.500 5.200 ;
  RECT 642.110 5.200 642.500 5.400 ;
  RECT 642.110 5.400 642.310 7.020 ;
  RECT 636.400 0.000 637.200 1.000 ;
  RECT 636.700 1.000 636.900 5.200 ;
  RECT 636.700 5.200 637.100 5.400 ;
  RECT 636.900 5.400 637.100 7.020 ;
  RECT 622.000 0.000 622.800 1.000 ;
  RECT 622.300 1.000 622.500 5.200 ;
  RECT 622.270 5.200 622.500 5.400 ;
  RECT 622.270 5.400 622.470 7.020 ;
  RECT 615.600 0.000 616.400 1.000 ;
  RECT 615.900 1.000 616.100 5.200 ;
  RECT 615.820 5.200 616.100 5.400 ;
  RECT 615.820 5.400 616.020 7.020 ;
  RECT 600.800 0.000 601.600 1.000 ;
  RECT 601.100 1.000 601.300 5.200 ;
  RECT 601.100 5.200 601.390 5.400 ;
  RECT 601.190 5.400 601.390 7.020 ;
  RECT 595.600 0.000 596.400 1.000 ;
  RECT 595.900 1.000 596.100 5.200 ;
  RECT 595.900 5.200 596.180 5.400 ;
  RECT 595.980 5.400 596.180 7.020 ;
  RECT 581.200 0.000 582.000 1.000 ;
  RECT 581.500 1.000 581.700 5.200 ;
  RECT 581.350 5.200 581.700 5.400 ;
  RECT 581.350 5.400 581.550 7.020 ;
  RECT 574.400 0.000 575.200 1.000 ;
  RECT 574.700 1.000 574.900 5.200 ;
  RECT 574.700 5.200 575.100 5.400 ;
  RECT 574.900 5.400 575.100 7.020 ;
  RECT 560.000 0.000 560.800 1.000 ;
  RECT 560.300 1.000 560.500 5.200 ;
  RECT 560.270 5.200 560.500 5.400 ;
  RECT 560.270 5.400 560.470 7.020 ;
  RECT 554.800 0.000 555.600 1.000 ;
  RECT 555.100 1.000 555.300 5.200 ;
  RECT 555.060 5.200 555.300 5.400 ;
  RECT 555.060 5.400 555.260 7.020 ;
  RECT 540.000 0.000 540.800 1.000 ;
  RECT 540.300 1.000 540.500 5.200 ;
  RECT 540.300 5.200 540.630 5.400 ;
  RECT 540.430 5.400 540.630 7.020 ;
  RECT 533.600 0.000 534.400 1.000 ;
  RECT 533.900 1.000 534.100 5.200 ;
  RECT 533.900 5.200 534.180 5.400 ;
  RECT 533.980 5.400 534.180 7.020 ;
  RECT 519.200 0.000 520.000 1.000 ;
  RECT 519.500 1.000 519.700 5.200 ;
  RECT 519.350 5.200 519.700 5.400 ;
  RECT 519.350 5.400 519.550 7.020 ;
  RECT 514.000 0.000 514.800 1.000 ;
  RECT 514.300 1.000 514.500 5.200 ;
  RECT 514.140 5.200 514.500 5.400 ;
  RECT 514.140 5.400 514.340 7.020 ;
  RECT 500.800 0.000 501.600 1.000 ;
  RECT 501.100 1.000 501.300 5.200 ;
  RECT 501.100 5.200 501.430 5.400 ;
  RECT 501.230 5.400 501.430 7.020 ;
  RECT 499.200 0.000 500.000 1.000 ;
  RECT 499.500 1.000 499.700 5.200 ;
  RECT 499.500 5.200 499.710 5.400 ;
  RECT 499.510 5.400 499.710 7.020 ;
  RECT 492.800 0.000 493.600 1.000 ;
  RECT 493.100 1.000 493.300 5.200 ;
  RECT 493.060 5.200 493.300 5.400 ;
  RECT 493.060 5.400 493.260 7.020 ;
  RECT 478.000 0.000 478.800 1.000 ;
  RECT 478.300 1.000 478.500 5.200 ;
  RECT 478.300 5.200 478.630 5.400 ;
  RECT 478.430 5.400 478.630 7.020 ;
  RECT 472.800 0.000 473.600 1.000 ;
  RECT 473.100 1.000 473.300 5.200 ;
  RECT 473.100 5.200 473.420 5.400 ;
  RECT 473.220 5.400 473.420 7.020 ;
  RECT 458.400 0.000 459.200 1.000 ;
  RECT 458.700 1.000 458.900 5.200 ;
  RECT 458.590 5.200 458.900 5.400 ;
  RECT 458.590 5.400 458.790 7.020 ;
  RECT 452.000 0.000 452.800 1.000 ;
  RECT 452.300 1.000 452.500 5.200 ;
  RECT 452.140 5.200 452.500 5.400 ;
  RECT 452.140 5.400 452.340 7.020 ;
  RECT 437.200 0.000 438.000 1.000 ;
  RECT 437.500 1.000 437.700 5.200 ;
  RECT 437.500 5.200 437.710 5.400 ;
  RECT 437.510 5.400 437.710 7.020 ;
  RECT 432.000 0.000 432.800 1.000 ;
  RECT 432.300 1.000 432.500 5.200 ;
  RECT 432.300 5.200 432.500 5.400 ;
  RECT 432.300 5.400 432.500 7.020 ;
  RECT 417.200 0.000 418.000 1.000 ;
  RECT 417.500 1.000 417.700 5.200 ;
  RECT 417.500 5.200 417.870 5.400 ;
  RECT 417.670 5.400 417.870 7.020 ;
  RECT 410.800 0.000 411.600 1.000 ;
  RECT 411.100 1.000 411.300 5.200 ;
  RECT 411.100 5.200 411.420 5.400 ;
  RECT 411.220 5.400 411.420 7.020 ;
  RECT 396.400 0.000 397.200 1.000 ;
  RECT 396.700 1.000 396.900 5.200 ;
  RECT 396.590 5.200 396.900 5.400 ;
  RECT 396.590 5.400 396.790 7.020 ;
  RECT 391.200 0.000 392.000 1.000 ;
  RECT 391.500 1.000 391.700 5.200 ;
  RECT 391.380 5.200 391.700 5.400 ;
  RECT 391.380 5.400 391.580 7.020 ;
  RECT 376.400 0.000 377.200 1.000 ;
  RECT 376.700 1.000 376.900 5.200 ;
  RECT 376.700 5.200 376.950 5.400 ;
  RECT 376.750 5.400 376.950 7.020 ;
  RECT 370.000 0.000 370.800 1.000 ;
  RECT 370.300 1.000 370.500 5.200 ;
  RECT 370.300 5.200 370.500 5.400 ;
  RECT 370.300 5.400 370.500 7.020 ;
  RECT 355.200 0.000 356.000 1.000 ;
  RECT 355.500 1.000 355.700 5.200 ;
  RECT 355.500 5.200 355.870 5.400 ;
  RECT 355.670 5.400 355.870 7.020 ;
  RECT 350.000 0.000 350.800 1.000 ;
  RECT 350.300 1.000 350.500 5.200 ;
  RECT 350.300 5.200 350.660 5.400 ;
  RECT 350.460 5.400 350.660 7.020 ;
  RECT 337.200 0.000 338.000 1.000 ;
  RECT 337.500 1.000 337.700 5.200 ;
  RECT 337.500 5.200 337.750 5.400 ;
  RECT 337.550 5.400 337.750 7.020 ;
  RECT 335.600 0.000 336.400 1.000 ;
  RECT 335.900 1.000 336.100 5.200 ;
  RECT 335.830 5.200 336.100 5.400 ;
  RECT 335.830 5.400 336.030 7.020 ;
  RECT 329.200 0.000 330.000 1.000 ;
  RECT 329.500 1.000 329.700 5.200 ;
  RECT 329.380 5.200 329.700 5.400 ;
  RECT 329.380 5.400 329.580 7.020 ;
  RECT 314.400 0.000 315.200 1.000 ;
  RECT 314.700 1.000 314.900 5.200 ;
  RECT 314.700 5.200 314.950 5.400 ;
  RECT 314.750 5.400 314.950 7.020 ;
  RECT 309.200 0.000 310.000 1.000 ;
  RECT 309.500 1.000 309.700 5.200 ;
  RECT 309.500 5.200 309.740 5.400 ;
  RECT 309.540 5.400 309.740 7.020 ;
  RECT 294.800 0.000 295.600 1.000 ;
  RECT 295.100 1.000 295.300 5.200 ;
  RECT 294.910 5.200 295.300 5.400 ;
  RECT 294.910 5.400 295.110 7.020 ;
  RECT 288.000 0.000 288.800 1.000 ;
  RECT 288.300 1.000 288.500 5.200 ;
  RECT 288.300 5.200 288.660 5.400 ;
  RECT 288.460 5.400 288.660 7.020 ;
  RECT 273.600 0.000 274.400 1.000 ;
  RECT 273.900 1.000 274.100 5.200 ;
  RECT 273.830 5.200 274.100 5.400 ;
  RECT 273.830 5.400 274.030 7.020 ;
  RECT 268.400 0.000 269.200 1.000 ;
  RECT 268.700 1.000 268.900 5.200 ;
  RECT 268.620 5.200 268.900 5.400 ;
  RECT 268.620 5.400 268.820 7.020 ;
  RECT 253.600 0.000 254.400 1.000 ;
  RECT 253.900 1.000 254.100 5.200 ;
  RECT 253.900 5.200 254.190 5.400 ;
  RECT 253.990 5.400 254.190 7.020 ;
  RECT 247.200 0.000 248.000 1.000 ;
  RECT 247.500 1.000 247.700 5.200 ;
  RECT 247.500 5.200 247.740 5.400 ;
  RECT 247.540 5.400 247.740 7.020 ;
  RECT 232.800 0.000 233.600 1.000 ;
  RECT 233.100 1.000 233.300 5.200 ;
  RECT 232.910 5.200 233.300 5.400 ;
  RECT 232.910 5.400 233.110 7.020 ;
  RECT 227.200 0.000 228.000 1.000 ;
  RECT 227.500 1.000 227.700 5.200 ;
  RECT 227.500 5.200 227.900 5.400 ;
  RECT 227.700 5.400 227.900 7.020 ;
  RECT 212.800 0.000 213.600 1.000 ;
  RECT 213.100 1.000 213.300 5.200 ;
  RECT 213.070 5.200 213.300 5.400 ;
  RECT 213.070 5.400 213.270 7.020 ;
  RECT 206.400 0.000 207.200 1.000 ;
  RECT 206.700 1.000 206.900 5.200 ;
  RECT 206.620 5.200 206.900 5.400 ;
  RECT 206.620 5.400 206.820 7.020 ;
  RECT 191.600 0.000 192.400 1.000 ;
  RECT 191.900 1.000 192.100 5.200 ;
  RECT 191.900 5.200 192.190 5.400 ;
  RECT 191.990 5.400 192.190 7.020 ;
  RECT 186.400 0.000 187.200 1.000 ;
  RECT 186.700 1.000 186.900 5.200 ;
  RECT 186.700 5.200 186.980 5.400 ;
  RECT 186.780 5.400 186.980 7.020 ;
  RECT 173.600 0.000 174.400 1.000 ;
  RECT 173.900 1.000 174.100 5.200 ;
  RECT 173.870 5.200 174.100 5.400 ;
  RECT 173.870 5.400 174.070 7.020 ;
  RECT 172.000 0.000 172.800 1.000 ;
  RECT 172.300 1.000 172.500 5.200 ;
  RECT 172.150 5.200 172.500 5.400 ;
  RECT 172.150 5.400 172.350 7.020 ;
  RECT 165.200 0.000 166.000 1.000 ;
  RECT 165.500 1.000 165.700 5.200 ;
  RECT 165.500 5.200 165.900 5.400 ;
  RECT 165.700 5.400 165.900 7.020 ;
  RECT 150.800 0.000 151.600 1.000 ;
  RECT 151.100 1.000 151.300 5.200 ;
  RECT 151.070 5.200 151.300 5.400 ;
  RECT 151.070 5.400 151.270 7.020 ;
  RECT 145.600 0.000 146.400 1.000 ;
  RECT 145.900 1.000 146.100 5.200 ;
  RECT 145.860 5.200 146.100 5.400 ;
  RECT 145.860 5.400 146.060 7.020 ;
  RECT 130.800 0.000 131.600 1.000 ;
  RECT 131.100 1.000 131.300 5.200 ;
  RECT 131.100 5.200 131.430 5.400 ;
  RECT 131.230 5.400 131.430 7.020 ;
  RECT 124.400 0.000 125.200 1.000 ;
  RECT 124.700 1.000 124.900 5.200 ;
  RECT 124.700 5.200 124.980 5.400 ;
  RECT 124.780 5.400 124.980 7.020 ;
  RECT 110.000 0.000 110.800 1.000 ;
  RECT 110.300 1.000 110.500 5.200 ;
  RECT 110.150 5.200 110.500 5.400 ;
  RECT 110.150 5.400 110.350 7.020 ;
  RECT 104.800 0.000 105.600 1.000 ;
  RECT 105.100 1.000 105.300 5.200 ;
  RECT 104.940 5.200 105.300 5.400 ;
  RECT 104.940 5.400 105.140 7.020 ;
  RECT 90.000 0.000 90.800 1.000 ;
  RECT 90.300 1.000 90.500 5.200 ;
  RECT 90.300 5.200 90.510 5.400 ;
  RECT 90.310 5.400 90.510 7.020 ;
  RECT 83.600 0.000 84.400 1.000 ;
  RECT 83.900 1.000 84.100 5.200 ;
  RECT 83.860 5.200 84.100 5.400 ;
  RECT 83.860 5.400 84.060 7.020 ;
  RECT 68.800 0.000 69.600 1.000 ;
  RECT 69.100 1.000 69.300 5.200 ;
  RECT 69.100 5.200 69.430 5.400 ;
  RECT 69.230 5.400 69.430 7.020 ;
  RECT 63.600 0.000 64.400 1.000 ;
  RECT 63.900 1.000 64.100 5.200 ;
  RECT 63.900 5.200 64.220 5.400 ;
  RECT 64.020 5.400 64.220 7.020 ;
  RECT 49.200 0.000 50.000 1.000 ;
  RECT 49.500 1.000 49.700 5.200 ;
  RECT 49.390 5.200 49.700 5.400 ;
  RECT 49.390 5.400 49.590 7.020 ;
  RECT 42.800 0.000 43.600 1.000 ;
  RECT 43.100 1.000 43.300 5.200 ;
  RECT 42.940 5.200 43.300 5.400 ;
  RECT 42.940 5.400 43.140 7.020 ;
  RECT 28.000 0.000 28.800 1.000 ;
  RECT 28.300 1.000 28.500 5.200 ;
  RECT 28.300 5.200 28.510 5.400 ;
  RECT 28.310 5.400 28.510 7.020 ;
  RECT 22.800 0.000 23.600 1.000 ;
  RECT 23.100 1.000 23.300 5.200 ;
  RECT 23.100 5.200 23.300 5.400 ;
  RECT 23.100 5.400 23.300 7.020 ;
  RECT 10.000 0.000 10.800 1.000 ;
  RECT 10.300 1.000 10.500 5.200 ;
  RECT 10.190 5.200 10.500 5.400 ;
  RECT 10.190 5.400 10.390 7.020 ;
  RECT 8.000 0.000 8.800 1.000 ;
  RECT 8.300 1.000 8.500 5.200 ;
  RECT 8.300 5.200 8.670 5.400 ;
  RECT 8.470 5.400 8.670 7.020 ;
  RECT 2687.520 9.570 2688.660 11.170 ;
  RECT 2687.520 14.200 2688.660 15.200 ;
  RECT 2687.520 18.730 2688.660 19.730 ;
  RECT 2687.520 21.230 2688.660 22.070 ;
  RECT 2687.520 24.170 2688.660 25.170 ;
  RECT 2687.520 36.320 2688.660 37.320 ;
  RECT 2687.520 39.480 2688.660 40.080 ;
  RECT 2687.520 45.560 2688.660 46.160 ;
  RECT 2687.520 57.100 2688.660 61.420 ;
  RECT 4.280 57.100 5.420 61.420 ;
  RECT 4.280 45.560 5.420 46.160 ;
  RECT 4.280 39.480 5.420 40.080 ;
  RECT 4.280 36.320 5.420 37.320 ;
  RECT 4.280 24.170 5.420 25.170 ;
  RECT 4.280 21.230 5.420 22.070 ;
  RECT 4.280 18.730 5.420 19.730 ;
  RECT 4.280 14.200 5.420 15.200 ;
  RECT 4.280 9.570 5.420 11.170 ;
  RECT 2687.520 559.940 2688.660 560.320 ;
  RECT 2687.520 552.020 2688.660 552.300 ;
  RECT 2687.520 548.340 2688.660 548.620 ;
  RECT 2687.520 544.660 2688.660 544.940 ;
  RECT 2687.520 540.980 2688.660 541.260 ;
  RECT 2687.520 537.300 2688.660 537.580 ;
  RECT 2687.520 533.620 2688.660 533.900 ;
  RECT 2687.520 529.940 2688.660 530.220 ;
  RECT 2687.520 526.260 2688.660 526.540 ;
  RECT 2687.520 522.580 2688.660 522.860 ;
  RECT 2687.520 518.900 2688.660 519.180 ;
  RECT 2687.520 515.220 2688.660 515.500 ;
  RECT 2687.520 511.540 2688.660 511.820 ;
  RECT 2687.520 507.860 2688.660 508.140 ;
  RECT 2687.520 504.180 2688.660 504.460 ;
  RECT 2687.520 500.500 2688.660 500.780 ;
  RECT 2687.520 496.820 2688.660 497.100 ;
  RECT 2687.520 493.140 2688.660 493.420 ;
  RECT 2687.520 489.460 2688.660 489.740 ;
  RECT 2687.520 485.780 2688.660 486.060 ;
  RECT 2687.520 482.100 2688.660 482.380 ;
  RECT 2687.520 478.420 2688.660 478.700 ;
  RECT 2687.520 474.740 2688.660 475.020 ;
  RECT 2687.520 471.060 2688.660 471.340 ;
  RECT 2687.520 467.380 2688.660 467.660 ;
  RECT 2687.520 463.700 2688.660 463.980 ;
  RECT 2687.520 460.020 2688.660 460.300 ;
  RECT 2687.520 456.340 2688.660 456.620 ;
  RECT 2687.520 452.660 2688.660 452.940 ;
  RECT 2687.520 448.980 2688.660 449.260 ;
  RECT 2687.520 445.300 2688.660 445.580 ;
  RECT 2687.520 441.620 2688.660 441.900 ;
  RECT 2687.520 437.940 2688.660 438.220 ;
  RECT 2687.520 434.260 2688.660 434.540 ;
  RECT 2687.520 430.580 2688.660 430.860 ;
  RECT 2687.520 426.900 2688.660 427.180 ;
  RECT 2687.520 423.220 2688.660 423.500 ;
  RECT 2687.520 419.540 2688.660 419.820 ;
  RECT 2687.520 415.860 2688.660 416.140 ;
  RECT 2687.520 412.180 2688.660 412.460 ;
  RECT 2687.520 408.500 2688.660 408.780 ;
  RECT 2687.520 404.820 2688.660 405.100 ;
  RECT 2687.520 401.140 2688.660 401.420 ;
  RECT 2687.520 397.460 2688.660 397.740 ;
  RECT 2687.520 393.780 2688.660 394.060 ;
  RECT 2687.520 390.100 2688.660 390.380 ;
  RECT 2687.520 386.420 2688.660 386.700 ;
  RECT 2687.520 382.740 2688.660 383.020 ;
  RECT 2687.520 379.060 2688.660 379.340 ;
  RECT 2687.520 375.380 2688.660 375.660 ;
  RECT 2687.520 371.700 2688.660 371.980 ;
  RECT 2687.520 368.020 2688.660 368.300 ;
  RECT 2687.520 364.340 2688.660 364.620 ;
  RECT 2687.520 360.660 2688.660 360.940 ;
  RECT 2687.520 356.980 2688.660 357.260 ;
  RECT 2687.520 353.300 2688.660 353.580 ;
  RECT 2687.520 349.620 2688.660 349.900 ;
  RECT 2687.520 345.940 2688.660 346.220 ;
  RECT 2687.520 342.260 2688.660 342.540 ;
  RECT 2687.520 338.580 2688.660 338.860 ;
  RECT 2687.520 334.900 2688.660 335.180 ;
  RECT 2687.520 331.220 2688.660 331.500 ;
  RECT 2687.520 327.540 2688.660 327.820 ;
  RECT 2687.520 323.860 2688.660 324.140 ;
  RECT 2687.520 320.180 2688.660 320.460 ;
  RECT 2687.520 316.500 2688.660 316.780 ;
  RECT 2687.520 312.820 2688.660 313.100 ;
  RECT 2687.520 309.140 2688.660 309.420 ;
  RECT 2687.520 305.460 2688.660 305.740 ;
  RECT 2687.520 301.780 2688.660 302.060 ;
  RECT 2687.520 298.100 2688.660 298.380 ;
  RECT 2687.520 294.420 2688.660 294.700 ;
  RECT 2687.520 290.740 2688.660 291.020 ;
  RECT 2687.520 287.060 2688.660 287.340 ;
  RECT 2687.520 283.380 2688.660 283.660 ;
  RECT 2687.520 279.700 2688.660 279.980 ;
  RECT 2687.520 276.020 2688.660 276.300 ;
  RECT 2687.520 272.340 2688.660 272.620 ;
  RECT 2687.520 268.660 2688.660 268.940 ;
  RECT 2687.520 264.980 2688.660 265.260 ;
  RECT 2687.520 261.300 2688.660 261.580 ;
  RECT 2687.520 257.620 2688.660 257.900 ;
  RECT 2687.520 253.940 2688.660 254.220 ;
  RECT 2687.520 250.260 2688.660 250.540 ;
  RECT 2687.520 246.580 2688.660 246.860 ;
  RECT 2687.520 242.900 2688.660 243.180 ;
  RECT 2687.520 239.220 2688.660 239.500 ;
  RECT 2687.520 235.540 2688.660 235.820 ;
  RECT 2687.520 231.860 2688.660 232.140 ;
  RECT 2687.520 228.180 2688.660 228.460 ;
  RECT 2687.520 224.500 2688.660 224.780 ;
  RECT 2687.520 220.820 2688.660 221.100 ;
  RECT 2687.520 217.140 2688.660 217.420 ;
  RECT 2687.520 213.460 2688.660 213.740 ;
  RECT 2687.520 209.780 2688.660 210.060 ;
  RECT 2687.520 206.100 2688.660 206.380 ;
  RECT 2687.520 202.420 2688.660 202.700 ;
  RECT 2687.520 198.740 2688.660 199.020 ;
  RECT 2687.520 195.060 2688.660 195.340 ;
  RECT 2687.520 191.380 2688.660 191.660 ;
  RECT 2687.520 187.700 2688.660 187.980 ;
  RECT 2687.520 184.020 2688.660 184.300 ;
  RECT 2687.520 180.340 2688.660 180.620 ;
  RECT 2687.520 176.660 2688.660 176.940 ;
  RECT 2687.520 172.980 2688.660 173.260 ;
  RECT 2687.520 169.300 2688.660 169.580 ;
  RECT 2687.520 165.620 2688.660 165.900 ;
  RECT 2687.520 161.940 2688.660 162.220 ;
  RECT 2687.520 158.260 2688.660 158.540 ;
  RECT 2687.520 154.580 2688.660 154.860 ;
  RECT 2687.520 150.900 2688.660 151.180 ;
  RECT 2687.520 147.220 2688.660 147.500 ;
  RECT 2687.520 143.540 2688.660 143.820 ;
  RECT 2687.520 139.860 2688.660 140.140 ;
  RECT 2687.520 136.180 2688.660 136.460 ;
  RECT 2687.520 132.500 2688.660 132.780 ;
  RECT 2687.520 128.820 2688.660 129.100 ;
  RECT 2687.520 125.140 2688.660 125.420 ;
  RECT 2687.520 121.460 2688.660 121.740 ;
  RECT 2687.520 117.780 2688.660 118.060 ;
  RECT 2687.520 114.100 2688.660 114.380 ;
  RECT 2687.520 110.420 2688.660 110.700 ;
  RECT 2687.520 106.740 2688.660 107.020 ;
  RECT 2687.520 103.060 2688.660 103.340 ;
  RECT 2687.520 99.380 2688.660 99.660 ;
  RECT 2687.520 95.700 2688.660 95.980 ;
  RECT 2687.520 92.020 2688.660 92.300 ;
  RECT 2687.520 88.340 2688.660 88.620 ;
  RECT 2687.520 84.660 2688.660 84.940 ;
  RECT 2687.520 80.980 2688.660 81.260 ;
  RECT 2687.520 77.300 2688.660 77.580 ;
  RECT 2687.520 73.620 2688.660 73.900 ;
  RECT 2687.520 69.940 2688.660 70.220 ;
  RECT 2687.520 65.600 2688.660 65.980 ;
  RECT 1376.820 560.510 1377.070 561.650 ;
  RECT 1417.740 560.510 1417.990 561.650 ;
  RECT 1458.660 560.510 1458.910 561.650 ;
  RECT 1499.580 560.510 1499.830 561.650 ;
  RECT 1540.500 560.510 1540.750 561.650 ;
  RECT 1581.420 560.510 1581.670 561.650 ;
  RECT 1622.340 560.510 1622.590 561.650 ;
  RECT 1663.260 560.510 1663.510 561.650 ;
  RECT 1704.180 560.510 1704.430 561.650 ;
  RECT 1745.100 560.510 1745.350 561.650 ;
  RECT 1786.020 560.510 1786.270 561.650 ;
  RECT 1826.940 560.510 1827.190 561.650 ;
  RECT 1867.860 560.510 1868.110 561.650 ;
  RECT 1908.780 560.510 1909.030 561.650 ;
  RECT 1949.700 560.510 1949.950 561.650 ;
  RECT 1990.620 560.510 1990.870 561.650 ;
  RECT 2031.540 560.510 2031.790 561.650 ;
  RECT 2072.460 560.510 2072.710 561.650 ;
  RECT 2113.380 560.510 2113.630 561.650 ;
  RECT 2154.300 560.510 2154.550 561.650 ;
  RECT 2195.220 560.510 2195.470 561.650 ;
  RECT 2236.140 560.510 2236.390 561.650 ;
  RECT 2277.060 560.510 2277.310 561.650 ;
  RECT 2317.980 560.510 2318.230 561.650 ;
  RECT 2358.900 560.510 2359.150 561.650 ;
  RECT 2399.820 560.510 2400.070 561.650 ;
  RECT 2440.740 560.510 2440.990 561.650 ;
  RECT 2481.660 560.510 2481.910 561.650 ;
  RECT 2522.580 560.510 2522.830 561.650 ;
  RECT 2563.500 560.510 2563.750 561.650 ;
  RECT 2604.420 560.510 2604.670 561.650 ;
  RECT 2645.340 560.510 2645.590 561.650 ;
  RECT 1359.810 560.510 1362.320 561.650 ;
  RECT 1347.390 560.510 1349.780 561.650 ;
  RECT 1339.880 560.510 1342.940 561.650 ;
  RECT 1364.060 560.510 1366.910 561.650 ;
  RECT 1368.360 560.510 1371.610 561.650 ;
  RECT 1337.160 560.510 1338.920 561.650 ;
  RECT 1319.820 560.510 1321.580 561.650 ;
  RECT 1323.820 560.510 1325.580 561.650 ;
  RECT 1327.820 560.510 1329.580 561.650 ;
  RECT 1331.820 560.510 1333.580 561.650 ;
  RECT 4.280 65.600 5.420 65.980 ;
  RECT 4.280 69.940 5.420 70.220 ;
  RECT 4.280 73.620 5.420 73.900 ;
  RECT 4.280 77.300 5.420 77.580 ;
  RECT 4.280 80.980 5.420 81.260 ;
  RECT 4.280 84.660 5.420 84.940 ;
  RECT 4.280 88.340 5.420 88.620 ;
  RECT 4.280 92.020 5.420 92.300 ;
  RECT 4.280 95.700 5.420 95.980 ;
  RECT 4.280 99.380 5.420 99.660 ;
  RECT 4.280 103.060 5.420 103.340 ;
  RECT 4.280 106.740 5.420 107.020 ;
  RECT 4.280 110.420 5.420 110.700 ;
  RECT 4.280 114.100 5.420 114.380 ;
  RECT 4.280 117.780 5.420 118.060 ;
  RECT 4.280 121.460 5.420 121.740 ;
  RECT 4.280 125.140 5.420 125.420 ;
  RECT 4.280 128.820 5.420 129.100 ;
  RECT 4.280 132.500 5.420 132.780 ;
  RECT 4.280 136.180 5.420 136.460 ;
  RECT 4.280 139.860 5.420 140.140 ;
  RECT 4.280 143.540 5.420 143.820 ;
  RECT 4.280 147.220 5.420 147.500 ;
  RECT 4.280 150.900 5.420 151.180 ;
  RECT 4.280 154.580 5.420 154.860 ;
  RECT 4.280 158.260 5.420 158.540 ;
  RECT 4.280 161.940 5.420 162.220 ;
  RECT 4.280 165.620 5.420 165.900 ;
  RECT 4.280 169.300 5.420 169.580 ;
  RECT 4.280 172.980 5.420 173.260 ;
  RECT 4.280 176.660 5.420 176.940 ;
  RECT 4.280 180.340 5.420 180.620 ;
  RECT 4.280 184.020 5.420 184.300 ;
  RECT 4.280 187.700 5.420 187.980 ;
  RECT 4.280 191.380 5.420 191.660 ;
  RECT 4.280 195.060 5.420 195.340 ;
  RECT 4.280 198.740 5.420 199.020 ;
  RECT 4.280 202.420 5.420 202.700 ;
  RECT 4.280 206.100 5.420 206.380 ;
  RECT 4.280 209.780 5.420 210.060 ;
  RECT 4.280 213.460 5.420 213.740 ;
  RECT 4.280 217.140 5.420 217.420 ;
  RECT 4.280 220.820 5.420 221.100 ;
  RECT 4.280 224.500 5.420 224.780 ;
  RECT 4.280 228.180 5.420 228.460 ;
  RECT 4.280 231.860 5.420 232.140 ;
  RECT 4.280 235.540 5.420 235.820 ;
  RECT 4.280 239.220 5.420 239.500 ;
  RECT 4.280 242.900 5.420 243.180 ;
  RECT 4.280 246.580 5.420 246.860 ;
  RECT 4.280 250.260 5.420 250.540 ;
  RECT 4.280 253.940 5.420 254.220 ;
  RECT 4.280 257.620 5.420 257.900 ;
  RECT 4.280 261.300 5.420 261.580 ;
  RECT 4.280 264.980 5.420 265.260 ;
  RECT 4.280 268.660 5.420 268.940 ;
  RECT 4.280 272.340 5.420 272.620 ;
  RECT 4.280 276.020 5.420 276.300 ;
  RECT 4.280 279.700 5.420 279.980 ;
  RECT 4.280 283.380 5.420 283.660 ;
  RECT 4.280 287.060 5.420 287.340 ;
  RECT 4.280 290.740 5.420 291.020 ;
  RECT 4.280 294.420 5.420 294.700 ;
  RECT 4.280 298.100 5.420 298.380 ;
  RECT 4.280 301.780 5.420 302.060 ;
  RECT 4.280 305.460 5.420 305.740 ;
  RECT 4.280 309.140 5.420 309.420 ;
  RECT 4.280 312.820 5.420 313.100 ;
  RECT 4.280 316.500 5.420 316.780 ;
  RECT 4.280 320.180 5.420 320.460 ;
  RECT 4.280 323.860 5.420 324.140 ;
  RECT 4.280 327.540 5.420 327.820 ;
  RECT 4.280 331.220 5.420 331.500 ;
  RECT 4.280 334.900 5.420 335.180 ;
  RECT 4.280 338.580 5.420 338.860 ;
  RECT 4.280 342.260 5.420 342.540 ;
  RECT 4.280 345.940 5.420 346.220 ;
  RECT 4.280 349.620 5.420 349.900 ;
  RECT 4.280 353.300 5.420 353.580 ;
  RECT 4.280 356.980 5.420 357.260 ;
  RECT 4.280 360.660 5.420 360.940 ;
  RECT 4.280 364.340 5.420 364.620 ;
  RECT 4.280 368.020 5.420 368.300 ;
  RECT 4.280 371.700 5.420 371.980 ;
  RECT 4.280 375.380 5.420 375.660 ;
  RECT 4.280 379.060 5.420 379.340 ;
  RECT 4.280 382.740 5.420 383.020 ;
  RECT 4.280 386.420 5.420 386.700 ;
  RECT 4.280 390.100 5.420 390.380 ;
  RECT 4.280 393.780 5.420 394.060 ;
  RECT 4.280 397.460 5.420 397.740 ;
  RECT 4.280 401.140 5.420 401.420 ;
  RECT 4.280 404.820 5.420 405.100 ;
  RECT 4.280 408.500 5.420 408.780 ;
  RECT 4.280 412.180 5.420 412.460 ;
  RECT 4.280 415.860 5.420 416.140 ;
  RECT 4.280 419.540 5.420 419.820 ;
  RECT 4.280 423.220 5.420 423.500 ;
  RECT 4.280 426.900 5.420 427.180 ;
  RECT 4.280 430.580 5.420 430.860 ;
  RECT 4.280 434.260 5.420 434.540 ;
  RECT 4.280 437.940 5.420 438.220 ;
  RECT 4.280 441.620 5.420 441.900 ;
  RECT 4.280 445.300 5.420 445.580 ;
  RECT 4.280 448.980 5.420 449.260 ;
  RECT 4.280 452.660 5.420 452.940 ;
  RECT 4.280 456.340 5.420 456.620 ;
  RECT 4.280 460.020 5.420 460.300 ;
  RECT 4.280 463.700 5.420 463.980 ;
  RECT 4.280 467.380 5.420 467.660 ;
  RECT 4.280 471.060 5.420 471.340 ;
  RECT 4.280 474.740 5.420 475.020 ;
  RECT 4.280 478.420 5.420 478.700 ;
  RECT 4.280 482.100 5.420 482.380 ;
  RECT 4.280 485.780 5.420 486.060 ;
  RECT 4.280 489.460 5.420 489.740 ;
  RECT 4.280 493.140 5.420 493.420 ;
  RECT 4.280 496.820 5.420 497.100 ;
  RECT 4.280 500.500 5.420 500.780 ;
  RECT 4.280 504.180 5.420 504.460 ;
  RECT 4.280 507.860 5.420 508.140 ;
  RECT 4.280 511.540 5.420 511.820 ;
  RECT 4.280 515.220 5.420 515.500 ;
  RECT 4.280 518.900 5.420 519.180 ;
  RECT 4.280 522.580 5.420 522.860 ;
  RECT 4.280 526.260 5.420 526.540 ;
  RECT 4.280 529.940 5.420 530.220 ;
  RECT 4.280 533.620 5.420 533.900 ;
  RECT 4.280 537.300 5.420 537.580 ;
  RECT 4.280 540.980 5.420 541.260 ;
  RECT 4.280 544.660 5.420 544.940 ;
  RECT 4.280 548.340 5.420 548.620 ;
  RECT 4.280 552.020 5.420 552.300 ;
  RECT 4.280 559.940 5.420 560.320 ;
  RECT 47.350 560.510 47.600 561.650 ;
  RECT 88.270 560.510 88.520 561.650 ;
  RECT 129.190 560.510 129.440 561.650 ;
  RECT 170.110 560.510 170.360 561.650 ;
  RECT 211.030 560.510 211.280 561.650 ;
  RECT 251.950 560.510 252.200 561.650 ;
  RECT 292.870 560.510 293.120 561.650 ;
  RECT 333.790 560.510 334.040 561.650 ;
  RECT 374.710 560.510 374.960 561.650 ;
  RECT 415.630 560.510 415.880 561.650 ;
  RECT 456.550 560.510 456.800 561.650 ;
  RECT 497.470 560.510 497.720 561.650 ;
  RECT 538.390 560.510 538.640 561.650 ;
  RECT 579.310 560.510 579.560 561.650 ;
  RECT 620.230 560.510 620.480 561.650 ;
  RECT 661.150 560.510 661.400 561.650 ;
  RECT 702.070 560.510 702.320 561.650 ;
  RECT 742.990 560.510 743.240 561.650 ;
  RECT 783.910 560.510 784.160 561.650 ;
  RECT 824.830 560.510 825.080 561.650 ;
  RECT 865.750 560.510 866.000 561.650 ;
  RECT 906.670 560.510 906.920 561.650 ;
  RECT 947.590 560.510 947.840 561.650 ;
  RECT 988.510 560.510 988.760 561.650 ;
  RECT 1029.430 560.510 1029.680 561.650 ;
  RECT 1070.350 560.510 1070.600 561.650 ;
  RECT 1111.270 560.510 1111.520 561.650 ;
  RECT 1152.190 560.510 1152.440 561.650 ;
  RECT 1193.110 560.510 1193.360 561.650 ;
  RECT 1234.030 560.510 1234.280 561.650 ;
  RECT 1274.950 560.510 1275.200 561.650 ;
  LAYER ME1 ;
  RECT 5.420 7.020 2687.520 560.510 ;
  RECT 2691.080 3.460 2692.940 564.070 ;
  RECT 0.000 3.460 1.860 564.070 ;
  RECT 1.860 564.070 2691.080 565.930 ;
  RECT 1.860 1.600 2691.080 3.460 ;
  RECT 2688.940 5.600 2690.800 561.930 ;
  RECT 2.140 5.600 4.000 561.930 ;
  RECT 4.000 561.930 2688.940 563.790 ;
  RECT 4.000 3.740 2688.940 5.600 ;
  RECT 2.140 561.930 4.000 563.790 ;
  RECT 0.000 564.070 1.860 565.930 ;
  RECT 2688.940 3.740 2690.800 5.600 ;
  RECT 2691.080 1.600 2692.940 3.460 ;
  RECT 2688.940 561.930 2690.800 563.790 ;
  RECT 2691.080 564.070 2692.940 565.930 ;
  RECT 2.140 3.740 4.000 5.600 ;
  RECT 0.000 1.600 1.860 3.460 ;
  RECT 2680.800 0.000 2681.600 1.000 ;
  RECT 2666.400 0.000 2667.200 1.000 ;
  RECT 2661.200 0.000 2662.000 1.000 ;
  RECT 2646.400 0.000 2647.200 1.000 ;
  RECT 2640.000 0.000 2640.800 1.000 ;
  RECT 2625.600 0.000 2626.400 1.000 ;
  RECT 2620.400 0.000 2621.200 1.000 ;
  RECT 2605.600 0.000 2606.400 1.000 ;
  RECT 2599.200 0.000 2600.000 1.000 ;
  RECT 2584.400 0.000 2585.200 1.000 ;
  RECT 2579.200 0.000 2580.000 1.000 ;
  RECT 2564.800 0.000 2565.600 1.000 ;
  RECT 2558.400 0.000 2559.200 1.000 ;
  RECT 2543.600 0.000 2544.400 1.000 ;
  RECT 2538.400 0.000 2539.200 1.000 ;
  RECT 2525.600 0.000 2526.400 1.000 ;
  RECT 2523.600 0.000 2524.400 1.000 ;
  RECT 2517.200 0.000 2518.000 1.000 ;
  RECT 2502.800 0.000 2503.600 1.000 ;
  RECT 2497.600 0.000 2498.400 1.000 ;
  RECT 2482.800 0.000 2483.600 1.000 ;
  RECT 2476.400 0.000 2477.200 1.000 ;
  RECT 2461.600 0.000 2462.400 1.000 ;
  RECT 2456.400 0.000 2457.200 1.000 ;
  RECT 2442.000 0.000 2442.800 1.000 ;
  RECT 2435.600 0.000 2436.400 1.000 ;
  RECT 2420.800 0.000 2421.600 1.000 ;
  RECT 2415.600 0.000 2416.400 1.000 ;
  RECT 2400.800 0.000 2401.600 1.000 ;
  RECT 2394.400 0.000 2395.200 1.000 ;
  RECT 2380.000 0.000 2380.800 1.000 ;
  RECT 2374.800 0.000 2375.600 1.000 ;
  RECT 2361.600 0.000 2362.400 1.000 ;
  RECT 2360.000 0.000 2360.800 1.000 ;
  RECT 2353.600 0.000 2354.400 1.000 ;
  RECT 2338.800 0.000 2339.600 1.000 ;
  RECT 2333.600 0.000 2334.400 1.000 ;
  RECT 2319.200 0.000 2320.000 1.000 ;
  RECT 2312.800 0.000 2313.600 1.000 ;
  RECT 2298.000 0.000 2298.800 1.000 ;
  RECT 2292.800 0.000 2293.600 1.000 ;
  RECT 2278.400 0.000 2279.200 1.000 ;
  RECT 2271.600 0.000 2272.400 1.000 ;
  RECT 2257.200 0.000 2258.000 1.000 ;
  RECT 2252.000 0.000 2252.800 1.000 ;
  RECT 2237.200 0.000 2238.000 1.000 ;
  RECT 2230.800 0.000 2231.600 1.000 ;
  RECT 2216.400 0.000 2217.200 1.000 ;
  RECT 2211.200 0.000 2212.000 1.000 ;
  RECT 2198.000 0.000 2198.800 1.000 ;
  RECT 2196.400 0.000 2197.200 1.000 ;
  RECT 2190.000 0.000 2190.800 1.000 ;
  RECT 2175.200 0.000 2176.000 1.000 ;
  RECT 2170.000 0.000 2170.800 1.000 ;
  RECT 2155.600 0.000 2156.400 1.000 ;
  RECT 2149.200 0.000 2150.000 1.000 ;
  RECT 2134.400 0.000 2135.200 1.000 ;
  RECT 2129.200 0.000 2130.000 1.000 ;
  RECT 2114.400 0.000 2115.200 1.000 ;
  RECT 2108.000 0.000 2108.800 1.000 ;
  RECT 2093.600 0.000 2094.400 1.000 ;
  RECT 2088.400 0.000 2089.200 1.000 ;
  RECT 2073.600 0.000 2074.400 1.000 ;
  RECT 2067.200 0.000 2068.000 1.000 ;
  RECT 2052.400 0.000 2053.200 1.000 ;
  RECT 2047.200 0.000 2048.000 1.000 ;
  RECT 2034.400 0.000 2035.200 1.000 ;
  RECT 2032.800 0.000 2033.600 1.000 ;
  RECT 2026.400 0.000 2027.200 1.000 ;
  RECT 2011.600 0.000 2012.400 1.000 ;
  RECT 2006.400 0.000 2007.200 1.000 ;
  RECT 1991.600 0.000 1992.400 1.000 ;
  RECT 1985.200 0.000 1986.000 1.000 ;
  RECT 1970.800 0.000 1971.600 1.000 ;
  RECT 1965.600 0.000 1966.400 1.000 ;
  RECT 1950.800 0.000 1951.600 1.000 ;
  RECT 1944.400 0.000 1945.200 1.000 ;
  RECT 1929.600 0.000 1930.400 1.000 ;
  RECT 1924.400 0.000 1925.200 1.000 ;
  RECT 1910.000 0.000 1910.800 1.000 ;
  RECT 1903.600 0.000 1904.400 1.000 ;
  RECT 1888.800 0.000 1889.600 1.000 ;
  RECT 1883.600 0.000 1884.400 1.000 ;
  RECT 1870.800 0.000 1871.600 1.000 ;
  RECT 1869.200 0.000 1870.000 1.000 ;
  RECT 1862.400 0.000 1863.200 1.000 ;
  RECT 1848.000 0.000 1848.800 1.000 ;
  RECT 1842.800 0.000 1843.600 1.000 ;
  RECT 1828.000 0.000 1828.800 1.000 ;
  RECT 1821.600 0.000 1822.400 1.000 ;
  RECT 1807.200 0.000 1808.000 1.000 ;
  RECT 1802.000 0.000 1802.800 1.000 ;
  RECT 1787.200 0.000 1788.000 1.000 ;
  RECT 1780.800 0.000 1781.600 1.000 ;
  RECT 1766.000 0.000 1766.800 1.000 ;
  RECT 1760.800 0.000 1761.600 1.000 ;
  RECT 1746.400 0.000 1747.200 1.000 ;
  RECT 1740.000 0.000 1740.800 1.000 ;
  RECT 1725.200 0.000 1726.000 1.000 ;
  RECT 1720.000 0.000 1720.800 1.000 ;
  RECT 1707.200 0.000 1708.000 1.000 ;
  RECT 1705.200 0.000 1706.000 1.000 ;
  RECT 1698.800 0.000 1699.600 1.000 ;
  RECT 1684.400 0.000 1685.200 1.000 ;
  RECT 1679.200 0.000 1680.000 1.000 ;
  RECT 1664.400 0.000 1665.200 1.000 ;
  RECT 1658.000 0.000 1658.800 1.000 ;
  RECT 1643.200 0.000 1644.000 1.000 ;
  RECT 1638.000 0.000 1638.800 1.000 ;
  RECT 1623.600 0.000 1624.400 1.000 ;
  RECT 1617.200 0.000 1618.000 1.000 ;
  RECT 1602.400 0.000 1603.200 1.000 ;
  RECT 1597.200 0.000 1598.000 1.000 ;
  RECT 1582.400 0.000 1583.200 1.000 ;
  RECT 1576.000 0.000 1576.800 1.000 ;
  RECT 1561.600 0.000 1562.400 1.000 ;
  RECT 1556.400 0.000 1557.200 1.000 ;
  RECT 1543.200 0.000 1544.000 1.000 ;
  RECT 1541.600 0.000 1542.400 1.000 ;
  RECT 1535.200 0.000 1536.000 1.000 ;
  RECT 1520.400 0.000 1521.200 1.000 ;
  RECT 1515.200 0.000 1516.000 1.000 ;
  RECT 1500.800 0.000 1501.600 1.000 ;
  RECT 1494.400 0.000 1495.200 1.000 ;
  RECT 1479.600 0.000 1480.400 1.000 ;
  RECT 1474.400 0.000 1475.200 1.000 ;
  RECT 1460.000 0.000 1460.800 1.000 ;
  RECT 1453.200 0.000 1454.000 1.000 ;
  RECT 1438.800 0.000 1439.600 1.000 ;
  RECT 1433.600 0.000 1434.400 1.000 ;
  RECT 1418.800 0.000 1419.600 1.000 ;
  RECT 1412.400 0.000 1413.200 1.000 ;
  RECT 1398.000 0.000 1398.800 1.000 ;
  RECT 1392.800 0.000 1393.600 1.000 ;
  RECT 1379.600 0.000 1380.400 1.000 ;
  RECT 1378.000 0.000 1378.800 1.000 ;
  RECT 1357.200 0.000 1358.000 1.000 ;
  RECT 1356.000 0.000 1356.800 1.000 ;
  RECT 1354.800 0.000 1355.600 1.000 ;
  RECT 1353.600 0.000 1354.400 1.000 ;
  RECT 1352.400 0.000 1353.200 1.000 ;
  RECT 1351.200 0.000 1352.000 1.000 ;
  RECT 1345.200 0.000 1346.000 1.000 ;
  RECT 1338.000 0.000 1338.800 1.000 ;
  RECT 1335.200 0.000 1336.000 1.000 ;
  RECT 1332.400 0.000 1333.200 1.000 ;
  RECT 1330.000 0.000 1330.800 1.000 ;
  RECT 1328.400 0.000 1329.200 1.000 ;
  RECT 1326.000 0.000 1326.800 1.000 ;
  RECT 1324.400 0.000 1325.200 1.000 ;
  RECT 1322.000 0.000 1322.800 1.000 ;
  RECT 1320.400 0.000 1321.200 1.000 ;
  RECT 1311.200 0.000 1312.000 1.000 ;
  RECT 1296.400 0.000 1297.200 1.000 ;
  RECT 1291.200 0.000 1292.000 1.000 ;
  RECT 1276.800 0.000 1277.600 1.000 ;
  RECT 1270.400 0.000 1271.200 1.000 ;
  RECT 1255.600 0.000 1256.400 1.000 ;
  RECT 1250.400 0.000 1251.200 1.000 ;
  RECT 1235.600 0.000 1236.400 1.000 ;
  RECT 1229.200 0.000 1230.000 1.000 ;
  RECT 1214.800 0.000 1215.600 1.000 ;
  RECT 1209.600 0.000 1210.400 1.000 ;
  RECT 1194.800 0.000 1195.600 1.000 ;
  RECT 1188.400 0.000 1189.200 1.000 ;
  RECT 1173.600 0.000 1174.400 1.000 ;
  RECT 1168.400 0.000 1169.200 1.000 ;
  RECT 1155.600 0.000 1156.400 1.000 ;
  RECT 1154.000 0.000 1154.800 1.000 ;
  RECT 1147.600 0.000 1148.400 1.000 ;
  RECT 1132.800 0.000 1133.600 1.000 ;
  RECT 1127.600 0.000 1128.400 1.000 ;
  RECT 1113.200 0.000 1114.000 1.000 ;
  RECT 1106.400 0.000 1107.200 1.000 ;
  RECT 1092.000 0.000 1092.800 1.000 ;
  RECT 1086.800 0.000 1087.600 1.000 ;
  RECT 1072.000 0.000 1072.800 1.000 ;
  RECT 1065.600 0.000 1066.400 1.000 ;
  RECT 1051.200 0.000 1052.000 1.000 ;
  RECT 1045.600 0.000 1046.400 1.000 ;
  RECT 1031.200 0.000 1032.000 1.000 ;
  RECT 1024.800 0.000 1025.600 1.000 ;
  RECT 1010.000 0.000 1010.800 1.000 ;
  RECT 1004.800 0.000 1005.600 1.000 ;
  RECT 992.000 0.000 992.800 1.000 ;
  RECT 990.400 0.000 991.200 1.000 ;
  RECT 983.600 0.000 984.400 1.000 ;
  RECT 969.200 0.000 970.000 1.000 ;
  RECT 964.000 0.000 964.800 1.000 ;
  RECT 949.200 0.000 950.000 1.000 ;
  RECT 942.800 0.000 943.600 1.000 ;
  RECT 928.400 0.000 929.200 1.000 ;
  RECT 923.200 0.000 924.000 1.000 ;
  RECT 908.400 0.000 909.200 1.000 ;
  RECT 902.000 0.000 902.800 1.000 ;
  RECT 887.200 0.000 888.000 1.000 ;
  RECT 882.000 0.000 882.800 1.000 ;
  RECT 867.600 0.000 868.400 1.000 ;
  RECT 861.200 0.000 862.000 1.000 ;
  RECT 846.400 0.000 847.200 1.000 ;
  RECT 841.200 0.000 842.000 1.000 ;
  RECT 828.400 0.000 829.200 1.000 ;
  RECT 826.400 0.000 827.200 1.000 ;
  RECT 820.000 0.000 820.800 1.000 ;
  RECT 805.600 0.000 806.400 1.000 ;
  RECT 800.400 0.000 801.200 1.000 ;
  RECT 785.600 0.000 786.400 1.000 ;
  RECT 779.200 0.000 780.000 1.000 ;
  RECT 764.400 0.000 765.200 1.000 ;
  RECT 759.200 0.000 760.000 1.000 ;
  RECT 744.800 0.000 745.600 1.000 ;
  RECT 738.400 0.000 739.200 1.000 ;
  RECT 723.600 0.000 724.400 1.000 ;
  RECT 718.400 0.000 719.200 1.000 ;
  RECT 704.000 0.000 704.800 1.000 ;
  RECT 697.200 0.000 698.000 1.000 ;
  RECT 682.800 0.000 683.600 1.000 ;
  RECT 677.600 0.000 678.400 1.000 ;
  RECT 664.800 0.000 665.600 1.000 ;
  RECT 662.800 0.000 663.600 1.000 ;
  RECT 656.400 0.000 657.200 1.000 ;
  RECT 642.000 0.000 642.800 1.000 ;
  RECT 636.400 0.000 637.200 1.000 ;
  RECT 622.000 0.000 622.800 1.000 ;
  RECT 615.600 0.000 616.400 1.000 ;
  RECT 600.800 0.000 601.600 1.000 ;
  RECT 595.600 0.000 596.400 1.000 ;
  RECT 581.200 0.000 582.000 1.000 ;
  RECT 574.400 0.000 575.200 1.000 ;
  RECT 560.000 0.000 560.800 1.000 ;
  RECT 554.800 0.000 555.600 1.000 ;
  RECT 540.000 0.000 540.800 1.000 ;
  RECT 533.600 0.000 534.400 1.000 ;
  RECT 519.200 0.000 520.000 1.000 ;
  RECT 514.000 0.000 514.800 1.000 ;
  RECT 500.800 0.000 501.600 1.000 ;
  RECT 499.200 0.000 500.000 1.000 ;
  RECT 492.800 0.000 493.600 1.000 ;
  RECT 478.000 0.000 478.800 1.000 ;
  RECT 472.800 0.000 473.600 1.000 ;
  RECT 458.400 0.000 459.200 1.000 ;
  RECT 452.000 0.000 452.800 1.000 ;
  RECT 437.200 0.000 438.000 1.000 ;
  RECT 432.000 0.000 432.800 1.000 ;
  RECT 417.200 0.000 418.000 1.000 ;
  RECT 410.800 0.000 411.600 1.000 ;
  RECT 396.400 0.000 397.200 1.000 ;
  RECT 391.200 0.000 392.000 1.000 ;
  RECT 376.400 0.000 377.200 1.000 ;
  RECT 370.000 0.000 370.800 1.000 ;
  RECT 355.200 0.000 356.000 1.000 ;
  RECT 350.000 0.000 350.800 1.000 ;
  RECT 337.200 0.000 338.000 1.000 ;
  RECT 335.600 0.000 336.400 1.000 ;
  RECT 329.200 0.000 330.000 1.000 ;
  RECT 314.400 0.000 315.200 1.000 ;
  RECT 309.200 0.000 310.000 1.000 ;
  RECT 294.800 0.000 295.600 1.000 ;
  RECT 288.000 0.000 288.800 1.000 ;
  RECT 273.600 0.000 274.400 1.000 ;
  RECT 268.400 0.000 269.200 1.000 ;
  RECT 253.600 0.000 254.400 1.000 ;
  RECT 247.200 0.000 248.000 1.000 ;
  RECT 232.800 0.000 233.600 1.000 ;
  RECT 227.200 0.000 228.000 1.000 ;
  RECT 212.800 0.000 213.600 1.000 ;
  RECT 206.400 0.000 207.200 1.000 ;
  RECT 191.600 0.000 192.400 1.000 ;
  RECT 186.400 0.000 187.200 1.000 ;
  RECT 173.600 0.000 174.400 1.000 ;
  RECT 172.000 0.000 172.800 1.000 ;
  RECT 165.200 0.000 166.000 1.000 ;
  RECT 150.800 0.000 151.600 1.000 ;
  RECT 145.600 0.000 146.400 1.000 ;
  RECT 130.800 0.000 131.600 1.000 ;
  RECT 124.400 0.000 125.200 1.000 ;
  RECT 110.000 0.000 110.800 1.000 ;
  RECT 104.800 0.000 105.600 1.000 ;
  RECT 90.000 0.000 90.800 1.000 ;
  RECT 83.600 0.000 84.400 1.000 ;
  RECT 68.800 0.000 69.600 1.000 ;
  RECT 63.600 0.000 64.400 1.000 ;
  RECT 49.200 0.000 50.000 1.000 ;
  RECT 42.800 0.000 43.600 1.000 ;
  RECT 28.000 0.000 28.800 1.000 ;
  RECT 22.800 0.000 23.600 1.000 ;
  RECT 10.000 0.000 10.800 1.000 ;
  RECT 8.000 0.000 8.800 1.000 ;
  LAYER VI2 ;
  RECT 2691.080 3.600 2692.940 563.930 ;
  LAYER VI1 ;
  RECT 2691.080 3.460 2692.940 564.070 ;
  LAYER VI2 ;
  RECT 0.000 3.600 1.860 563.930 ;
  LAYER VI1 ;
  RECT 0.000 3.460 1.860 564.070 ;
  LAYER VI2 ;
  RECT 2.000 564.070 2690.940 565.930 ;
  LAYER VI1 ;
  RECT 1.860 564.070 2691.080 565.930 ;
  LAYER VI2 ;
  RECT 2682.600 1.600 2690.940 3.460 ;
  LAYER VI2 ;
  RECT 2668.200 1.600 2680.280 3.460 ;
  LAYER VI2 ;
  RECT 2663.000 1.600 2665.650 3.460 ;
  LAYER VI2 ;
  RECT 2648.200 1.600 2660.440 3.460 ;
  LAYER VI2 ;
  RECT 2641.800 1.600 2645.810 3.460 ;
  LAYER VI2 ;
  RECT 2627.400 1.600 2639.360 3.460 ;
  LAYER VI2 ;
  RECT 2622.200 1.600 2624.730 3.460 ;
  LAYER VI2 ;
  RECT 2607.400 1.600 2619.520 3.460 ;
  LAYER VI2 ;
  RECT 2601.000 1.600 2604.890 3.460 ;
  LAYER VI2 ;
  RECT 2586.200 1.600 2598.440 3.460 ;
  LAYER VI2 ;
  RECT 2581.000 1.600 2583.810 3.460 ;
  LAYER VI2 ;
  RECT 2566.600 1.600 2578.600 3.460 ;
  LAYER VI2 ;
  RECT 2560.200 1.600 2563.970 3.460 ;
  LAYER VI2 ;
  RECT 2545.400 1.600 2557.520 3.460 ;
  LAYER VI2 ;
  RECT 2540.200 1.600 2542.890 3.460 ;
  LAYER VI2 ;
  RECT 2527.400 1.600 2537.680 3.460 ;
  LAYER VI2 ;
  RECT 2519.000 1.600 2523.050 3.460 ;
  LAYER VI2 ;
  RECT 2504.600 1.600 2516.600 3.460 ;
  LAYER VI2 ;
  RECT 2499.400 1.600 2501.970 3.460 ;
  LAYER VI2 ;
  RECT 2484.600 1.600 2496.760 3.460 ;
  LAYER VI2 ;
  RECT 2478.200 1.600 2482.130 3.460 ;
  LAYER VI2 ;
  RECT 2463.400 1.600 2475.680 3.460 ;
  LAYER VI2 ;
  RECT 2458.200 1.600 2461.050 3.460 ;
  LAYER VI2 ;
  RECT 2443.800 1.600 2455.840 3.460 ;
  LAYER VI2 ;
  RECT 2437.400 1.600 2441.210 3.460 ;
  LAYER VI2 ;
  RECT 2422.600 1.600 2434.760 3.460 ;
  LAYER VI2 ;
  RECT 2417.400 1.600 2420.130 3.460 ;
  LAYER VI2 ;
  RECT 2402.600 1.600 2414.920 3.460 ;
  LAYER VI2 ;
  RECT 2396.200 1.600 2400.290 3.460 ;
  LAYER VI2 ;
  RECT 2381.800 1.600 2393.840 3.460 ;
  LAYER VI2 ;
  RECT 2376.600 1.600 2379.210 3.460 ;
  LAYER VI2 ;
  RECT 2363.400 1.600 2374.000 3.460 ;
  LAYER VI2 ;
  RECT 2355.400 1.600 2359.370 3.460 ;
  LAYER VI2 ;
  RECT 2340.600 1.600 2352.920 3.460 ;
  LAYER VI2 ;
  RECT 2335.400 1.600 2338.290 3.460 ;
  LAYER VI2 ;
  RECT 2321.000 1.600 2333.080 3.460 ;
  LAYER VI2 ;
  RECT 2314.600 1.600 2318.450 3.460 ;
  LAYER VI2 ;
  RECT 2299.800 1.600 2312.000 3.460 ;
  LAYER VI2 ;
  RECT 2294.600 1.600 2297.370 3.460 ;
  LAYER VI2 ;
  RECT 2280.200 1.600 2292.160 3.460 ;
  LAYER VI2 ;
  RECT 2273.400 1.600 2277.530 3.460 ;
  LAYER VI2 ;
  RECT 2259.000 1.600 2271.080 3.460 ;
  LAYER VI2 ;
  RECT 2253.800 1.600 2256.450 3.460 ;
  LAYER VI2 ;
  RECT 2239.000 1.600 2251.240 3.460 ;
  LAYER VI2 ;
  RECT 2232.600 1.600 2236.610 3.460 ;
  LAYER VI2 ;
  RECT 2218.200 1.600 2230.160 3.460 ;
  LAYER VI2 ;
  RECT 2213.000 1.600 2215.530 3.460 ;
  LAYER VI2 ;
  RECT 2199.800 1.600 2210.320 3.460 ;
  LAYER VI2 ;
  RECT 2191.800 1.600 2195.690 3.460 ;
  LAYER VI2 ;
  RECT 2177.000 1.600 2189.240 3.460 ;
  LAYER VI2 ;
  RECT 2171.800 1.600 2174.610 3.460 ;
  LAYER VI2 ;
  RECT 2157.400 1.600 2169.400 3.460 ;
  LAYER VI2 ;
  RECT 2151.000 1.600 2154.770 3.460 ;
  LAYER VI2 ;
  RECT 2136.200 1.600 2148.320 3.460 ;
  LAYER VI2 ;
  RECT 2131.000 1.600 2133.690 3.460 ;
  LAYER VI2 ;
  RECT 2116.200 1.600 2128.480 3.460 ;
  LAYER VI2 ;
  RECT 2109.800 1.600 2113.850 3.460 ;
  LAYER VI2 ;
  RECT 2095.400 1.600 2107.400 3.460 ;
  LAYER VI2 ;
  RECT 2090.200 1.600 2092.770 3.460 ;
  LAYER VI2 ;
  RECT 2075.400 1.600 2087.560 3.460 ;
  LAYER VI2 ;
  RECT 2069.000 1.600 2072.930 3.460 ;
  LAYER VI2 ;
  RECT 2054.200 1.600 2066.480 3.460 ;
  LAYER VI2 ;
  RECT 2049.000 1.600 2051.850 3.460 ;
  LAYER VI2 ;
  RECT 2036.200 1.600 2046.640 3.460 ;
  LAYER VI2 ;
  RECT 2028.200 1.600 2032.010 3.460 ;
  LAYER VI2 ;
  RECT 2013.400 1.600 2025.560 3.460 ;
  LAYER VI2 ;
  RECT 2008.200 1.600 2010.930 3.460 ;
  LAYER VI2 ;
  RECT 1993.400 1.600 2005.720 3.460 ;
  LAYER VI2 ;
  RECT 1987.000 1.600 1991.090 3.460 ;
  LAYER VI2 ;
  RECT 1972.600 1.600 1984.640 3.460 ;
  LAYER VI2 ;
  RECT 1967.400 1.600 1970.010 3.460 ;
  LAYER VI2 ;
  RECT 1952.600 1.600 1964.800 3.460 ;
  LAYER VI2 ;
  RECT 1946.200 1.600 1950.170 3.460 ;
  LAYER VI2 ;
  RECT 1931.400 1.600 1943.720 3.460 ;
  LAYER VI2 ;
  RECT 1926.200 1.600 1929.090 3.460 ;
  LAYER VI2 ;
  RECT 1911.800 1.600 1923.880 3.460 ;
  LAYER VI2 ;
  RECT 1905.400 1.600 1909.250 3.460 ;
  LAYER VI2 ;
  RECT 1890.600 1.600 1902.800 3.460 ;
  LAYER VI2 ;
  RECT 1885.400 1.600 1888.170 3.460 ;
  LAYER VI2 ;
  RECT 1872.600 1.600 1882.960 3.460 ;
  LAYER VI2 ;
  RECT 1864.200 1.600 1868.330 3.460 ;
  LAYER VI2 ;
  RECT 1849.800 1.600 1861.880 3.460 ;
  LAYER VI2 ;
  RECT 1844.600 1.600 1847.250 3.460 ;
  LAYER VI2 ;
  RECT 1829.800 1.600 1842.040 3.460 ;
  LAYER VI2 ;
  RECT 1823.400 1.600 1827.410 3.460 ;
  LAYER VI2 ;
  RECT 1809.000 1.600 1820.960 3.460 ;
  LAYER VI2 ;
  RECT 1803.800 1.600 1806.330 3.460 ;
  LAYER VI2 ;
  RECT 1789.000 1.600 1801.120 3.460 ;
  LAYER VI2 ;
  RECT 1782.600 1.600 1786.490 3.460 ;
  LAYER VI2 ;
  RECT 1767.800 1.600 1780.040 3.460 ;
  LAYER VI2 ;
  RECT 1762.600 1.600 1765.410 3.460 ;
  LAYER VI2 ;
  RECT 1748.200 1.600 1760.200 3.460 ;
  LAYER VI2 ;
  RECT 1741.800 1.600 1745.570 3.460 ;
  LAYER VI2 ;
  RECT 1727.000 1.600 1739.120 3.460 ;
  LAYER VI2 ;
  RECT 1721.800 1.600 1724.490 3.460 ;
  LAYER VI2 ;
  RECT 1709.000 1.600 1719.280 3.460 ;
  LAYER VI2 ;
  RECT 1700.600 1.600 1704.650 3.460 ;
  LAYER VI2 ;
  RECT 1686.200 1.600 1698.200 3.460 ;
  LAYER VI2 ;
  RECT 1681.000 1.600 1683.570 3.460 ;
  LAYER VI2 ;
  RECT 1666.200 1.600 1678.360 3.460 ;
  LAYER VI2 ;
  RECT 1659.800 1.600 1663.730 3.460 ;
  LAYER VI2 ;
  RECT 1645.000 1.600 1657.280 3.460 ;
  LAYER VI2 ;
  RECT 1639.800 1.600 1642.650 3.460 ;
  LAYER VI2 ;
  RECT 1625.400 1.600 1637.440 3.460 ;
  LAYER VI2 ;
  RECT 1619.000 1.600 1622.810 3.460 ;
  LAYER VI2 ;
  RECT 1604.200 1.600 1616.360 3.460 ;
  LAYER VI2 ;
  RECT 1599.000 1.600 1601.730 3.460 ;
  LAYER VI2 ;
  RECT 1584.200 1.600 1596.520 3.460 ;
  LAYER VI2 ;
  RECT 1577.800 1.600 1581.890 3.460 ;
  LAYER VI2 ;
  RECT 1563.400 1.600 1575.440 3.460 ;
  LAYER VI2 ;
  RECT 1558.200 1.600 1560.810 3.460 ;
  LAYER VI2 ;
  RECT 1545.000 1.600 1555.600 3.460 ;
  LAYER VI2 ;
  RECT 1537.000 1.600 1540.970 3.460 ;
  LAYER VI2 ;
  RECT 1522.200 1.600 1534.520 3.460 ;
  LAYER VI2 ;
  RECT 1517.000 1.600 1519.890 3.460 ;
  LAYER VI2 ;
  RECT 1502.600 1.600 1514.680 3.460 ;
  LAYER VI2 ;
  RECT 1496.200 1.600 1500.050 3.460 ;
  LAYER VI2 ;
  RECT 1481.400 1.600 1493.600 3.460 ;
  LAYER VI2 ;
  RECT 1476.200 1.600 1478.970 3.460 ;
  LAYER VI2 ;
  RECT 1461.800 1.600 1473.760 3.460 ;
  LAYER VI2 ;
  RECT 1455.000 1.600 1459.130 3.460 ;
  LAYER VI2 ;
  RECT 1440.600 1.600 1452.680 3.460 ;
  LAYER VI2 ;
  RECT 1435.400 1.600 1438.050 3.460 ;
  LAYER VI2 ;
  RECT 1420.600 1.600 1432.840 3.460 ;
  LAYER VI2 ;
  RECT 1414.200 1.600 1418.210 3.460 ;
  LAYER VI2 ;
  RECT 1399.800 1.600 1411.760 3.460 ;
  LAYER VI2 ;
  RECT 1394.600 1.600 1397.130 3.460 ;
  LAYER VI2 ;
  RECT 1381.400 1.600 1391.920 3.460 ;
  LAYER VI2 ;
  RECT 1359.000 1.600 1377.290 3.460 ;
  LAYER VI2 ;
  RECT 1347.000 1.600 1350.450 3.460 ;
  LAYER VI2 ;
  RECT 1339.800 1.600 1344.480 3.460 ;
  LAYER VI2 ;
  RECT 1313.000 1.600 1319.840 3.460 ;
  LAYER VI2 ;
  RECT 1298.200 1.600 1310.460 3.460 ;
  LAYER VI2 ;
  RECT 1293.000 1.600 1295.830 3.460 ;
  LAYER VI2 ;
  RECT 1278.600 1.600 1290.620 3.460 ;
  LAYER VI2 ;
  RECT 1272.200 1.600 1275.990 3.460 ;
  LAYER VI2 ;
  RECT 1257.400 1.600 1269.540 3.460 ;
  LAYER VI2 ;
  RECT 1252.200 1.600 1254.910 3.460 ;
  LAYER VI2 ;
  RECT 1237.400 1.600 1249.700 3.460 ;
  LAYER VI2 ;
  RECT 1231.000 1.600 1235.070 3.460 ;
  LAYER VI2 ;
  RECT 1216.600 1.600 1228.620 3.460 ;
  LAYER VI2 ;
  RECT 1211.400 1.600 1213.990 3.460 ;
  LAYER VI2 ;
  RECT 1196.600 1.600 1208.780 3.460 ;
  LAYER VI2 ;
  RECT 1190.200 1.600 1194.150 3.460 ;
  LAYER VI2 ;
  RECT 1175.400 1.600 1187.700 3.460 ;
  LAYER VI2 ;
  RECT 1170.200 1.600 1173.070 3.460 ;
  LAYER VI2 ;
  RECT 1157.400 1.600 1167.860 3.460 ;
  LAYER VI2 ;
  RECT 1149.400 1.600 1153.230 3.460 ;
  LAYER VI2 ;
  RECT 1134.600 1.600 1146.780 3.460 ;
  LAYER VI2 ;
  RECT 1129.400 1.600 1132.150 3.460 ;
  LAYER VI2 ;
  RECT 1115.000 1.600 1126.940 3.460 ;
  LAYER VI2 ;
  RECT 1108.200 1.600 1112.310 3.460 ;
  LAYER VI2 ;
  RECT 1093.800 1.600 1105.860 3.460 ;
  LAYER VI2 ;
  RECT 1088.600 1.600 1091.230 3.460 ;
  LAYER VI2 ;
  RECT 1073.800 1.600 1086.020 3.460 ;
  LAYER VI2 ;
  RECT 1067.400 1.600 1071.390 3.460 ;
  LAYER VI2 ;
  RECT 1053.000 1.600 1064.940 3.460 ;
  LAYER VI2 ;
  RECT 1047.400 1.600 1050.310 3.460 ;
  LAYER VI2 ;
  RECT 1033.000 1.600 1045.100 3.460 ;
  LAYER VI2 ;
  RECT 1026.600 1.600 1030.470 3.460 ;
  LAYER VI2 ;
  RECT 1011.800 1.600 1024.020 3.460 ;
  LAYER VI2 ;
  RECT 1006.600 1.600 1009.390 3.460 ;
  LAYER VI2 ;
  RECT 993.800 1.600 1004.180 3.460 ;
  LAYER VI2 ;
  RECT 985.400 1.600 989.550 3.460 ;
  LAYER VI2 ;
  RECT 971.000 1.600 983.100 3.460 ;
  LAYER VI2 ;
  RECT 965.800 1.600 968.470 3.460 ;
  LAYER VI2 ;
  RECT 951.000 1.600 963.260 3.460 ;
  LAYER VI2 ;
  RECT 944.600 1.600 948.630 3.460 ;
  LAYER VI2 ;
  RECT 930.200 1.600 942.180 3.460 ;
  LAYER VI2 ;
  RECT 925.000 1.600 927.550 3.460 ;
  LAYER VI2 ;
  RECT 910.200 1.600 922.340 3.460 ;
  LAYER VI2 ;
  RECT 903.800 1.600 907.710 3.460 ;
  LAYER VI2 ;
  RECT 889.000 1.600 901.260 3.460 ;
  LAYER VI2 ;
  RECT 883.800 1.600 886.630 3.460 ;
  LAYER VI2 ;
  RECT 869.400 1.600 881.420 3.460 ;
  LAYER VI2 ;
  RECT 863.000 1.600 866.790 3.460 ;
  LAYER VI2 ;
  RECT 848.200 1.600 860.340 3.460 ;
  LAYER VI2 ;
  RECT 843.000 1.600 845.710 3.460 ;
  LAYER VI2 ;
  RECT 830.200 1.600 840.500 3.460 ;
  LAYER VI2 ;
  RECT 821.800 1.600 825.870 3.460 ;
  LAYER VI2 ;
  RECT 807.400 1.600 819.420 3.460 ;
  LAYER VI2 ;
  RECT 802.200 1.600 804.790 3.460 ;
  LAYER VI2 ;
  RECT 787.400 1.600 799.580 3.460 ;
  LAYER VI2 ;
  RECT 781.000 1.600 784.950 3.460 ;
  LAYER VI2 ;
  RECT 766.200 1.600 778.500 3.460 ;
  LAYER VI2 ;
  RECT 761.000 1.600 763.870 3.460 ;
  LAYER VI2 ;
  RECT 746.600 1.600 758.660 3.460 ;
  LAYER VI2 ;
  RECT 740.200 1.600 744.030 3.460 ;
  LAYER VI2 ;
  RECT 725.400 1.600 737.580 3.460 ;
  LAYER VI2 ;
  RECT 720.200 1.600 722.950 3.460 ;
  LAYER VI2 ;
  RECT 705.800 1.600 717.740 3.460 ;
  LAYER VI2 ;
  RECT 699.000 1.600 703.110 3.460 ;
  LAYER VI2 ;
  RECT 684.600 1.600 696.660 3.460 ;
  LAYER VI2 ;
  RECT 679.400 1.600 682.030 3.460 ;
  LAYER VI2 ;
  RECT 666.600 1.600 676.820 3.460 ;
  LAYER VI2 ;
  RECT 658.200 1.600 662.190 3.460 ;
  LAYER VI2 ;
  RECT 643.800 1.600 655.740 3.460 ;
  LAYER VI2 ;
  RECT 638.200 1.600 641.110 3.460 ;
  LAYER VI2 ;
  RECT 623.800 1.600 635.900 3.460 ;
  LAYER VI2 ;
  RECT 617.400 1.600 621.270 3.460 ;
  LAYER VI2 ;
  RECT 602.600 1.600 614.820 3.460 ;
  LAYER VI2 ;
  RECT 597.400 1.600 600.190 3.460 ;
  LAYER VI2 ;
  RECT 583.000 1.600 594.980 3.460 ;
  LAYER VI2 ;
  RECT 576.200 1.600 580.350 3.460 ;
  LAYER VI2 ;
  RECT 561.800 1.600 573.900 3.460 ;
  LAYER VI2 ;
  RECT 556.600 1.600 559.270 3.460 ;
  LAYER VI2 ;
  RECT 541.800 1.600 554.060 3.460 ;
  LAYER VI2 ;
  RECT 535.400 1.600 539.430 3.460 ;
  LAYER VI2 ;
  RECT 521.000 1.600 532.980 3.460 ;
  LAYER VI2 ;
  RECT 515.800 1.600 518.350 3.460 ;
  LAYER VI2 ;
  RECT 502.600 1.600 513.140 3.460 ;
  LAYER VI2 ;
  RECT 494.600 1.600 498.510 3.460 ;
  LAYER VI2 ;
  RECT 479.800 1.600 492.060 3.460 ;
  LAYER VI2 ;
  RECT 474.600 1.600 477.430 3.460 ;
  LAYER VI2 ;
  RECT 460.200 1.600 472.220 3.460 ;
  LAYER VI2 ;
  RECT 453.800 1.600 457.590 3.460 ;
  LAYER VI2 ;
  RECT 439.000 1.600 451.140 3.460 ;
  LAYER VI2 ;
  RECT 433.800 1.600 436.510 3.460 ;
  LAYER VI2 ;
  RECT 419.000 1.600 431.300 3.460 ;
  LAYER VI2 ;
  RECT 412.600 1.600 416.670 3.460 ;
  LAYER VI2 ;
  RECT 398.200 1.600 410.220 3.460 ;
  LAYER VI2 ;
  RECT 393.000 1.600 395.590 3.460 ;
  LAYER VI2 ;
  RECT 378.200 1.600 390.380 3.460 ;
  LAYER VI2 ;
  RECT 371.800 1.600 375.750 3.460 ;
  LAYER VI2 ;
  RECT 357.000 1.600 369.300 3.460 ;
  LAYER VI2 ;
  RECT 351.800 1.600 354.670 3.460 ;
  LAYER VI2 ;
  RECT 339.000 1.600 349.460 3.460 ;
  LAYER VI2 ;
  RECT 331.000 1.600 334.830 3.460 ;
  LAYER VI2 ;
  RECT 316.200 1.600 328.380 3.460 ;
  LAYER VI2 ;
  RECT 311.000 1.600 313.750 3.460 ;
  LAYER VI2 ;
  RECT 296.600 1.600 308.540 3.460 ;
  LAYER VI2 ;
  RECT 289.800 1.600 293.910 3.460 ;
  LAYER VI2 ;
  RECT 275.400 1.600 287.460 3.460 ;
  LAYER VI2 ;
  RECT 270.200 1.600 272.830 3.460 ;
  LAYER VI2 ;
  RECT 255.400 1.600 267.620 3.460 ;
  LAYER VI2 ;
  RECT 249.000 1.600 252.990 3.460 ;
  LAYER VI2 ;
  RECT 234.600 1.600 246.540 3.460 ;
  LAYER VI2 ;
  RECT 229.000 1.600 231.910 3.460 ;
  LAYER VI2 ;
  RECT 214.600 1.600 226.700 3.460 ;
  LAYER VI2 ;
  RECT 208.200 1.600 212.070 3.460 ;
  LAYER VI2 ;
  RECT 193.400 1.600 205.620 3.460 ;
  LAYER VI2 ;
  RECT 188.200 1.600 190.990 3.460 ;
  LAYER VI2 ;
  RECT 175.400 1.600 185.780 3.460 ;
  LAYER VI2 ;
  RECT 167.000 1.600 171.150 3.460 ;
  LAYER VI2 ;
  RECT 152.600 1.600 164.700 3.460 ;
  LAYER VI2 ;
  RECT 147.400 1.600 150.070 3.460 ;
  LAYER VI2 ;
  RECT 132.600 1.600 144.860 3.460 ;
  LAYER VI2 ;
  RECT 126.200 1.600 130.230 3.460 ;
  LAYER VI2 ;
  RECT 111.800 1.600 123.780 3.460 ;
  LAYER VI2 ;
  RECT 106.600 1.600 109.150 3.460 ;
  LAYER VI2 ;
  RECT 91.800 1.600 103.940 3.460 ;
  LAYER VI2 ;
  RECT 85.400 1.600 89.310 3.460 ;
  LAYER VI2 ;
  RECT 70.600 1.600 82.860 3.460 ;
  LAYER VI2 ;
  RECT 65.400 1.600 68.230 3.460 ;
  LAYER VI2 ;
  RECT 51.000 1.600 63.020 3.460 ;
  LAYER VI2 ;
  RECT 44.600 1.600 48.390 3.460 ;
  LAYER VI2 ;
  RECT 29.800 1.600 41.940 3.460 ;
  LAYER VI2 ;
  RECT 24.600 1.600 27.310 3.460 ;
  LAYER VI2 ;
  RECT 11.800 1.600 22.100 3.460 ;
  LAYER VI2 ;
  RECT 2.000 1.600 7.470 3.460 ;
  LAYER VI1 ;
  RECT 2682.600 1.600 2691.080 3.460 ;
  LAYER VI1 ;
  RECT 2668.200 1.600 2680.280 3.460 ;
  LAYER VI1 ;
  RECT 2663.000 1.600 2665.650 3.460 ;
  LAYER VI1 ;
  RECT 2648.200 1.600 2660.440 3.460 ;
  LAYER VI1 ;
  RECT 2641.800 1.600 2645.810 3.460 ;
  LAYER VI1 ;
  RECT 2627.400 1.600 2639.360 3.460 ;
  LAYER VI1 ;
  RECT 2622.200 1.600 2624.730 3.460 ;
  LAYER VI1 ;
  RECT 2607.400 1.600 2619.520 3.460 ;
  LAYER VI1 ;
  RECT 2601.000 1.600 2604.890 3.460 ;
  LAYER VI1 ;
  RECT 2586.200 1.600 2598.440 3.460 ;
  LAYER VI1 ;
  RECT 2581.000 1.600 2583.810 3.460 ;
  LAYER VI1 ;
  RECT 2566.600 1.600 2578.600 3.460 ;
  LAYER VI1 ;
  RECT 2560.200 1.600 2563.970 3.460 ;
  LAYER VI1 ;
  RECT 2545.400 1.600 2557.520 3.460 ;
  LAYER VI1 ;
  RECT 2540.200 1.600 2542.890 3.460 ;
  LAYER VI1 ;
  RECT 2527.400 1.600 2537.680 3.460 ;
  LAYER VI1 ;
  RECT 2519.000 1.600 2523.050 3.460 ;
  LAYER VI1 ;
  RECT 2504.600 1.600 2516.600 3.460 ;
  LAYER VI1 ;
  RECT 2499.400 1.600 2501.970 3.460 ;
  LAYER VI1 ;
  RECT 2484.600 1.600 2496.760 3.460 ;
  LAYER VI1 ;
  RECT 2478.200 1.600 2482.130 3.460 ;
  LAYER VI1 ;
  RECT 2463.400 1.600 2475.680 3.460 ;
  LAYER VI1 ;
  RECT 2458.200 1.600 2461.050 3.460 ;
  LAYER VI1 ;
  RECT 2443.800 1.600 2455.840 3.460 ;
  LAYER VI1 ;
  RECT 2437.400 1.600 2441.210 3.460 ;
  LAYER VI1 ;
  RECT 2422.600 1.600 2434.760 3.460 ;
  LAYER VI1 ;
  RECT 2417.400 1.600 2420.130 3.460 ;
  LAYER VI1 ;
  RECT 2402.600 1.600 2414.920 3.460 ;
  LAYER VI1 ;
  RECT 2396.200 1.600 2400.290 3.460 ;
  LAYER VI1 ;
  RECT 2381.800 1.600 2393.840 3.460 ;
  LAYER VI1 ;
  RECT 2376.600 1.600 2379.210 3.460 ;
  LAYER VI1 ;
  RECT 2363.400 1.600 2374.000 3.460 ;
  LAYER VI1 ;
  RECT 2355.400 1.600 2359.370 3.460 ;
  LAYER VI1 ;
  RECT 2340.600 1.600 2352.920 3.460 ;
  LAYER VI1 ;
  RECT 2335.400 1.600 2338.290 3.460 ;
  LAYER VI1 ;
  RECT 2321.000 1.600 2333.080 3.460 ;
  LAYER VI1 ;
  RECT 2314.600 1.600 2318.450 3.460 ;
  LAYER VI1 ;
  RECT 2299.800 1.600 2312.000 3.460 ;
  LAYER VI1 ;
  RECT 2294.600 1.600 2297.370 3.460 ;
  LAYER VI1 ;
  RECT 2280.200 1.600 2292.160 3.460 ;
  LAYER VI1 ;
  RECT 2273.400 1.600 2277.530 3.460 ;
  LAYER VI1 ;
  RECT 2259.000 1.600 2271.080 3.460 ;
  LAYER VI1 ;
  RECT 2253.800 1.600 2256.450 3.460 ;
  LAYER VI1 ;
  RECT 2239.000 1.600 2251.240 3.460 ;
  LAYER VI1 ;
  RECT 2232.600 1.600 2236.610 3.460 ;
  LAYER VI1 ;
  RECT 2218.200 1.600 2230.160 3.460 ;
  LAYER VI1 ;
  RECT 2213.000 1.600 2215.530 3.460 ;
  LAYER VI1 ;
  RECT 2199.800 1.600 2210.320 3.460 ;
  LAYER VI1 ;
  RECT 2191.800 1.600 2195.690 3.460 ;
  LAYER VI1 ;
  RECT 2177.000 1.600 2189.240 3.460 ;
  LAYER VI1 ;
  RECT 2171.800 1.600 2174.610 3.460 ;
  LAYER VI1 ;
  RECT 2157.400 1.600 2169.400 3.460 ;
  LAYER VI1 ;
  RECT 2151.000 1.600 2154.770 3.460 ;
  LAYER VI1 ;
  RECT 2136.200 1.600 2148.320 3.460 ;
  LAYER VI1 ;
  RECT 2131.000 1.600 2133.690 3.460 ;
  LAYER VI1 ;
  RECT 2116.200 1.600 2128.480 3.460 ;
  LAYER VI1 ;
  RECT 2109.800 1.600 2113.850 3.460 ;
  LAYER VI1 ;
  RECT 2095.400 1.600 2107.400 3.460 ;
  LAYER VI1 ;
  RECT 2090.200 1.600 2092.770 3.460 ;
  LAYER VI1 ;
  RECT 2075.400 1.600 2087.560 3.460 ;
  LAYER VI1 ;
  RECT 2069.000 1.600 2072.930 3.460 ;
  LAYER VI1 ;
  RECT 2054.200 1.600 2066.480 3.460 ;
  LAYER VI1 ;
  RECT 2049.000 1.600 2051.850 3.460 ;
  LAYER VI1 ;
  RECT 2036.200 1.600 2046.640 3.460 ;
  LAYER VI1 ;
  RECT 2028.200 1.600 2032.010 3.460 ;
  LAYER VI1 ;
  RECT 2013.400 1.600 2025.560 3.460 ;
  LAYER VI1 ;
  RECT 2008.200 1.600 2010.930 3.460 ;
  LAYER VI1 ;
  RECT 1993.400 1.600 2005.720 3.460 ;
  LAYER VI1 ;
  RECT 1987.000 1.600 1991.090 3.460 ;
  LAYER VI1 ;
  RECT 1972.600 1.600 1984.640 3.460 ;
  LAYER VI1 ;
  RECT 1967.400 1.600 1970.010 3.460 ;
  LAYER VI1 ;
  RECT 1952.600 1.600 1964.800 3.460 ;
  LAYER VI1 ;
  RECT 1946.200 1.600 1950.170 3.460 ;
  LAYER VI1 ;
  RECT 1931.400 1.600 1943.720 3.460 ;
  LAYER VI1 ;
  RECT 1926.200 1.600 1929.090 3.460 ;
  LAYER VI1 ;
  RECT 1911.800 1.600 1923.880 3.460 ;
  LAYER VI1 ;
  RECT 1905.400 1.600 1909.250 3.460 ;
  LAYER VI1 ;
  RECT 1890.600 1.600 1902.800 3.460 ;
  LAYER VI1 ;
  RECT 1885.400 1.600 1888.170 3.460 ;
  LAYER VI1 ;
  RECT 1872.600 1.600 1882.960 3.460 ;
  LAYER VI1 ;
  RECT 1864.200 1.600 1868.330 3.460 ;
  LAYER VI1 ;
  RECT 1849.800 1.600 1861.880 3.460 ;
  LAYER VI1 ;
  RECT 1844.600 1.600 1847.250 3.460 ;
  LAYER VI1 ;
  RECT 1829.800 1.600 1842.040 3.460 ;
  LAYER VI1 ;
  RECT 1823.400 1.600 1827.410 3.460 ;
  LAYER VI1 ;
  RECT 1809.000 1.600 1820.960 3.460 ;
  LAYER VI1 ;
  RECT 1803.800 1.600 1806.330 3.460 ;
  LAYER VI1 ;
  RECT 1789.000 1.600 1801.120 3.460 ;
  LAYER VI1 ;
  RECT 1782.600 1.600 1786.490 3.460 ;
  LAYER VI1 ;
  RECT 1767.800 1.600 1780.040 3.460 ;
  LAYER VI1 ;
  RECT 1762.600 1.600 1765.410 3.460 ;
  LAYER VI1 ;
  RECT 1748.200 1.600 1760.200 3.460 ;
  LAYER VI1 ;
  RECT 1741.800 1.600 1745.570 3.460 ;
  LAYER VI1 ;
  RECT 1727.000 1.600 1739.120 3.460 ;
  LAYER VI1 ;
  RECT 1721.800 1.600 1724.490 3.460 ;
  LAYER VI1 ;
  RECT 1709.000 1.600 1719.280 3.460 ;
  LAYER VI1 ;
  RECT 1700.600 1.600 1704.650 3.460 ;
  LAYER VI1 ;
  RECT 1686.200 1.600 1698.200 3.460 ;
  LAYER VI1 ;
  RECT 1681.000 1.600 1683.570 3.460 ;
  LAYER VI1 ;
  RECT 1666.200 1.600 1678.360 3.460 ;
  LAYER VI1 ;
  RECT 1659.800 1.600 1663.730 3.460 ;
  LAYER VI1 ;
  RECT 1645.000 1.600 1657.280 3.460 ;
  LAYER VI1 ;
  RECT 1639.800 1.600 1642.650 3.460 ;
  LAYER VI1 ;
  RECT 1625.400 1.600 1637.440 3.460 ;
  LAYER VI1 ;
  RECT 1619.000 1.600 1622.810 3.460 ;
  LAYER VI1 ;
  RECT 1604.200 1.600 1616.360 3.460 ;
  LAYER VI1 ;
  RECT 1599.000 1.600 1601.730 3.460 ;
  LAYER VI1 ;
  RECT 1584.200 1.600 1596.520 3.460 ;
  LAYER VI1 ;
  RECT 1577.800 1.600 1581.890 3.460 ;
  LAYER VI1 ;
  RECT 1563.400 1.600 1575.440 3.460 ;
  LAYER VI1 ;
  RECT 1558.200 1.600 1560.810 3.460 ;
  LAYER VI1 ;
  RECT 1545.000 1.600 1555.600 3.460 ;
  LAYER VI1 ;
  RECT 1537.000 1.600 1540.970 3.460 ;
  LAYER VI1 ;
  RECT 1522.200 1.600 1534.520 3.460 ;
  LAYER VI1 ;
  RECT 1517.000 1.600 1519.890 3.460 ;
  LAYER VI1 ;
  RECT 1502.600 1.600 1514.680 3.460 ;
  LAYER VI1 ;
  RECT 1496.200 1.600 1500.050 3.460 ;
  LAYER VI1 ;
  RECT 1481.400 1.600 1493.600 3.460 ;
  LAYER VI1 ;
  RECT 1476.200 1.600 1478.970 3.460 ;
  LAYER VI1 ;
  RECT 1461.800 1.600 1473.760 3.460 ;
  LAYER VI1 ;
  RECT 1455.000 1.600 1459.130 3.460 ;
  LAYER VI1 ;
  RECT 1440.600 1.600 1452.680 3.460 ;
  LAYER VI1 ;
  RECT 1435.400 1.600 1438.050 3.460 ;
  LAYER VI1 ;
  RECT 1420.600 1.600 1432.840 3.460 ;
  LAYER VI1 ;
  RECT 1414.200 1.600 1418.210 3.460 ;
  LAYER VI1 ;
  RECT 1399.800 1.600 1411.760 3.460 ;
  LAYER VI1 ;
  RECT 1394.600 1.600 1397.130 3.460 ;
  LAYER VI1 ;
  RECT 1381.400 1.600 1391.920 3.460 ;
  LAYER VI1 ;
  RECT 1359.000 1.600 1377.290 3.460 ;
  LAYER VI1 ;
  RECT 1347.000 1.600 1350.450 3.460 ;
  LAYER VI1 ;
  RECT 1339.800 1.600 1344.480 3.460 ;
  LAYER VI1 ;
  RECT 1313.000 1.600 1319.840 3.460 ;
  LAYER VI1 ;
  RECT 1298.200 1.600 1310.460 3.460 ;
  LAYER VI1 ;
  RECT 1293.000 1.600 1295.830 3.460 ;
  LAYER VI1 ;
  RECT 1278.600 1.600 1290.620 3.460 ;
  LAYER VI1 ;
  RECT 1272.200 1.600 1275.990 3.460 ;
  LAYER VI1 ;
  RECT 1257.400 1.600 1269.540 3.460 ;
  LAYER VI1 ;
  RECT 1252.200 1.600 1254.910 3.460 ;
  LAYER VI1 ;
  RECT 1237.400 1.600 1249.700 3.460 ;
  LAYER VI1 ;
  RECT 1231.000 1.600 1235.070 3.460 ;
  LAYER VI1 ;
  RECT 1216.600 1.600 1228.620 3.460 ;
  LAYER VI1 ;
  RECT 1211.400 1.600 1213.990 3.460 ;
  LAYER VI1 ;
  RECT 1196.600 1.600 1208.780 3.460 ;
  LAYER VI1 ;
  RECT 1190.200 1.600 1194.150 3.460 ;
  LAYER VI1 ;
  RECT 1175.400 1.600 1187.700 3.460 ;
  LAYER VI1 ;
  RECT 1170.200 1.600 1173.070 3.460 ;
  LAYER VI1 ;
  RECT 1157.400 1.600 1167.860 3.460 ;
  LAYER VI1 ;
  RECT 1149.400 1.600 1153.230 3.460 ;
  LAYER VI1 ;
  RECT 1134.600 1.600 1146.780 3.460 ;
  LAYER VI1 ;
  RECT 1129.400 1.600 1132.150 3.460 ;
  LAYER VI1 ;
  RECT 1115.000 1.600 1126.940 3.460 ;
  LAYER VI1 ;
  RECT 1108.200 1.600 1112.310 3.460 ;
  LAYER VI1 ;
  RECT 1093.800 1.600 1105.860 3.460 ;
  LAYER VI1 ;
  RECT 1088.600 1.600 1091.230 3.460 ;
  LAYER VI1 ;
  RECT 1073.800 1.600 1086.020 3.460 ;
  LAYER VI1 ;
  RECT 1067.400 1.600 1071.390 3.460 ;
  LAYER VI1 ;
  RECT 1053.000 1.600 1064.940 3.460 ;
  LAYER VI1 ;
  RECT 1047.400 1.600 1050.310 3.460 ;
  LAYER VI1 ;
  RECT 1033.000 1.600 1045.100 3.460 ;
  LAYER VI1 ;
  RECT 1026.600 1.600 1030.470 3.460 ;
  LAYER VI1 ;
  RECT 1011.800 1.600 1024.020 3.460 ;
  LAYER VI1 ;
  RECT 1006.600 1.600 1009.390 3.460 ;
  LAYER VI1 ;
  RECT 993.800 1.600 1004.180 3.460 ;
  LAYER VI1 ;
  RECT 985.400 1.600 989.550 3.460 ;
  LAYER VI1 ;
  RECT 971.000 1.600 983.100 3.460 ;
  LAYER VI1 ;
  RECT 965.800 1.600 968.470 3.460 ;
  LAYER VI1 ;
  RECT 951.000 1.600 963.260 3.460 ;
  LAYER VI1 ;
  RECT 944.600 1.600 948.630 3.460 ;
  LAYER VI1 ;
  RECT 930.200 1.600 942.180 3.460 ;
  LAYER VI1 ;
  RECT 925.000 1.600 927.550 3.460 ;
  LAYER VI1 ;
  RECT 910.200 1.600 922.340 3.460 ;
  LAYER VI1 ;
  RECT 903.800 1.600 907.710 3.460 ;
  LAYER VI1 ;
  RECT 889.000 1.600 901.260 3.460 ;
  LAYER VI1 ;
  RECT 883.800 1.600 886.630 3.460 ;
  LAYER VI1 ;
  RECT 869.400 1.600 881.420 3.460 ;
  LAYER VI1 ;
  RECT 863.000 1.600 866.790 3.460 ;
  LAYER VI1 ;
  RECT 848.200 1.600 860.340 3.460 ;
  LAYER VI1 ;
  RECT 843.000 1.600 845.710 3.460 ;
  LAYER VI1 ;
  RECT 830.200 1.600 840.500 3.460 ;
  LAYER VI1 ;
  RECT 821.800 1.600 825.870 3.460 ;
  LAYER VI1 ;
  RECT 807.400 1.600 819.420 3.460 ;
  LAYER VI1 ;
  RECT 802.200 1.600 804.790 3.460 ;
  LAYER VI1 ;
  RECT 787.400 1.600 799.580 3.460 ;
  LAYER VI1 ;
  RECT 781.000 1.600 784.950 3.460 ;
  LAYER VI1 ;
  RECT 766.200 1.600 778.500 3.460 ;
  LAYER VI1 ;
  RECT 761.000 1.600 763.870 3.460 ;
  LAYER VI1 ;
  RECT 746.600 1.600 758.660 3.460 ;
  LAYER VI1 ;
  RECT 740.200 1.600 744.030 3.460 ;
  LAYER VI1 ;
  RECT 725.400 1.600 737.580 3.460 ;
  LAYER VI1 ;
  RECT 720.200 1.600 722.950 3.460 ;
  LAYER VI1 ;
  RECT 705.800 1.600 717.740 3.460 ;
  LAYER VI1 ;
  RECT 699.000 1.600 703.110 3.460 ;
  LAYER VI1 ;
  RECT 684.600 1.600 696.660 3.460 ;
  LAYER VI1 ;
  RECT 679.400 1.600 682.030 3.460 ;
  LAYER VI1 ;
  RECT 666.600 1.600 676.820 3.460 ;
  LAYER VI1 ;
  RECT 658.200 1.600 662.190 3.460 ;
  LAYER VI1 ;
  RECT 643.800 1.600 655.740 3.460 ;
  LAYER VI1 ;
  RECT 638.200 1.600 641.110 3.460 ;
  LAYER VI1 ;
  RECT 623.800 1.600 635.900 3.460 ;
  LAYER VI1 ;
  RECT 617.400 1.600 621.270 3.460 ;
  LAYER VI1 ;
  RECT 602.600 1.600 614.820 3.460 ;
  LAYER VI1 ;
  RECT 597.400 1.600 600.190 3.460 ;
  LAYER VI1 ;
  RECT 583.000 1.600 594.980 3.460 ;
  LAYER VI1 ;
  RECT 576.200 1.600 580.350 3.460 ;
  LAYER VI1 ;
  RECT 561.800 1.600 573.900 3.460 ;
  LAYER VI1 ;
  RECT 556.600 1.600 559.270 3.460 ;
  LAYER VI1 ;
  RECT 541.800 1.600 554.060 3.460 ;
  LAYER VI1 ;
  RECT 535.400 1.600 539.430 3.460 ;
  LAYER VI1 ;
  RECT 521.000 1.600 532.980 3.460 ;
  LAYER VI1 ;
  RECT 515.800 1.600 518.350 3.460 ;
  LAYER VI1 ;
  RECT 502.600 1.600 513.140 3.460 ;
  LAYER VI1 ;
  RECT 494.600 1.600 498.510 3.460 ;
  LAYER VI1 ;
  RECT 479.800 1.600 492.060 3.460 ;
  LAYER VI1 ;
  RECT 474.600 1.600 477.430 3.460 ;
  LAYER VI1 ;
  RECT 460.200 1.600 472.220 3.460 ;
  LAYER VI1 ;
  RECT 453.800 1.600 457.590 3.460 ;
  LAYER VI1 ;
  RECT 439.000 1.600 451.140 3.460 ;
  LAYER VI1 ;
  RECT 433.800 1.600 436.510 3.460 ;
  LAYER VI1 ;
  RECT 419.000 1.600 431.300 3.460 ;
  LAYER VI1 ;
  RECT 412.600 1.600 416.670 3.460 ;
  LAYER VI1 ;
  RECT 398.200 1.600 410.220 3.460 ;
  LAYER VI1 ;
  RECT 393.000 1.600 395.590 3.460 ;
  LAYER VI1 ;
  RECT 378.200 1.600 390.380 3.460 ;
  LAYER VI1 ;
  RECT 371.800 1.600 375.750 3.460 ;
  LAYER VI1 ;
  RECT 357.000 1.600 369.300 3.460 ;
  LAYER VI1 ;
  RECT 351.800 1.600 354.670 3.460 ;
  LAYER VI1 ;
  RECT 339.000 1.600 349.460 3.460 ;
  LAYER VI1 ;
  RECT 331.000 1.600 334.830 3.460 ;
  LAYER VI1 ;
  RECT 316.200 1.600 328.380 3.460 ;
  LAYER VI1 ;
  RECT 311.000 1.600 313.750 3.460 ;
  LAYER VI1 ;
  RECT 296.600 1.600 308.540 3.460 ;
  LAYER VI1 ;
  RECT 289.800 1.600 293.910 3.460 ;
  LAYER VI1 ;
  RECT 275.400 1.600 287.460 3.460 ;
  LAYER VI1 ;
  RECT 270.200 1.600 272.830 3.460 ;
  LAYER VI1 ;
  RECT 255.400 1.600 267.620 3.460 ;
  LAYER VI1 ;
  RECT 249.000 1.600 252.990 3.460 ;
  LAYER VI1 ;
  RECT 234.600 1.600 246.540 3.460 ;
  LAYER VI1 ;
  RECT 229.000 1.600 231.910 3.460 ;
  LAYER VI1 ;
  RECT 214.600 1.600 226.700 3.460 ;
  LAYER VI1 ;
  RECT 208.200 1.600 212.070 3.460 ;
  LAYER VI1 ;
  RECT 193.400 1.600 205.620 3.460 ;
  LAYER VI1 ;
  RECT 188.200 1.600 190.990 3.460 ;
  LAYER VI1 ;
  RECT 175.400 1.600 185.780 3.460 ;
  LAYER VI1 ;
  RECT 167.000 1.600 171.150 3.460 ;
  LAYER VI1 ;
  RECT 152.600 1.600 164.700 3.460 ;
  LAYER VI1 ;
  RECT 147.400 1.600 150.070 3.460 ;
  LAYER VI1 ;
  RECT 132.600 1.600 144.860 3.460 ;
  LAYER VI1 ;
  RECT 126.200 1.600 130.230 3.460 ;
  LAYER VI1 ;
  RECT 111.800 1.600 123.780 3.460 ;
  LAYER VI1 ;
  RECT 106.600 1.600 109.150 3.460 ;
  LAYER VI1 ;
  RECT 91.800 1.600 103.940 3.460 ;
  LAYER VI1 ;
  RECT 85.400 1.600 89.310 3.460 ;
  LAYER VI1 ;
  RECT 70.600 1.600 82.860 3.460 ;
  LAYER VI1 ;
  RECT 65.400 1.600 68.230 3.460 ;
  LAYER VI1 ;
  RECT 51.000 1.600 63.020 3.460 ;
  LAYER VI1 ;
  RECT 44.600 1.600 48.390 3.460 ;
  LAYER VI1 ;
  RECT 29.800 1.600 41.940 3.460 ;
  LAYER VI1 ;
  RECT 24.600 1.600 27.310 3.460 ;
  LAYER VI1 ;
  RECT 11.800 1.600 22.100 3.460 ;
  LAYER VI1 ;
  RECT 1.860 1.600 7.470 3.460 ;
  LAYER VI3 ;
  RECT 2688.940 555.000 2690.660 561.930 ;
  LAYER VI3 ;
  RECT 2688.940 64.930 2690.660 67.240 ;
  LAYER VI3 ;
  RECT 2688.940 44.080 2690.660 61.260 ;
  LAYER VI3 ;
  RECT 2688.940 39.620 2690.660 41.480 ;
  LAYER VI3 ;
  RECT 2688.940 29.870 2690.660 33.520 ;
  LAYER VI3 ;
  RECT 2688.940 24.270 2690.660 26.870 ;
  LAYER VI3 ;
  RECT 2688.940 18.130 2690.660 21.270 ;
  LAYER VI3 ;
  RECT 2688.940 5.600 2690.660 11.230 ;
  LAYER VI2 ;
  RECT 2688.940 555.000 2690.660 561.930 ;
  LAYER VI2 ;
  RECT 2688.940 64.930 2690.660 67.240 ;
  LAYER VI2 ;
  RECT 2688.940 44.080 2690.660 61.260 ;
  LAYER VI2 ;
  RECT 2688.940 39.620 2690.660 41.480 ;
  LAYER VI2 ;
  RECT 2688.940 29.870 2690.660 33.520 ;
  LAYER VI2 ;
  RECT 2688.940 24.270 2690.660 26.870 ;
  LAYER VI2 ;
  RECT 2688.940 18.130 2690.660 21.270 ;
  LAYER VI2 ;
  RECT 2688.940 5.600 2690.660 11.230 ;
  LAYER VI1 ;
  RECT 2688.940 5.600 2690.800 561.930 ;
  LAYER VI3 ;
  RECT 2.280 555.000 4.000 561.930 ;
  LAYER VI3 ;
  RECT 2.280 64.930 4.000 67.240 ;
  LAYER VI3 ;
  RECT 2.280 44.080 4.000 61.260 ;
  LAYER VI3 ;
  RECT 2.280 39.620 4.000 41.480 ;
  LAYER VI3 ;
  RECT 2.280 29.870 4.000 33.520 ;
  LAYER VI3 ;
  RECT 2.280 24.270 4.000 26.870 ;
  LAYER VI3 ;
  RECT 2.280 18.130 4.000 21.270 ;
  LAYER VI3 ;
  RECT 2.280 5.600 4.000 11.230 ;
  LAYER VI2 ;
  RECT 2.280 555.000 4.000 561.930 ;
  LAYER VI2 ;
  RECT 2.280 64.930 4.000 67.240 ;
  LAYER VI2 ;
  RECT 2.280 44.080 4.000 61.260 ;
  LAYER VI2 ;
  RECT 2.280 39.620 4.000 41.480 ;
  LAYER VI2 ;
  RECT 2.280 29.870 4.000 33.520 ;
  LAYER VI2 ;
  RECT 2.280 24.270 4.000 26.870 ;
  LAYER VI2 ;
  RECT 2.280 18.130 4.000 21.270 ;
  LAYER VI2 ;
  RECT 2.280 5.600 4.000 11.230 ;
  LAYER VI1 ;
  RECT 2.140 5.600 4.000 561.930 ;
  LAYER VI3 ;
  RECT 2646.020 561.930 2688.940 563.650 ;
  LAYER VI3 ;
  RECT 2605.100 561.930 2643.770 563.650 ;
  LAYER VI3 ;
  RECT 2564.180 561.930 2602.850 563.650 ;
  LAYER VI3 ;
  RECT 2523.260 561.930 2561.930 563.650 ;
  LAYER VI3 ;
  RECT 2482.340 561.930 2521.010 563.650 ;
  LAYER VI3 ;
  RECT 2441.420 561.930 2480.090 563.650 ;
  LAYER VI3 ;
  RECT 2400.500 561.930 2439.170 563.650 ;
  LAYER VI3 ;
  RECT 2359.580 561.930 2398.250 563.650 ;
  LAYER VI3 ;
  RECT 2318.660 561.930 2357.330 563.650 ;
  LAYER VI3 ;
  RECT 2277.740 561.930 2316.410 563.650 ;
  LAYER VI3 ;
  RECT 2236.820 561.930 2275.490 563.650 ;
  LAYER VI3 ;
  RECT 2195.900 561.930 2234.570 563.650 ;
  LAYER VI3 ;
  RECT 2154.980 561.930 2193.650 563.650 ;
  LAYER VI3 ;
  RECT 2114.060 561.930 2152.730 563.650 ;
  LAYER VI3 ;
  RECT 2073.140 561.930 2111.810 563.650 ;
  LAYER VI3 ;
  RECT 2032.220 561.930 2070.890 563.650 ;
  LAYER VI3 ;
  RECT 1991.300 561.930 2029.970 563.650 ;
  LAYER VI3 ;
  RECT 1950.380 561.930 1989.050 563.650 ;
  LAYER VI3 ;
  RECT 1909.460 561.930 1948.130 563.650 ;
  LAYER VI3 ;
  RECT 1868.540 561.930 1907.210 563.650 ;
  LAYER VI3 ;
  RECT 1827.620 561.930 1866.290 563.650 ;
  LAYER VI3 ;
  RECT 1786.700 561.930 1825.370 563.650 ;
  LAYER VI3 ;
  RECT 1745.780 561.930 1784.450 563.650 ;
  LAYER VI3 ;
  RECT 1704.860 561.930 1743.530 563.650 ;
  LAYER VI3 ;
  RECT 1663.940 561.930 1702.610 563.650 ;
  LAYER VI3 ;
  RECT 1623.020 561.930 1661.690 563.650 ;
  LAYER VI3 ;
  RECT 1582.100 561.930 1620.770 563.650 ;
  LAYER VI3 ;
  RECT 1541.180 561.930 1579.850 563.650 ;
  LAYER VI3 ;
  RECT 1500.260 561.930 1538.930 563.650 ;
  LAYER VI3 ;
  RECT 1459.340 561.930 1498.010 563.650 ;
  LAYER VI3 ;
  RECT 1418.420 561.930 1457.090 563.650 ;
  LAYER VI3 ;
  RECT 1377.500 561.930 1416.170 563.650 ;
  LAYER VI3 ;
  RECT 1358.760 561.930 1371.760 563.650 ;
  LAYER VI3 ;
  RECT 1347.630 561.930 1352.440 563.650 ;
  LAYER VI3 ;
  RECT 1337.920 561.930 1342.440 563.650 ;
  LAYER VI3 ;
  RECT 1332.580 561.930 1334.160 563.650 ;
  LAYER VI3 ;
  RECT 1276.770 561.930 1315.800 563.650 ;
  LAYER VI3 ;
  RECT 1235.850 561.930 1274.520 563.650 ;
  LAYER VI3 ;
  RECT 1194.930 561.930 1233.600 563.650 ;
  LAYER VI3 ;
  RECT 1154.010 561.930 1192.680 563.650 ;
  LAYER VI3 ;
  RECT 1113.090 561.930 1151.760 563.650 ;
  LAYER VI3 ;
  RECT 1072.170 561.930 1110.840 563.650 ;
  LAYER VI3 ;
  RECT 1031.250 561.930 1069.920 563.650 ;
  LAYER VI3 ;
  RECT 990.330 561.930 1029.000 563.650 ;
  LAYER VI3 ;
  RECT 949.410 561.930 988.080 563.650 ;
  LAYER VI3 ;
  RECT 908.490 561.930 947.160 563.650 ;
  LAYER VI3 ;
  RECT 867.570 561.930 906.240 563.650 ;
  LAYER VI3 ;
  RECT 826.650 561.930 865.320 563.650 ;
  LAYER VI3 ;
  RECT 785.730 561.930 824.400 563.650 ;
  LAYER VI3 ;
  RECT 744.810 561.930 783.480 563.650 ;
  LAYER VI3 ;
  RECT 703.890 561.930 742.560 563.650 ;
  LAYER VI3 ;
  RECT 662.970 561.930 701.640 563.650 ;
  LAYER VI3 ;
  RECT 622.050 561.930 660.720 563.650 ;
  LAYER VI3 ;
  RECT 581.130 561.930 619.800 563.650 ;
  LAYER VI3 ;
  RECT 540.210 561.930 578.880 563.650 ;
  LAYER VI3 ;
  RECT 499.290 561.930 537.960 563.650 ;
  LAYER VI3 ;
  RECT 458.370 561.930 497.040 563.650 ;
  LAYER VI3 ;
  RECT 417.450 561.930 456.120 563.650 ;
  LAYER VI3 ;
  RECT 376.530 561.930 415.200 563.650 ;
  LAYER VI3 ;
  RECT 335.610 561.930 374.280 563.650 ;
  LAYER VI3 ;
  RECT 294.690 561.930 333.360 563.650 ;
  LAYER VI3 ;
  RECT 253.770 561.930 292.440 563.650 ;
  LAYER VI3 ;
  RECT 212.850 561.930 251.520 563.650 ;
  LAYER VI3 ;
  RECT 171.930 561.930 210.600 563.650 ;
  LAYER VI3 ;
  RECT 131.010 561.930 169.680 563.650 ;
  LAYER VI3 ;
  RECT 90.090 561.930 128.760 563.650 ;
  LAYER VI3 ;
  RECT 49.170 561.930 87.840 563.650 ;
  LAYER VI3 ;
  RECT 4.000 561.930 46.920 563.650 ;
  LAYER VI2 ;
  RECT 2646.020 561.930 2688.940 563.650 ;
  LAYER VI2 ;
  RECT 2605.100 561.930 2643.770 563.650 ;
  LAYER VI2 ;
  RECT 2564.180 561.930 2602.850 563.650 ;
  LAYER VI2 ;
  RECT 2523.260 561.930 2561.930 563.650 ;
  LAYER VI2 ;
  RECT 2482.340 561.930 2521.010 563.650 ;
  LAYER VI2 ;
  RECT 2441.420 561.930 2480.090 563.650 ;
  LAYER VI2 ;
  RECT 2400.500 561.930 2439.170 563.650 ;
  LAYER VI2 ;
  RECT 2359.580 561.930 2398.250 563.650 ;
  LAYER VI2 ;
  RECT 2318.660 561.930 2357.330 563.650 ;
  LAYER VI2 ;
  RECT 2277.740 561.930 2316.410 563.650 ;
  LAYER VI2 ;
  RECT 2236.820 561.930 2275.490 563.650 ;
  LAYER VI2 ;
  RECT 2195.900 561.930 2234.570 563.650 ;
  LAYER VI2 ;
  RECT 2154.980 561.930 2193.650 563.650 ;
  LAYER VI2 ;
  RECT 2114.060 561.930 2152.730 563.650 ;
  LAYER VI2 ;
  RECT 2073.140 561.930 2111.810 563.650 ;
  LAYER VI2 ;
  RECT 2032.220 561.930 2070.890 563.650 ;
  LAYER VI2 ;
  RECT 1991.300 561.930 2029.970 563.650 ;
  LAYER VI2 ;
  RECT 1950.380 561.930 1989.050 563.650 ;
  LAYER VI2 ;
  RECT 1909.460 561.930 1948.130 563.650 ;
  LAYER VI2 ;
  RECT 1868.540 561.930 1907.210 563.650 ;
  LAYER VI2 ;
  RECT 1827.620 561.930 1866.290 563.650 ;
  LAYER VI2 ;
  RECT 1786.700 561.930 1825.370 563.650 ;
  LAYER VI2 ;
  RECT 1745.780 561.930 1784.450 563.650 ;
  LAYER VI2 ;
  RECT 1704.860 561.930 1743.530 563.650 ;
  LAYER VI2 ;
  RECT 1663.940 561.930 1702.610 563.650 ;
  LAYER VI2 ;
  RECT 1623.020 561.930 1661.690 563.650 ;
  LAYER VI2 ;
  RECT 1582.100 561.930 1620.770 563.650 ;
  LAYER VI2 ;
  RECT 1541.180 561.930 1579.850 563.650 ;
  LAYER VI2 ;
  RECT 1500.260 561.930 1538.930 563.650 ;
  LAYER VI2 ;
  RECT 1459.340 561.930 1498.010 563.650 ;
  LAYER VI2 ;
  RECT 1418.420 561.930 1457.090 563.650 ;
  LAYER VI2 ;
  RECT 1377.500 561.930 1416.170 563.650 ;
  LAYER VI2 ;
  RECT 1358.760 561.930 1371.760 563.650 ;
  LAYER VI2 ;
  RECT 1347.630 561.930 1352.440 563.650 ;
  LAYER VI2 ;
  RECT 1337.920 561.930 1342.440 563.650 ;
  LAYER VI2 ;
  RECT 1332.580 561.930 1334.160 563.650 ;
  LAYER VI2 ;
  RECT 1276.770 561.930 1315.800 563.650 ;
  LAYER VI2 ;
  RECT 1235.850 561.930 1274.520 563.650 ;
  LAYER VI2 ;
  RECT 1194.930 561.930 1233.600 563.650 ;
  LAYER VI2 ;
  RECT 1154.010 561.930 1192.680 563.650 ;
  LAYER VI2 ;
  RECT 1113.090 561.930 1151.760 563.650 ;
  LAYER VI2 ;
  RECT 1072.170 561.930 1110.840 563.650 ;
  LAYER VI2 ;
  RECT 1031.250 561.930 1069.920 563.650 ;
  LAYER VI2 ;
  RECT 990.330 561.930 1029.000 563.650 ;
  LAYER VI2 ;
  RECT 949.410 561.930 988.080 563.650 ;
  LAYER VI2 ;
  RECT 908.490 561.930 947.160 563.650 ;
  LAYER VI2 ;
  RECT 867.570 561.930 906.240 563.650 ;
  LAYER VI2 ;
  RECT 826.650 561.930 865.320 563.650 ;
  LAYER VI2 ;
  RECT 785.730 561.930 824.400 563.650 ;
  LAYER VI2 ;
  RECT 744.810 561.930 783.480 563.650 ;
  LAYER VI2 ;
  RECT 703.890 561.930 742.560 563.650 ;
  LAYER VI2 ;
  RECT 662.970 561.930 701.640 563.650 ;
  LAYER VI2 ;
  RECT 622.050 561.930 660.720 563.650 ;
  LAYER VI2 ;
  RECT 581.130 561.930 619.800 563.650 ;
  LAYER VI2 ;
  RECT 540.210 561.930 578.880 563.650 ;
  LAYER VI2 ;
  RECT 499.290 561.930 537.960 563.650 ;
  LAYER VI2 ;
  RECT 458.370 561.930 497.040 563.650 ;
  LAYER VI2 ;
  RECT 417.450 561.930 456.120 563.650 ;
  LAYER VI2 ;
  RECT 376.530 561.930 415.200 563.650 ;
  LAYER VI2 ;
  RECT 335.610 561.930 374.280 563.650 ;
  LAYER VI2 ;
  RECT 294.690 561.930 333.360 563.650 ;
  LAYER VI2 ;
  RECT 253.770 561.930 292.440 563.650 ;
  LAYER VI2 ;
  RECT 212.850 561.930 251.520 563.650 ;
  LAYER VI2 ;
  RECT 171.930 561.930 210.600 563.650 ;
  LAYER VI2 ;
  RECT 131.010 561.930 169.680 563.650 ;
  LAYER VI2 ;
  RECT 90.090 561.930 128.760 563.650 ;
  LAYER VI2 ;
  RECT 49.170 561.930 87.840 563.650 ;
  LAYER VI2 ;
  RECT 4.000 561.930 46.920 563.650 ;
  LAYER VI1 ;
  RECT 4.000 561.930 2688.940 563.790 ;
  LAYER VI3 ;
  RECT 2675.540 3.880 2685.380 5.600 ;
  LAYER VI3 ;
  RECT 2655.700 3.880 2665.540 5.600 ;
  LAYER VI3 ;
  RECT 2634.620 3.880 2645.700 5.600 ;
  LAYER VI3 ;
  RECT 2614.780 3.880 2624.620 5.600 ;
  LAYER VI3 ;
  RECT 2593.700 3.880 2604.780 5.600 ;
  LAYER VI3 ;
  RECT 2573.860 3.880 2583.700 5.600 ;
  LAYER VI3 ;
  RECT 2552.780 3.880 2563.860 5.600 ;
  LAYER VI3 ;
  RECT 2532.940 3.880 2542.780 5.600 ;
  LAYER VI3 ;
  RECT 2511.860 3.880 2522.940 5.600 ;
  LAYER VI3 ;
  RECT 2492.020 3.880 2501.860 5.600 ;
  LAYER VI3 ;
  RECT 2470.940 3.880 2482.020 5.600 ;
  LAYER VI3 ;
  RECT 2451.100 3.880 2460.940 5.600 ;
  LAYER VI3 ;
  RECT 2430.020 3.880 2441.100 5.600 ;
  LAYER VI3 ;
  RECT 2410.180 3.880 2420.020 5.600 ;
  LAYER VI3 ;
  RECT 2389.100 3.880 2400.180 5.600 ;
  LAYER VI3 ;
  RECT 2369.260 3.880 2379.100 5.600 ;
  LAYER VI3 ;
  RECT 2348.180 3.880 2359.260 5.600 ;
  LAYER VI3 ;
  RECT 2328.340 3.880 2338.180 5.600 ;
  LAYER VI3 ;
  RECT 2307.260 3.880 2318.340 5.600 ;
  LAYER VI3 ;
  RECT 2287.420 3.880 2297.260 5.600 ;
  LAYER VI3 ;
  RECT 2266.340 3.880 2277.420 5.600 ;
  LAYER VI3 ;
  RECT 2246.500 3.880 2256.340 5.600 ;
  LAYER VI3 ;
  RECT 2225.420 3.880 2236.500 5.600 ;
  LAYER VI3 ;
  RECT 2205.580 3.880 2215.420 5.600 ;
  LAYER VI3 ;
  RECT 2184.500 3.880 2195.580 5.600 ;
  LAYER VI3 ;
  RECT 2164.660 3.880 2174.500 5.600 ;
  LAYER VI3 ;
  RECT 2143.580 3.880 2154.660 5.600 ;
  LAYER VI3 ;
  RECT 2123.740 3.880 2133.580 5.600 ;
  LAYER VI3 ;
  RECT 2102.660 3.880 2113.740 5.600 ;
  LAYER VI3 ;
  RECT 2082.820 3.880 2092.660 5.600 ;
  LAYER VI3 ;
  RECT 2061.740 3.880 2072.820 5.600 ;
  LAYER VI3 ;
  RECT 2041.900 3.880 2051.740 5.600 ;
  LAYER VI3 ;
  RECT 2020.820 3.880 2031.900 5.600 ;
  LAYER VI3 ;
  RECT 2000.980 3.880 2010.820 5.600 ;
  LAYER VI3 ;
  RECT 1979.900 3.880 1990.980 5.600 ;
  LAYER VI3 ;
  RECT 1960.060 3.880 1969.900 5.600 ;
  LAYER VI3 ;
  RECT 1938.980 3.880 1950.060 5.600 ;
  LAYER VI3 ;
  RECT 1919.140 3.880 1928.980 5.600 ;
  LAYER VI3 ;
  RECT 1898.060 3.880 1909.140 5.600 ;
  LAYER VI3 ;
  RECT 1878.220 3.880 1888.060 5.600 ;
  LAYER VI3 ;
  RECT 1857.140 3.880 1868.220 5.600 ;
  LAYER VI3 ;
  RECT 1837.300 3.880 1847.140 5.600 ;
  LAYER VI3 ;
  RECT 1816.220 3.880 1827.300 5.600 ;
  LAYER VI3 ;
  RECT 1796.380 3.880 1806.220 5.600 ;
  LAYER VI3 ;
  RECT 1775.300 3.880 1786.380 5.600 ;
  LAYER VI3 ;
  RECT 1755.460 3.880 1765.300 5.600 ;
  LAYER VI3 ;
  RECT 1734.380 3.880 1745.460 5.600 ;
  LAYER VI3 ;
  RECT 1714.540 3.880 1724.380 5.600 ;
  LAYER VI3 ;
  RECT 1693.460 3.880 1704.540 5.600 ;
  LAYER VI3 ;
  RECT 1673.620 3.880 1683.460 5.600 ;
  LAYER VI3 ;
  RECT 1652.540 3.880 1663.620 5.600 ;
  LAYER VI3 ;
  RECT 1632.700 3.880 1642.540 5.600 ;
  LAYER VI3 ;
  RECT 1611.620 3.880 1622.700 5.600 ;
  LAYER VI3 ;
  RECT 1591.780 3.880 1601.620 5.600 ;
  LAYER VI3 ;
  RECT 1570.700 3.880 1581.780 5.600 ;
  LAYER VI3 ;
  RECT 1550.860 3.880 1560.700 5.600 ;
  LAYER VI3 ;
  RECT 1529.780 3.880 1540.860 5.600 ;
  LAYER VI3 ;
  RECT 1509.940 3.880 1519.780 5.600 ;
  LAYER VI3 ;
  RECT 1488.860 3.880 1499.940 5.600 ;
  LAYER VI3 ;
  RECT 1469.020 3.880 1478.860 5.600 ;
  LAYER VI3 ;
  RECT 1447.940 3.880 1459.020 5.600 ;
  LAYER VI3 ;
  RECT 1428.100 3.880 1437.940 5.600 ;
  LAYER VI3 ;
  RECT 1407.020 3.880 1418.100 5.600 ;
  LAYER VI3 ;
  RECT 1387.180 3.880 1397.020 5.600 ;
  LAYER VI3 ;
  RECT 1359.210 3.880 1377.180 5.600 ;
  LAYER VI3 ;
  RECT 1347.890 3.880 1351.290 5.600 ;
  LAYER VI3 ;
  RECT 1337.920 3.880 1342.440 5.600 ;
  LAYER VI3 ;
  RECT 1332.580 3.880 1334.160 5.600 ;
  LAYER VI3 ;
  RECT 1305.720 3.880 1316.820 5.600 ;
  LAYER VI3 ;
  RECT 1285.880 3.880 1295.720 5.600 ;
  LAYER VI3 ;
  RECT 1264.800 3.880 1275.880 5.600 ;
  LAYER VI3 ;
  RECT 1244.960 3.880 1254.800 5.600 ;
  LAYER VI3 ;
  RECT 1223.880 3.880 1234.960 5.600 ;
  LAYER VI3 ;
  RECT 1204.040 3.880 1213.880 5.600 ;
  LAYER VI3 ;
  RECT 1182.960 3.880 1194.040 5.600 ;
  LAYER VI3 ;
  RECT 1163.120 3.880 1172.960 5.600 ;
  LAYER VI3 ;
  RECT 1142.040 3.880 1153.120 5.600 ;
  LAYER VI3 ;
  RECT 1122.200 3.880 1132.040 5.600 ;
  LAYER VI3 ;
  RECT 1101.120 3.880 1112.200 5.600 ;
  LAYER VI3 ;
  RECT 1081.280 3.880 1091.120 5.600 ;
  LAYER VI3 ;
  RECT 1060.200 3.880 1071.280 5.600 ;
  LAYER VI3 ;
  RECT 1040.360 3.880 1050.200 5.600 ;
  LAYER VI3 ;
  RECT 1019.280 3.880 1030.360 5.600 ;
  LAYER VI3 ;
  RECT 999.440 3.880 1009.280 5.600 ;
  LAYER VI3 ;
  RECT 978.360 3.880 989.440 5.600 ;
  LAYER VI3 ;
  RECT 958.520 3.880 968.360 5.600 ;
  LAYER VI3 ;
  RECT 937.440 3.880 948.520 5.600 ;
  LAYER VI3 ;
  RECT 917.600 3.880 927.440 5.600 ;
  LAYER VI3 ;
  RECT 896.520 3.880 907.600 5.600 ;
  LAYER VI3 ;
  RECT 876.680 3.880 886.520 5.600 ;
  LAYER VI3 ;
  RECT 855.600 3.880 866.680 5.600 ;
  LAYER VI3 ;
  RECT 835.760 3.880 845.600 5.600 ;
  LAYER VI3 ;
  RECT 814.680 3.880 825.760 5.600 ;
  LAYER VI3 ;
  RECT 794.840 3.880 804.680 5.600 ;
  LAYER VI3 ;
  RECT 773.760 3.880 784.840 5.600 ;
  LAYER VI3 ;
  RECT 753.920 3.880 763.760 5.600 ;
  LAYER VI3 ;
  RECT 732.840 3.880 743.920 5.600 ;
  LAYER VI3 ;
  RECT 713.000 3.880 722.840 5.600 ;
  LAYER VI3 ;
  RECT 691.920 3.880 703.000 5.600 ;
  LAYER VI3 ;
  RECT 672.080 3.880 681.920 5.600 ;
  LAYER VI3 ;
  RECT 651.000 3.880 662.080 5.600 ;
  LAYER VI3 ;
  RECT 631.160 3.880 641.000 5.600 ;
  LAYER VI3 ;
  RECT 610.080 3.880 621.160 5.600 ;
  LAYER VI3 ;
  RECT 590.240 3.880 600.080 5.600 ;
  LAYER VI3 ;
  RECT 569.160 3.880 580.240 5.600 ;
  LAYER VI3 ;
  RECT 549.320 3.880 559.160 5.600 ;
  LAYER VI3 ;
  RECT 528.240 3.880 539.320 5.600 ;
  LAYER VI3 ;
  RECT 508.400 3.880 518.240 5.600 ;
  LAYER VI3 ;
  RECT 487.320 3.880 498.400 5.600 ;
  LAYER VI3 ;
  RECT 467.480 3.880 477.320 5.600 ;
  LAYER VI3 ;
  RECT 446.400 3.880 457.480 5.600 ;
  LAYER VI3 ;
  RECT 426.560 3.880 436.400 5.600 ;
  LAYER VI3 ;
  RECT 405.480 3.880 416.560 5.600 ;
  LAYER VI3 ;
  RECT 385.640 3.880 395.480 5.600 ;
  LAYER VI3 ;
  RECT 364.560 3.880 375.640 5.600 ;
  LAYER VI3 ;
  RECT 344.720 3.880 354.560 5.600 ;
  LAYER VI3 ;
  RECT 323.640 3.880 334.720 5.600 ;
  LAYER VI3 ;
  RECT 303.800 3.880 313.640 5.600 ;
  LAYER VI3 ;
  RECT 282.720 3.880 293.800 5.600 ;
  LAYER VI3 ;
  RECT 262.880 3.880 272.720 5.600 ;
  LAYER VI3 ;
  RECT 241.800 3.880 252.880 5.600 ;
  LAYER VI3 ;
  RECT 221.960 3.880 231.800 5.600 ;
  LAYER VI3 ;
  RECT 200.880 3.880 211.960 5.600 ;
  LAYER VI3 ;
  RECT 181.040 3.880 190.880 5.600 ;
  LAYER VI3 ;
  RECT 159.960 3.880 171.040 5.600 ;
  LAYER VI3 ;
  RECT 140.120 3.880 149.960 5.600 ;
  LAYER VI3 ;
  RECT 119.040 3.880 130.120 5.600 ;
  LAYER VI3 ;
  RECT 99.200 3.880 109.040 5.600 ;
  LAYER VI3 ;
  RECT 78.120 3.880 89.200 5.600 ;
  LAYER VI3 ;
  RECT 58.280 3.880 68.120 5.600 ;
  LAYER VI3 ;
  RECT 37.200 3.880 48.280 5.600 ;
  LAYER VI3 ;
  RECT 17.360 3.880 27.200 5.600 ;
  LAYER VI2 ;
  RECT 2682.600 3.880 2685.380 5.600 ;
  LAYER VI2 ;
  RECT 2675.540 3.880 2680.280 5.600 ;
  LAYER VI2 ;
  RECT 2663.000 3.880 2665.540 5.600 ;
  LAYER VI2 ;
  RECT 2655.700 3.880 2660.440 5.600 ;
  LAYER VI2 ;
  RECT 2641.800 3.880 2645.700 5.600 ;
  LAYER VI2 ;
  RECT 2634.620 3.880 2639.360 5.600 ;
  LAYER VI2 ;
  RECT 2622.200 3.880 2624.620 5.600 ;
  LAYER VI2 ;
  RECT 2614.780 3.880 2619.520 5.600 ;
  LAYER VI2 ;
  RECT 2601.000 3.880 2604.780 5.600 ;
  LAYER VI2 ;
  RECT 2593.700 3.880 2598.440 5.600 ;
  LAYER VI2 ;
  RECT 2581.000 3.880 2583.700 5.600 ;
  LAYER VI2 ;
  RECT 2573.860 3.880 2578.600 5.600 ;
  LAYER VI2 ;
  RECT 2560.200 3.880 2563.860 5.600 ;
  LAYER VI2 ;
  RECT 2552.780 3.880 2557.520 5.600 ;
  LAYER VI2 ;
  RECT 2540.200 3.880 2542.780 5.600 ;
  LAYER VI2 ;
  RECT 2532.940 3.880 2537.680 5.600 ;
  LAYER VI2 ;
  RECT 2519.000 3.880 2522.940 5.600 ;
  LAYER VI2 ;
  RECT 2511.860 3.880 2516.600 5.600 ;
  LAYER VI2 ;
  RECT 2499.400 3.880 2501.860 5.600 ;
  LAYER VI2 ;
  RECT 2492.020 3.880 2496.760 5.600 ;
  LAYER VI2 ;
  RECT 2478.200 3.880 2482.020 5.600 ;
  LAYER VI2 ;
  RECT 2470.940 3.880 2475.680 5.600 ;
  LAYER VI2 ;
  RECT 2458.200 3.880 2460.940 5.600 ;
  LAYER VI2 ;
  RECT 2451.100 3.880 2455.840 5.600 ;
  LAYER VI2 ;
  RECT 2437.400 3.880 2441.100 5.600 ;
  LAYER VI2 ;
  RECT 2430.020 3.880 2434.760 5.600 ;
  LAYER VI2 ;
  RECT 2417.400 3.880 2420.020 5.600 ;
  LAYER VI2 ;
  RECT 2410.180 3.880 2414.920 5.600 ;
  LAYER VI2 ;
  RECT 2396.200 3.880 2400.180 5.600 ;
  LAYER VI2 ;
  RECT 2389.100 3.880 2393.840 5.600 ;
  LAYER VI2 ;
  RECT 2376.600 3.880 2379.100 5.600 ;
  LAYER VI2 ;
  RECT 2369.260 3.880 2374.000 5.600 ;
  LAYER VI2 ;
  RECT 2355.400 3.880 2359.260 5.600 ;
  LAYER VI2 ;
  RECT 2348.180 3.880 2352.920 5.600 ;
  LAYER VI2 ;
  RECT 2335.400 3.880 2338.180 5.600 ;
  LAYER VI2 ;
  RECT 2328.340 3.880 2333.080 5.600 ;
  LAYER VI2 ;
  RECT 2314.600 3.880 2318.340 5.600 ;
  LAYER VI2 ;
  RECT 2307.260 3.880 2312.000 5.600 ;
  LAYER VI2 ;
  RECT 2294.600 3.880 2297.260 5.600 ;
  LAYER VI2 ;
  RECT 2287.420 3.880 2292.160 5.600 ;
  LAYER VI2 ;
  RECT 2273.400 3.880 2277.420 5.600 ;
  LAYER VI2 ;
  RECT 2266.340 3.880 2271.080 5.600 ;
  LAYER VI2 ;
  RECT 2253.800 3.880 2256.340 5.600 ;
  LAYER VI2 ;
  RECT 2246.500 3.880 2251.240 5.600 ;
  LAYER VI2 ;
  RECT 2232.600 3.880 2236.500 5.600 ;
  LAYER VI2 ;
  RECT 2225.420 3.880 2230.160 5.600 ;
  LAYER VI2 ;
  RECT 2213.000 3.880 2215.420 5.600 ;
  LAYER VI2 ;
  RECT 2205.580 3.880 2210.320 5.600 ;
  LAYER VI2 ;
  RECT 2191.800 3.880 2195.580 5.600 ;
  LAYER VI2 ;
  RECT 2184.500 3.880 2189.240 5.600 ;
  LAYER VI2 ;
  RECT 2171.800 3.880 2174.500 5.600 ;
  LAYER VI2 ;
  RECT 2164.660 3.880 2169.400 5.600 ;
  LAYER VI2 ;
  RECT 2151.000 3.880 2154.660 5.600 ;
  LAYER VI2 ;
  RECT 2143.580 3.880 2148.320 5.600 ;
  LAYER VI2 ;
  RECT 2131.000 3.880 2133.580 5.600 ;
  LAYER VI2 ;
  RECT 2123.740 3.880 2128.480 5.600 ;
  LAYER VI2 ;
  RECT 2109.800 3.880 2113.740 5.600 ;
  LAYER VI2 ;
  RECT 2102.660 3.880 2107.400 5.600 ;
  LAYER VI2 ;
  RECT 2090.200 3.880 2092.660 5.600 ;
  LAYER VI2 ;
  RECT 2082.820 3.880 2087.560 5.600 ;
  LAYER VI2 ;
  RECT 2069.000 3.880 2072.820 5.600 ;
  LAYER VI2 ;
  RECT 2061.740 3.880 2066.480 5.600 ;
  LAYER VI2 ;
  RECT 2049.000 3.880 2051.740 5.600 ;
  LAYER VI2 ;
  RECT 2041.900 3.880 2046.640 5.600 ;
  LAYER VI2 ;
  RECT 2028.200 3.880 2031.900 5.600 ;
  LAYER VI2 ;
  RECT 2020.820 3.880 2025.560 5.600 ;
  LAYER VI2 ;
  RECT 2008.200 3.880 2010.820 5.600 ;
  LAYER VI2 ;
  RECT 2000.980 3.880 2005.720 5.600 ;
  LAYER VI2 ;
  RECT 1987.000 3.880 1990.980 5.600 ;
  LAYER VI2 ;
  RECT 1979.900 3.880 1984.640 5.600 ;
  LAYER VI2 ;
  RECT 1967.400 3.880 1969.900 5.600 ;
  LAYER VI2 ;
  RECT 1960.060 3.880 1964.800 5.600 ;
  LAYER VI2 ;
  RECT 1946.200 3.880 1950.060 5.600 ;
  LAYER VI2 ;
  RECT 1938.980 3.880 1943.720 5.600 ;
  LAYER VI2 ;
  RECT 1926.200 3.880 1928.980 5.600 ;
  LAYER VI2 ;
  RECT 1919.140 3.880 1923.880 5.600 ;
  LAYER VI2 ;
  RECT 1905.400 3.880 1909.140 5.600 ;
  LAYER VI2 ;
  RECT 1898.060 3.880 1902.800 5.600 ;
  LAYER VI2 ;
  RECT 1885.400 3.880 1888.060 5.600 ;
  LAYER VI2 ;
  RECT 1878.220 3.880 1882.960 5.600 ;
  LAYER VI2 ;
  RECT 1864.200 3.880 1868.220 5.600 ;
  LAYER VI2 ;
  RECT 1857.140 3.880 1861.880 5.600 ;
  LAYER VI2 ;
  RECT 1844.600 3.880 1847.140 5.600 ;
  LAYER VI2 ;
  RECT 1837.300 3.880 1842.040 5.600 ;
  LAYER VI2 ;
  RECT 1823.400 3.880 1827.300 5.600 ;
  LAYER VI2 ;
  RECT 1816.220 3.880 1820.960 5.600 ;
  LAYER VI2 ;
  RECT 1803.800 3.880 1806.220 5.600 ;
  LAYER VI2 ;
  RECT 1796.380 3.880 1801.120 5.600 ;
  LAYER VI2 ;
  RECT 1782.600 3.880 1786.380 5.600 ;
  LAYER VI2 ;
  RECT 1775.300 3.880 1780.040 5.600 ;
  LAYER VI2 ;
  RECT 1762.600 3.880 1765.300 5.600 ;
  LAYER VI2 ;
  RECT 1755.460 3.880 1760.200 5.600 ;
  LAYER VI2 ;
  RECT 1741.800 3.880 1745.460 5.600 ;
  LAYER VI2 ;
  RECT 1734.380 3.880 1739.120 5.600 ;
  LAYER VI2 ;
  RECT 1721.800 3.880 1724.380 5.600 ;
  LAYER VI2 ;
  RECT 1714.540 3.880 1719.280 5.600 ;
  LAYER VI2 ;
  RECT 1700.600 3.880 1704.540 5.600 ;
  LAYER VI2 ;
  RECT 1693.460 3.880 1698.200 5.600 ;
  LAYER VI2 ;
  RECT 1681.000 3.880 1683.460 5.600 ;
  LAYER VI2 ;
  RECT 1673.620 3.880 1678.360 5.600 ;
  LAYER VI2 ;
  RECT 1659.800 3.880 1663.620 5.600 ;
  LAYER VI2 ;
  RECT 1652.540 3.880 1657.280 5.600 ;
  LAYER VI2 ;
  RECT 1639.800 3.880 1642.540 5.600 ;
  LAYER VI2 ;
  RECT 1632.700 3.880 1637.440 5.600 ;
  LAYER VI2 ;
  RECT 1619.000 3.880 1622.700 5.600 ;
  LAYER VI2 ;
  RECT 1611.620 3.880 1616.360 5.600 ;
  LAYER VI2 ;
  RECT 1599.000 3.880 1601.620 5.600 ;
  LAYER VI2 ;
  RECT 1591.780 3.880 1596.520 5.600 ;
  LAYER VI2 ;
  RECT 1577.800 3.880 1581.780 5.600 ;
  LAYER VI2 ;
  RECT 1570.700 3.880 1575.440 5.600 ;
  LAYER VI2 ;
  RECT 1558.200 3.880 1560.700 5.600 ;
  LAYER VI2 ;
  RECT 1550.860 3.880 1555.600 5.600 ;
  LAYER VI2 ;
  RECT 1537.000 3.880 1540.860 5.600 ;
  LAYER VI2 ;
  RECT 1529.780 3.880 1534.520 5.600 ;
  LAYER VI2 ;
  RECT 1517.000 3.880 1519.780 5.600 ;
  LAYER VI2 ;
  RECT 1509.940 3.880 1514.680 5.600 ;
  LAYER VI2 ;
  RECT 1496.200 3.880 1499.940 5.600 ;
  LAYER VI2 ;
  RECT 1488.860 3.880 1493.600 5.600 ;
  LAYER VI2 ;
  RECT 1476.200 3.880 1478.860 5.600 ;
  LAYER VI2 ;
  RECT 1469.020 3.880 1473.760 5.600 ;
  LAYER VI2 ;
  RECT 1455.000 3.880 1459.020 5.600 ;
  LAYER VI2 ;
  RECT 1447.940 3.880 1452.680 5.600 ;
  LAYER VI2 ;
  RECT 1435.400 3.880 1437.940 5.600 ;
  LAYER VI2 ;
  RECT 1428.100 3.880 1432.840 5.600 ;
  LAYER VI2 ;
  RECT 1414.200 3.880 1418.100 5.600 ;
  LAYER VI2 ;
  RECT 1407.020 3.880 1411.760 5.600 ;
  LAYER VI2 ;
  RECT 1394.600 3.880 1397.020 5.600 ;
  LAYER VI2 ;
  RECT 1387.180 3.880 1391.920 5.600 ;
  LAYER VI2 ;
  RECT 1359.210 3.880 1377.180 5.600 ;
  LAYER VI2 ;
  RECT 1347.890 3.880 1350.450 5.600 ;
  LAYER VI2 ;
  RECT 1339.800 3.880 1342.440 5.600 ;
  LAYER VI2 ;
  RECT 1313.000 3.880 1316.820 5.600 ;
  LAYER VI2 ;
  RECT 1305.720 3.880 1310.460 5.600 ;
  LAYER VI2 ;
  RECT 1293.000 3.880 1295.720 5.600 ;
  LAYER VI2 ;
  RECT 1285.880 3.880 1290.620 5.600 ;
  LAYER VI2 ;
  RECT 1272.200 3.880 1275.880 5.600 ;
  LAYER VI2 ;
  RECT 1264.800 3.880 1269.540 5.600 ;
  LAYER VI2 ;
  RECT 1252.200 3.880 1254.800 5.600 ;
  LAYER VI2 ;
  RECT 1244.960 3.880 1249.700 5.600 ;
  LAYER VI2 ;
  RECT 1231.000 3.880 1234.960 5.600 ;
  LAYER VI2 ;
  RECT 1223.880 3.880 1228.620 5.600 ;
  LAYER VI2 ;
  RECT 1211.400 3.880 1213.880 5.600 ;
  LAYER VI2 ;
  RECT 1204.040 3.880 1208.780 5.600 ;
  LAYER VI2 ;
  RECT 1190.200 3.880 1194.040 5.600 ;
  LAYER VI2 ;
  RECT 1182.960 3.880 1187.700 5.600 ;
  LAYER VI2 ;
  RECT 1170.200 3.880 1172.960 5.600 ;
  LAYER VI2 ;
  RECT 1163.120 3.880 1167.860 5.600 ;
  LAYER VI2 ;
  RECT 1149.400 3.880 1153.120 5.600 ;
  LAYER VI2 ;
  RECT 1142.040 3.880 1146.780 5.600 ;
  LAYER VI2 ;
  RECT 1129.400 3.880 1132.040 5.600 ;
  LAYER VI2 ;
  RECT 1122.200 3.880 1126.940 5.600 ;
  LAYER VI2 ;
  RECT 1108.200 3.880 1112.200 5.600 ;
  LAYER VI2 ;
  RECT 1101.120 3.880 1105.860 5.600 ;
  LAYER VI2 ;
  RECT 1088.600 3.880 1091.120 5.600 ;
  LAYER VI2 ;
  RECT 1081.280 3.880 1086.020 5.600 ;
  LAYER VI2 ;
  RECT 1067.400 3.880 1071.280 5.600 ;
  LAYER VI2 ;
  RECT 1060.200 3.880 1064.940 5.600 ;
  LAYER VI2 ;
  RECT 1047.400 3.880 1050.200 5.600 ;
  LAYER VI2 ;
  RECT 1040.360 3.880 1045.100 5.600 ;
  LAYER VI2 ;
  RECT 1026.600 3.880 1030.360 5.600 ;
  LAYER VI2 ;
  RECT 1019.280 3.880 1024.020 5.600 ;
  LAYER VI2 ;
  RECT 1006.600 3.880 1009.280 5.600 ;
  LAYER VI2 ;
  RECT 999.440 3.880 1004.180 5.600 ;
  LAYER VI2 ;
  RECT 985.400 3.880 989.440 5.600 ;
  LAYER VI2 ;
  RECT 978.360 3.880 983.100 5.600 ;
  LAYER VI2 ;
  RECT 965.800 3.880 968.360 5.600 ;
  LAYER VI2 ;
  RECT 958.520 3.880 963.260 5.600 ;
  LAYER VI2 ;
  RECT 944.600 3.880 948.520 5.600 ;
  LAYER VI2 ;
  RECT 937.440 3.880 942.180 5.600 ;
  LAYER VI2 ;
  RECT 925.000 3.880 927.440 5.600 ;
  LAYER VI2 ;
  RECT 917.600 3.880 922.340 5.600 ;
  LAYER VI2 ;
  RECT 903.800 3.880 907.600 5.600 ;
  LAYER VI2 ;
  RECT 896.520 3.880 901.260 5.600 ;
  LAYER VI2 ;
  RECT 883.800 3.880 886.520 5.600 ;
  LAYER VI2 ;
  RECT 876.680 3.880 881.420 5.600 ;
  LAYER VI2 ;
  RECT 863.000 3.880 866.680 5.600 ;
  LAYER VI2 ;
  RECT 855.600 3.880 860.340 5.600 ;
  LAYER VI2 ;
  RECT 843.000 3.880 845.600 5.600 ;
  LAYER VI2 ;
  RECT 835.760 3.880 840.500 5.600 ;
  LAYER VI2 ;
  RECT 821.800 3.880 825.760 5.600 ;
  LAYER VI2 ;
  RECT 814.680 3.880 819.420 5.600 ;
  LAYER VI2 ;
  RECT 802.200 3.880 804.680 5.600 ;
  LAYER VI2 ;
  RECT 794.840 3.880 799.580 5.600 ;
  LAYER VI2 ;
  RECT 781.000 3.880 784.840 5.600 ;
  LAYER VI2 ;
  RECT 773.760 3.880 778.500 5.600 ;
  LAYER VI2 ;
  RECT 761.000 3.880 763.760 5.600 ;
  LAYER VI2 ;
  RECT 753.920 3.880 758.660 5.600 ;
  LAYER VI2 ;
  RECT 740.200 3.880 743.920 5.600 ;
  LAYER VI2 ;
  RECT 732.840 3.880 737.580 5.600 ;
  LAYER VI2 ;
  RECT 720.200 3.880 722.840 5.600 ;
  LAYER VI2 ;
  RECT 713.000 3.880 717.740 5.600 ;
  LAYER VI2 ;
  RECT 699.000 3.880 703.000 5.600 ;
  LAYER VI2 ;
  RECT 691.920 3.880 696.660 5.600 ;
  LAYER VI2 ;
  RECT 679.400 3.880 681.920 5.600 ;
  LAYER VI2 ;
  RECT 672.080 3.880 676.820 5.600 ;
  LAYER VI2 ;
  RECT 658.200 3.880 662.080 5.600 ;
  LAYER VI2 ;
  RECT 651.000 3.880 655.740 5.600 ;
  LAYER VI2 ;
  RECT 638.200 3.880 641.000 5.600 ;
  LAYER VI2 ;
  RECT 631.160 3.880 635.900 5.600 ;
  LAYER VI2 ;
  RECT 617.400 3.880 621.160 5.600 ;
  LAYER VI2 ;
  RECT 610.080 3.880 614.820 5.600 ;
  LAYER VI2 ;
  RECT 597.400 3.880 600.080 5.600 ;
  LAYER VI2 ;
  RECT 590.240 3.880 594.980 5.600 ;
  LAYER VI2 ;
  RECT 576.200 3.880 580.240 5.600 ;
  LAYER VI2 ;
  RECT 569.160 3.880 573.900 5.600 ;
  LAYER VI2 ;
  RECT 556.600 3.880 559.160 5.600 ;
  LAYER VI2 ;
  RECT 549.320 3.880 554.060 5.600 ;
  LAYER VI2 ;
  RECT 535.400 3.880 539.320 5.600 ;
  LAYER VI2 ;
  RECT 528.240 3.880 532.980 5.600 ;
  LAYER VI2 ;
  RECT 515.800 3.880 518.240 5.600 ;
  LAYER VI2 ;
  RECT 508.400 3.880 513.140 5.600 ;
  LAYER VI2 ;
  RECT 494.600 3.880 498.400 5.600 ;
  LAYER VI2 ;
  RECT 487.320 3.880 492.060 5.600 ;
  LAYER VI2 ;
  RECT 474.600 3.880 477.320 5.600 ;
  LAYER VI2 ;
  RECT 467.480 3.880 472.220 5.600 ;
  LAYER VI2 ;
  RECT 453.800 3.880 457.480 5.600 ;
  LAYER VI2 ;
  RECT 446.400 3.880 451.140 5.600 ;
  LAYER VI2 ;
  RECT 433.800 3.880 436.400 5.600 ;
  LAYER VI2 ;
  RECT 426.560 3.880 431.300 5.600 ;
  LAYER VI2 ;
  RECT 412.600 3.880 416.560 5.600 ;
  LAYER VI2 ;
  RECT 405.480 3.880 410.220 5.600 ;
  LAYER VI2 ;
  RECT 393.000 3.880 395.480 5.600 ;
  LAYER VI2 ;
  RECT 385.640 3.880 390.380 5.600 ;
  LAYER VI2 ;
  RECT 371.800 3.880 375.640 5.600 ;
  LAYER VI2 ;
  RECT 364.560 3.880 369.300 5.600 ;
  LAYER VI2 ;
  RECT 351.800 3.880 354.560 5.600 ;
  LAYER VI2 ;
  RECT 344.720 3.880 349.460 5.600 ;
  LAYER VI2 ;
  RECT 331.000 3.880 334.720 5.600 ;
  LAYER VI2 ;
  RECT 323.640 3.880 328.380 5.600 ;
  LAYER VI2 ;
  RECT 311.000 3.880 313.640 5.600 ;
  LAYER VI2 ;
  RECT 303.800 3.880 308.540 5.600 ;
  LAYER VI2 ;
  RECT 289.800 3.880 293.800 5.600 ;
  LAYER VI2 ;
  RECT 282.720 3.880 287.460 5.600 ;
  LAYER VI2 ;
  RECT 270.200 3.880 272.720 5.600 ;
  LAYER VI2 ;
  RECT 262.880 3.880 267.620 5.600 ;
  LAYER VI2 ;
  RECT 249.000 3.880 252.880 5.600 ;
  LAYER VI2 ;
  RECT 241.800 3.880 246.540 5.600 ;
  LAYER VI2 ;
  RECT 229.000 3.880 231.800 5.600 ;
  LAYER VI2 ;
  RECT 221.960 3.880 226.700 5.600 ;
  LAYER VI2 ;
  RECT 208.200 3.880 211.960 5.600 ;
  LAYER VI2 ;
  RECT 200.880 3.880 205.620 5.600 ;
  LAYER VI2 ;
  RECT 188.200 3.880 190.880 5.600 ;
  LAYER VI2 ;
  RECT 181.040 3.880 185.780 5.600 ;
  LAYER VI2 ;
  RECT 167.000 3.880 171.040 5.600 ;
  LAYER VI2 ;
  RECT 159.960 3.880 164.700 5.600 ;
  LAYER VI2 ;
  RECT 147.400 3.880 149.960 5.600 ;
  LAYER VI2 ;
  RECT 140.120 3.880 144.860 5.600 ;
  LAYER VI2 ;
  RECT 126.200 3.880 130.120 5.600 ;
  LAYER VI2 ;
  RECT 119.040 3.880 123.780 5.600 ;
  LAYER VI2 ;
  RECT 106.600 3.880 109.040 5.600 ;
  LAYER VI2 ;
  RECT 99.200 3.880 103.940 5.600 ;
  LAYER VI2 ;
  RECT 85.400 3.880 89.200 5.600 ;
  LAYER VI2 ;
  RECT 78.120 3.880 82.860 5.600 ;
  LAYER VI2 ;
  RECT 65.400 3.880 68.120 5.600 ;
  LAYER VI2 ;
  RECT 58.280 3.880 63.020 5.600 ;
  LAYER VI2 ;
  RECT 44.600 3.880 48.280 5.600 ;
  LAYER VI2 ;
  RECT 37.200 3.880 41.940 5.600 ;
  LAYER VI2 ;
  RECT 24.600 3.880 27.200 5.600 ;
  LAYER VI2 ;
  RECT 17.360 3.880 22.100 5.600 ;
  LAYER VI1 ;
  RECT 2682.600 3.740 2688.940 5.600 ;
  LAYER VI1 ;
  RECT 2668.200 3.740 2680.280 5.600 ;
  LAYER VI1 ;
  RECT 2663.000 3.740 2665.650 5.600 ;
  LAYER VI1 ;
  RECT 2648.200 3.740 2660.440 5.600 ;
  LAYER VI1 ;
  RECT 2641.800 3.740 2645.810 5.600 ;
  LAYER VI1 ;
  RECT 2627.400 3.740 2639.360 5.600 ;
  LAYER VI1 ;
  RECT 2622.200 3.740 2624.730 5.600 ;
  LAYER VI1 ;
  RECT 2607.400 3.740 2619.520 5.600 ;
  LAYER VI1 ;
  RECT 2601.000 3.740 2604.890 5.600 ;
  LAYER VI1 ;
  RECT 2586.200 3.740 2598.440 5.600 ;
  LAYER VI1 ;
  RECT 2581.000 3.740 2583.810 5.600 ;
  LAYER VI1 ;
  RECT 2566.600 3.740 2578.600 5.600 ;
  LAYER VI1 ;
  RECT 2560.200 3.740 2563.970 5.600 ;
  LAYER VI1 ;
  RECT 2545.400 3.740 2557.520 5.600 ;
  LAYER VI1 ;
  RECT 2540.200 3.740 2542.890 5.600 ;
  LAYER VI1 ;
  RECT 2527.400 3.740 2537.680 5.600 ;
  LAYER VI1 ;
  RECT 2519.000 3.740 2523.050 5.600 ;
  LAYER VI1 ;
  RECT 2504.600 3.740 2516.600 5.600 ;
  LAYER VI1 ;
  RECT 2499.400 3.740 2501.970 5.600 ;
  LAYER VI1 ;
  RECT 2484.600 3.740 2496.760 5.600 ;
  LAYER VI1 ;
  RECT 2478.200 3.740 2482.130 5.600 ;
  LAYER VI1 ;
  RECT 2463.400 3.740 2475.680 5.600 ;
  LAYER VI1 ;
  RECT 2458.200 3.740 2461.050 5.600 ;
  LAYER VI1 ;
  RECT 2443.800 3.740 2455.840 5.600 ;
  LAYER VI1 ;
  RECT 2437.400 3.740 2441.210 5.600 ;
  LAYER VI1 ;
  RECT 2422.600 3.740 2434.760 5.600 ;
  LAYER VI1 ;
  RECT 2417.400 3.740 2420.130 5.600 ;
  LAYER VI1 ;
  RECT 2402.600 3.740 2414.920 5.600 ;
  LAYER VI1 ;
  RECT 2396.200 3.740 2400.290 5.600 ;
  LAYER VI1 ;
  RECT 2381.800 3.740 2393.840 5.600 ;
  LAYER VI1 ;
  RECT 2376.600 3.740 2379.210 5.600 ;
  LAYER VI1 ;
  RECT 2363.400 3.740 2374.000 5.600 ;
  LAYER VI1 ;
  RECT 2355.400 3.740 2359.370 5.600 ;
  LAYER VI1 ;
  RECT 2340.600 3.740 2352.920 5.600 ;
  LAYER VI1 ;
  RECT 2335.400 3.740 2338.290 5.600 ;
  LAYER VI1 ;
  RECT 2321.000 3.740 2333.080 5.600 ;
  LAYER VI1 ;
  RECT 2314.600 3.740 2318.450 5.600 ;
  LAYER VI1 ;
  RECT 2299.800 3.740 2312.000 5.600 ;
  LAYER VI1 ;
  RECT 2294.600 3.740 2297.370 5.600 ;
  LAYER VI1 ;
  RECT 2280.200 3.740 2292.160 5.600 ;
  LAYER VI1 ;
  RECT 2273.400 3.740 2277.530 5.600 ;
  LAYER VI1 ;
  RECT 2259.000 3.740 2271.080 5.600 ;
  LAYER VI1 ;
  RECT 2253.800 3.740 2256.450 5.600 ;
  LAYER VI1 ;
  RECT 2239.000 3.740 2251.240 5.600 ;
  LAYER VI1 ;
  RECT 2232.600 3.740 2236.610 5.600 ;
  LAYER VI1 ;
  RECT 2218.200 3.740 2230.160 5.600 ;
  LAYER VI1 ;
  RECT 2213.000 3.740 2215.530 5.600 ;
  LAYER VI1 ;
  RECT 2199.800 3.740 2210.320 5.600 ;
  LAYER VI1 ;
  RECT 2191.800 3.740 2195.690 5.600 ;
  LAYER VI1 ;
  RECT 2177.000 3.740 2189.240 5.600 ;
  LAYER VI1 ;
  RECT 2171.800 3.740 2174.610 5.600 ;
  LAYER VI1 ;
  RECT 2157.400 3.740 2169.400 5.600 ;
  LAYER VI1 ;
  RECT 2151.000 3.740 2154.770 5.600 ;
  LAYER VI1 ;
  RECT 2136.200 3.740 2148.320 5.600 ;
  LAYER VI1 ;
  RECT 2131.000 3.740 2133.690 5.600 ;
  LAYER VI1 ;
  RECT 2116.200 3.740 2128.480 5.600 ;
  LAYER VI1 ;
  RECT 2109.800 3.740 2113.850 5.600 ;
  LAYER VI1 ;
  RECT 2095.400 3.740 2107.400 5.600 ;
  LAYER VI1 ;
  RECT 2090.200 3.740 2092.770 5.600 ;
  LAYER VI1 ;
  RECT 2075.400 3.740 2087.560 5.600 ;
  LAYER VI1 ;
  RECT 2069.000 3.740 2072.930 5.600 ;
  LAYER VI1 ;
  RECT 2054.200 3.740 2066.480 5.600 ;
  LAYER VI1 ;
  RECT 2049.000 3.740 2051.850 5.600 ;
  LAYER VI1 ;
  RECT 2036.200 3.740 2046.640 5.600 ;
  LAYER VI1 ;
  RECT 2028.200 3.740 2032.010 5.600 ;
  LAYER VI1 ;
  RECT 2013.400 3.740 2025.560 5.600 ;
  LAYER VI1 ;
  RECT 2008.200 3.740 2010.930 5.600 ;
  LAYER VI1 ;
  RECT 1993.400 3.740 2005.720 5.600 ;
  LAYER VI1 ;
  RECT 1987.000 3.740 1991.090 5.600 ;
  LAYER VI1 ;
  RECT 1972.600 3.740 1984.640 5.600 ;
  LAYER VI1 ;
  RECT 1967.400 3.740 1970.010 5.600 ;
  LAYER VI1 ;
  RECT 1952.600 3.740 1964.800 5.600 ;
  LAYER VI1 ;
  RECT 1946.200 3.740 1950.170 5.600 ;
  LAYER VI1 ;
  RECT 1931.400 3.740 1943.720 5.600 ;
  LAYER VI1 ;
  RECT 1926.200 3.740 1929.090 5.600 ;
  LAYER VI1 ;
  RECT 1911.800 3.740 1923.880 5.600 ;
  LAYER VI1 ;
  RECT 1905.400 3.740 1909.250 5.600 ;
  LAYER VI1 ;
  RECT 1890.600 3.740 1902.800 5.600 ;
  LAYER VI1 ;
  RECT 1885.400 3.740 1888.170 5.600 ;
  LAYER VI1 ;
  RECT 1872.600 3.740 1882.960 5.600 ;
  LAYER VI1 ;
  RECT 1864.200 3.740 1868.330 5.600 ;
  LAYER VI1 ;
  RECT 1849.800 3.740 1861.880 5.600 ;
  LAYER VI1 ;
  RECT 1844.600 3.740 1847.250 5.600 ;
  LAYER VI1 ;
  RECT 1829.800 3.740 1842.040 5.600 ;
  LAYER VI1 ;
  RECT 1823.400 3.740 1827.410 5.600 ;
  LAYER VI1 ;
  RECT 1809.000 3.740 1820.960 5.600 ;
  LAYER VI1 ;
  RECT 1803.800 3.740 1806.330 5.600 ;
  LAYER VI1 ;
  RECT 1789.000 3.740 1801.120 5.600 ;
  LAYER VI1 ;
  RECT 1782.600 3.740 1786.490 5.600 ;
  LAYER VI1 ;
  RECT 1767.800 3.740 1780.040 5.600 ;
  LAYER VI1 ;
  RECT 1762.600 3.740 1765.410 5.600 ;
  LAYER VI1 ;
  RECT 1748.200 3.740 1760.200 5.600 ;
  LAYER VI1 ;
  RECT 1741.800 3.740 1745.570 5.600 ;
  LAYER VI1 ;
  RECT 1727.000 3.740 1739.120 5.600 ;
  LAYER VI1 ;
  RECT 1721.800 3.740 1724.490 5.600 ;
  LAYER VI1 ;
  RECT 1709.000 3.740 1719.280 5.600 ;
  LAYER VI1 ;
  RECT 1700.600 3.740 1704.650 5.600 ;
  LAYER VI1 ;
  RECT 1686.200 3.740 1698.200 5.600 ;
  LAYER VI1 ;
  RECT 1681.000 3.740 1683.570 5.600 ;
  LAYER VI1 ;
  RECT 1666.200 3.740 1678.360 5.600 ;
  LAYER VI1 ;
  RECT 1659.800 3.740 1663.730 5.600 ;
  LAYER VI1 ;
  RECT 1645.000 3.740 1657.280 5.600 ;
  LAYER VI1 ;
  RECT 1639.800 3.740 1642.650 5.600 ;
  LAYER VI1 ;
  RECT 1625.400 3.740 1637.440 5.600 ;
  LAYER VI1 ;
  RECT 1619.000 3.740 1622.810 5.600 ;
  LAYER VI1 ;
  RECT 1604.200 3.740 1616.360 5.600 ;
  LAYER VI1 ;
  RECT 1599.000 3.740 1601.730 5.600 ;
  LAYER VI1 ;
  RECT 1584.200 3.740 1596.520 5.600 ;
  LAYER VI1 ;
  RECT 1577.800 3.740 1581.890 5.600 ;
  LAYER VI1 ;
  RECT 1563.400 3.740 1575.440 5.600 ;
  LAYER VI1 ;
  RECT 1558.200 3.740 1560.810 5.600 ;
  LAYER VI1 ;
  RECT 1545.000 3.740 1555.600 5.600 ;
  LAYER VI1 ;
  RECT 1537.000 3.740 1540.970 5.600 ;
  LAYER VI1 ;
  RECT 1522.200 3.740 1534.520 5.600 ;
  LAYER VI1 ;
  RECT 1517.000 3.740 1519.890 5.600 ;
  LAYER VI1 ;
  RECT 1502.600 3.740 1514.680 5.600 ;
  LAYER VI1 ;
  RECT 1496.200 3.740 1500.050 5.600 ;
  LAYER VI1 ;
  RECT 1481.400 3.740 1493.600 5.600 ;
  LAYER VI1 ;
  RECT 1476.200 3.740 1478.970 5.600 ;
  LAYER VI1 ;
  RECT 1461.800 3.740 1473.760 5.600 ;
  LAYER VI1 ;
  RECT 1455.000 3.740 1459.130 5.600 ;
  LAYER VI1 ;
  RECT 1440.600 3.740 1452.680 5.600 ;
  LAYER VI1 ;
  RECT 1435.400 3.740 1438.050 5.600 ;
  LAYER VI1 ;
  RECT 1420.600 3.740 1432.840 5.600 ;
  LAYER VI1 ;
  RECT 1414.200 3.740 1418.210 5.600 ;
  LAYER VI1 ;
  RECT 1399.800 3.740 1411.760 5.600 ;
  LAYER VI1 ;
  RECT 1394.600 3.740 1397.130 5.600 ;
  LAYER VI1 ;
  RECT 1381.400 3.740 1391.920 5.600 ;
  LAYER VI1 ;
  RECT 1359.000 3.740 1377.290 5.600 ;
  LAYER VI1 ;
  RECT 1347.000 3.740 1350.450 5.600 ;
  LAYER VI1 ;
  RECT 1339.800 3.740 1344.480 5.600 ;
  LAYER VI1 ;
  RECT 1313.000 3.740 1319.840 5.600 ;
  LAYER VI1 ;
  RECT 1298.200 3.740 1310.460 5.600 ;
  LAYER VI1 ;
  RECT 1293.000 3.740 1295.830 5.600 ;
  LAYER VI1 ;
  RECT 1278.600 3.740 1290.620 5.600 ;
  LAYER VI1 ;
  RECT 1272.200 3.740 1275.990 5.600 ;
  LAYER VI1 ;
  RECT 1257.400 3.740 1269.540 5.600 ;
  LAYER VI1 ;
  RECT 1252.200 3.740 1254.910 5.600 ;
  LAYER VI1 ;
  RECT 1237.400 3.740 1249.700 5.600 ;
  LAYER VI1 ;
  RECT 1231.000 3.740 1235.070 5.600 ;
  LAYER VI1 ;
  RECT 1216.600 3.740 1228.620 5.600 ;
  LAYER VI1 ;
  RECT 1211.400 3.740 1213.990 5.600 ;
  LAYER VI1 ;
  RECT 1196.600 3.740 1208.780 5.600 ;
  LAYER VI1 ;
  RECT 1190.200 3.740 1194.150 5.600 ;
  LAYER VI1 ;
  RECT 1175.400 3.740 1187.700 5.600 ;
  LAYER VI1 ;
  RECT 1170.200 3.740 1173.070 5.600 ;
  LAYER VI1 ;
  RECT 1157.400 3.740 1167.860 5.600 ;
  LAYER VI1 ;
  RECT 1149.400 3.740 1153.230 5.600 ;
  LAYER VI1 ;
  RECT 1134.600 3.740 1146.780 5.600 ;
  LAYER VI1 ;
  RECT 1129.400 3.740 1132.150 5.600 ;
  LAYER VI1 ;
  RECT 1115.000 3.740 1126.940 5.600 ;
  LAYER VI1 ;
  RECT 1108.200 3.740 1112.310 5.600 ;
  LAYER VI1 ;
  RECT 1093.800 3.740 1105.860 5.600 ;
  LAYER VI1 ;
  RECT 1088.600 3.740 1091.230 5.600 ;
  LAYER VI1 ;
  RECT 1073.800 3.740 1086.020 5.600 ;
  LAYER VI1 ;
  RECT 1067.400 3.740 1071.390 5.600 ;
  LAYER VI1 ;
  RECT 1053.000 3.740 1064.940 5.600 ;
  LAYER VI1 ;
  RECT 1047.400 3.740 1050.310 5.600 ;
  LAYER VI1 ;
  RECT 1033.000 3.740 1045.100 5.600 ;
  LAYER VI1 ;
  RECT 1026.600 3.740 1030.470 5.600 ;
  LAYER VI1 ;
  RECT 1011.800 3.740 1024.020 5.600 ;
  LAYER VI1 ;
  RECT 1006.600 3.740 1009.390 5.600 ;
  LAYER VI1 ;
  RECT 993.800 3.740 1004.180 5.600 ;
  LAYER VI1 ;
  RECT 985.400 3.740 989.550 5.600 ;
  LAYER VI1 ;
  RECT 971.000 3.740 983.100 5.600 ;
  LAYER VI1 ;
  RECT 965.800 3.740 968.470 5.600 ;
  LAYER VI1 ;
  RECT 951.000 3.740 963.260 5.600 ;
  LAYER VI1 ;
  RECT 944.600 3.740 948.630 5.600 ;
  LAYER VI1 ;
  RECT 930.200 3.740 942.180 5.600 ;
  LAYER VI1 ;
  RECT 925.000 3.740 927.550 5.600 ;
  LAYER VI1 ;
  RECT 910.200 3.740 922.340 5.600 ;
  LAYER VI1 ;
  RECT 903.800 3.740 907.710 5.600 ;
  LAYER VI1 ;
  RECT 889.000 3.740 901.260 5.600 ;
  LAYER VI1 ;
  RECT 883.800 3.740 886.630 5.600 ;
  LAYER VI1 ;
  RECT 869.400 3.740 881.420 5.600 ;
  LAYER VI1 ;
  RECT 863.000 3.740 866.790 5.600 ;
  LAYER VI1 ;
  RECT 848.200 3.740 860.340 5.600 ;
  LAYER VI1 ;
  RECT 843.000 3.740 845.710 5.600 ;
  LAYER VI1 ;
  RECT 830.200 3.740 840.500 5.600 ;
  LAYER VI1 ;
  RECT 821.800 3.740 825.870 5.600 ;
  LAYER VI1 ;
  RECT 807.400 3.740 819.420 5.600 ;
  LAYER VI1 ;
  RECT 802.200 3.740 804.790 5.600 ;
  LAYER VI1 ;
  RECT 787.400 3.740 799.580 5.600 ;
  LAYER VI1 ;
  RECT 781.000 3.740 784.950 5.600 ;
  LAYER VI1 ;
  RECT 766.200 3.740 778.500 5.600 ;
  LAYER VI1 ;
  RECT 761.000 3.740 763.870 5.600 ;
  LAYER VI1 ;
  RECT 746.600 3.740 758.660 5.600 ;
  LAYER VI1 ;
  RECT 740.200 3.740 744.030 5.600 ;
  LAYER VI1 ;
  RECT 725.400 3.740 737.580 5.600 ;
  LAYER VI1 ;
  RECT 720.200 3.740 722.950 5.600 ;
  LAYER VI1 ;
  RECT 705.800 3.740 717.740 5.600 ;
  LAYER VI1 ;
  RECT 699.000 3.740 703.110 5.600 ;
  LAYER VI1 ;
  RECT 684.600 3.740 696.660 5.600 ;
  LAYER VI1 ;
  RECT 679.400 3.740 682.030 5.600 ;
  LAYER VI1 ;
  RECT 666.600 3.740 676.820 5.600 ;
  LAYER VI1 ;
  RECT 658.200 3.740 662.190 5.600 ;
  LAYER VI1 ;
  RECT 643.800 3.740 655.740 5.600 ;
  LAYER VI1 ;
  RECT 638.200 3.740 641.110 5.600 ;
  LAYER VI1 ;
  RECT 623.800 3.740 635.900 5.600 ;
  LAYER VI1 ;
  RECT 617.400 3.740 621.270 5.600 ;
  LAYER VI1 ;
  RECT 602.600 3.740 614.820 5.600 ;
  LAYER VI1 ;
  RECT 597.400 3.740 600.190 5.600 ;
  LAYER VI1 ;
  RECT 583.000 3.740 594.980 5.600 ;
  LAYER VI1 ;
  RECT 576.200 3.740 580.350 5.600 ;
  LAYER VI1 ;
  RECT 561.800 3.740 573.900 5.600 ;
  LAYER VI1 ;
  RECT 556.600 3.740 559.270 5.600 ;
  LAYER VI1 ;
  RECT 541.800 3.740 554.060 5.600 ;
  LAYER VI1 ;
  RECT 535.400 3.740 539.430 5.600 ;
  LAYER VI1 ;
  RECT 521.000 3.740 532.980 5.600 ;
  LAYER VI1 ;
  RECT 515.800 3.740 518.350 5.600 ;
  LAYER VI1 ;
  RECT 502.600 3.740 513.140 5.600 ;
  LAYER VI1 ;
  RECT 494.600 3.740 498.510 5.600 ;
  LAYER VI1 ;
  RECT 479.800 3.740 492.060 5.600 ;
  LAYER VI1 ;
  RECT 474.600 3.740 477.430 5.600 ;
  LAYER VI1 ;
  RECT 460.200 3.740 472.220 5.600 ;
  LAYER VI1 ;
  RECT 453.800 3.740 457.590 5.600 ;
  LAYER VI1 ;
  RECT 439.000 3.740 451.140 5.600 ;
  LAYER VI1 ;
  RECT 433.800 3.740 436.510 5.600 ;
  LAYER VI1 ;
  RECT 419.000 3.740 431.300 5.600 ;
  LAYER VI1 ;
  RECT 412.600 3.740 416.670 5.600 ;
  LAYER VI1 ;
  RECT 398.200 3.740 410.220 5.600 ;
  LAYER VI1 ;
  RECT 393.000 3.740 395.590 5.600 ;
  LAYER VI1 ;
  RECT 378.200 3.740 390.380 5.600 ;
  LAYER VI1 ;
  RECT 371.800 3.740 375.750 5.600 ;
  LAYER VI1 ;
  RECT 357.000 3.740 369.300 5.600 ;
  LAYER VI1 ;
  RECT 351.800 3.740 354.670 5.600 ;
  LAYER VI1 ;
  RECT 339.000 3.740 349.460 5.600 ;
  LAYER VI1 ;
  RECT 331.000 3.740 334.830 5.600 ;
  LAYER VI1 ;
  RECT 316.200 3.740 328.380 5.600 ;
  LAYER VI1 ;
  RECT 311.000 3.740 313.750 5.600 ;
  LAYER VI1 ;
  RECT 296.600 3.740 308.540 5.600 ;
  LAYER VI1 ;
  RECT 289.800 3.740 293.910 5.600 ;
  LAYER VI1 ;
  RECT 275.400 3.740 287.460 5.600 ;
  LAYER VI1 ;
  RECT 270.200 3.740 272.830 5.600 ;
  LAYER VI1 ;
  RECT 255.400 3.740 267.620 5.600 ;
  LAYER VI1 ;
  RECT 249.000 3.740 252.990 5.600 ;
  LAYER VI1 ;
  RECT 234.600 3.740 246.540 5.600 ;
  LAYER VI1 ;
  RECT 229.000 3.740 231.910 5.600 ;
  LAYER VI1 ;
  RECT 214.600 3.740 226.700 5.600 ;
  LAYER VI1 ;
  RECT 208.200 3.740 212.070 5.600 ;
  LAYER VI1 ;
  RECT 193.400 3.740 205.620 5.600 ;
  LAYER VI1 ;
  RECT 188.200 3.740 190.990 5.600 ;
  LAYER VI1 ;
  RECT 175.400 3.740 185.780 5.600 ;
  LAYER VI1 ;
  RECT 167.000 3.740 171.150 5.600 ;
  LAYER VI1 ;
  RECT 152.600 3.740 164.700 5.600 ;
  LAYER VI1 ;
  RECT 147.400 3.740 150.070 5.600 ;
  LAYER VI1 ;
  RECT 132.600 3.740 144.860 5.600 ;
  LAYER VI1 ;
  RECT 126.200 3.740 130.230 5.600 ;
  LAYER VI1 ;
  RECT 111.800 3.740 123.780 5.600 ;
  LAYER VI1 ;
  RECT 106.600 3.740 109.150 5.600 ;
  LAYER VI1 ;
  RECT 91.800 3.740 103.940 5.600 ;
  LAYER VI1 ;
  RECT 85.400 3.740 89.310 5.600 ;
  LAYER VI1 ;
  RECT 70.600 3.740 82.860 5.600 ;
  LAYER VI1 ;
  RECT 65.400 3.740 68.230 5.600 ;
  LAYER VI1 ;
  RECT 51.000 3.740 63.020 5.600 ;
  LAYER VI1 ;
  RECT 44.600 3.740 48.390 5.600 ;
  LAYER VI1 ;
  RECT 29.800 3.740 41.940 5.600 ;
  LAYER VI1 ;
  RECT 24.600 3.740 27.310 5.600 ;
  LAYER VI1 ;
  RECT 11.800 3.740 22.100 5.600 ;
  LAYER VI1 ;
  RECT 4.000 3.740 7.470 5.600 ;
  LAYER VI3 ;
  RECT 2.280 561.930 4.000 563.650 ;
  LAYER VI2 ;
  RECT 2.280 561.930 4.000 563.650 ;
  LAYER VI1 ;
  RECT 2.140 561.930 4.000 563.790 ;
  LAYER VI2 ;
  RECT 0.000 564.070 1.860 565.930 ;
  LAYER VI1 ;
  RECT 0.000 564.070 1.860 565.930 ;
  LAYER VI3 ;
  RECT 2688.940 3.880 2690.660 5.600 ;
  LAYER VI2 ;
  RECT 2688.940 3.880 2690.660 5.600 ;
  LAYER VI1 ;
  RECT 2688.940 3.740 2690.800 5.600 ;
  LAYER VI2 ;
  RECT 2691.080 1.600 2692.940 3.460 ;
  LAYER VI1 ;
  RECT 2691.080 1.600 2692.940 3.460 ;
  LAYER VI3 ;
  RECT 2688.940 561.930 2690.660 563.650 ;
  LAYER VI2 ;
  RECT 2688.940 561.930 2690.660 563.650 ;
  LAYER VI1 ;
  RECT 2688.940 561.930 2690.800 563.790 ;
  LAYER VI2 ;
  RECT 2691.080 564.070 2692.940 565.930 ;
  LAYER VI1 ;
  RECT 2691.080 564.070 2692.940 565.930 ;
  LAYER VI3 ;
  RECT 2.280 3.880 4.000 5.600 ;
  LAYER VI2 ;
  RECT 2.280 3.880 4.000 5.600 ;
  LAYER VI1 ;
  RECT 2.140 3.740 4.000 5.600 ;
  LAYER VI2 ;
  RECT 0.000 1.600 1.860 3.460 ;
  LAYER VI1 ;
  RECT 0.000 1.600 1.860 3.460 ;
  LAYER VI1 ;
  RECT 2680.800 0.200 2681.600 1.000 ;
  LAYER VI2 ;
  RECT 2680.800 0.200 2681.600 1.000 ;
  LAYER VI3 ;
  RECT 2680.800 0.200 2681.600 1.000 ;
  LAYER VI1 ;
  RECT 2666.400 0.200 2667.200 1.000 ;
  LAYER VI2 ;
  RECT 2666.400 0.200 2667.200 1.000 ;
  LAYER VI3 ;
  RECT 2666.400 0.200 2667.200 1.000 ;
  LAYER VI1 ;
  RECT 2661.200 0.200 2662.000 1.000 ;
  LAYER VI2 ;
  RECT 2661.200 0.200 2662.000 1.000 ;
  LAYER VI3 ;
  RECT 2661.200 0.200 2662.000 1.000 ;
  LAYER VI1 ;
  RECT 2646.400 0.200 2647.200 1.000 ;
  LAYER VI2 ;
  RECT 2646.400 0.200 2647.200 1.000 ;
  LAYER VI3 ;
  RECT 2646.400 0.200 2647.200 1.000 ;
  LAYER VI1 ;
  RECT 2640.000 0.200 2640.800 1.000 ;
  LAYER VI2 ;
  RECT 2640.000 0.200 2640.800 1.000 ;
  LAYER VI3 ;
  RECT 2640.000 0.200 2640.800 1.000 ;
  LAYER VI1 ;
  RECT 2625.600 0.200 2626.400 1.000 ;
  LAYER VI2 ;
  RECT 2625.600 0.200 2626.400 1.000 ;
  LAYER VI3 ;
  RECT 2625.600 0.200 2626.400 1.000 ;
  LAYER VI1 ;
  RECT 2620.400 0.200 2621.200 1.000 ;
  LAYER VI2 ;
  RECT 2620.400 0.200 2621.200 1.000 ;
  LAYER VI3 ;
  RECT 2620.400 0.200 2621.200 1.000 ;
  LAYER VI1 ;
  RECT 2605.600 0.200 2606.400 1.000 ;
  LAYER VI2 ;
  RECT 2605.600 0.200 2606.400 1.000 ;
  LAYER VI3 ;
  RECT 2605.600 0.200 2606.400 1.000 ;
  LAYER VI1 ;
  RECT 2599.200 0.200 2600.000 1.000 ;
  LAYER VI2 ;
  RECT 2599.200 0.200 2600.000 1.000 ;
  LAYER VI3 ;
  RECT 2599.200 0.200 2600.000 1.000 ;
  LAYER VI1 ;
  RECT 2584.400 0.200 2585.200 1.000 ;
  LAYER VI2 ;
  RECT 2584.400 0.200 2585.200 1.000 ;
  LAYER VI3 ;
  RECT 2584.400 0.200 2585.200 1.000 ;
  LAYER VI1 ;
  RECT 2579.200 0.200 2580.000 1.000 ;
  LAYER VI2 ;
  RECT 2579.200 0.200 2580.000 1.000 ;
  LAYER VI3 ;
  RECT 2579.200 0.200 2580.000 1.000 ;
  LAYER VI1 ;
  RECT 2564.800 0.200 2565.600 1.000 ;
  LAYER VI2 ;
  RECT 2564.800 0.200 2565.600 1.000 ;
  LAYER VI3 ;
  RECT 2564.800 0.200 2565.600 1.000 ;
  LAYER VI1 ;
  RECT 2558.400 0.200 2559.200 1.000 ;
  LAYER VI2 ;
  RECT 2558.400 0.200 2559.200 1.000 ;
  LAYER VI3 ;
  RECT 2558.400 0.200 2559.200 1.000 ;
  LAYER VI1 ;
  RECT 2543.600 0.200 2544.400 1.000 ;
  LAYER VI2 ;
  RECT 2543.600 0.200 2544.400 1.000 ;
  LAYER VI3 ;
  RECT 2543.600 0.200 2544.400 1.000 ;
  LAYER VI1 ;
  RECT 2538.400 0.200 2539.200 1.000 ;
  LAYER VI2 ;
  RECT 2538.400 0.200 2539.200 1.000 ;
  LAYER VI3 ;
  RECT 2538.400 0.200 2539.200 1.000 ;
  LAYER VI1 ;
  RECT 2525.600 0.200 2526.400 1.000 ;
  LAYER VI2 ;
  RECT 2525.600 0.200 2526.400 1.000 ;
  LAYER VI3 ;
  RECT 2525.600 0.200 2526.400 1.000 ;
  LAYER VI1 ;
  RECT 2523.600 0.200 2524.400 1.000 ;
  LAYER VI2 ;
  RECT 2523.600 0.200 2524.400 1.000 ;
  LAYER VI3 ;
  RECT 2523.600 0.200 2524.400 1.000 ;
  LAYER VI1 ;
  RECT 2517.200 0.200 2518.000 1.000 ;
  LAYER VI2 ;
  RECT 2517.200 0.200 2518.000 1.000 ;
  LAYER VI3 ;
  RECT 2517.200 0.200 2518.000 1.000 ;
  LAYER VI1 ;
  RECT 2502.800 0.200 2503.600 1.000 ;
  LAYER VI2 ;
  RECT 2502.800 0.200 2503.600 1.000 ;
  LAYER VI3 ;
  RECT 2502.800 0.200 2503.600 1.000 ;
  LAYER VI1 ;
  RECT 2497.600 0.200 2498.400 1.000 ;
  LAYER VI2 ;
  RECT 2497.600 0.200 2498.400 1.000 ;
  LAYER VI3 ;
  RECT 2497.600 0.200 2498.400 1.000 ;
  LAYER VI1 ;
  RECT 2482.800 0.200 2483.600 1.000 ;
  LAYER VI2 ;
  RECT 2482.800 0.200 2483.600 1.000 ;
  LAYER VI3 ;
  RECT 2482.800 0.200 2483.600 1.000 ;
  LAYER VI1 ;
  RECT 2476.400 0.200 2477.200 1.000 ;
  LAYER VI2 ;
  RECT 2476.400 0.200 2477.200 1.000 ;
  LAYER VI3 ;
  RECT 2476.400 0.200 2477.200 1.000 ;
  LAYER VI1 ;
  RECT 2461.600 0.200 2462.400 1.000 ;
  LAYER VI2 ;
  RECT 2461.600 0.200 2462.400 1.000 ;
  LAYER VI3 ;
  RECT 2461.600 0.200 2462.400 1.000 ;
  LAYER VI1 ;
  RECT 2456.400 0.200 2457.200 1.000 ;
  LAYER VI2 ;
  RECT 2456.400 0.200 2457.200 1.000 ;
  LAYER VI3 ;
  RECT 2456.400 0.200 2457.200 1.000 ;
  LAYER VI1 ;
  RECT 2442.000 0.200 2442.800 1.000 ;
  LAYER VI2 ;
  RECT 2442.000 0.200 2442.800 1.000 ;
  LAYER VI3 ;
  RECT 2442.000 0.200 2442.800 1.000 ;
  LAYER VI1 ;
  RECT 2435.600 0.200 2436.400 1.000 ;
  LAYER VI2 ;
  RECT 2435.600 0.200 2436.400 1.000 ;
  LAYER VI3 ;
  RECT 2435.600 0.200 2436.400 1.000 ;
  LAYER VI1 ;
  RECT 2420.800 0.200 2421.600 1.000 ;
  LAYER VI2 ;
  RECT 2420.800 0.200 2421.600 1.000 ;
  LAYER VI3 ;
  RECT 2420.800 0.200 2421.600 1.000 ;
  LAYER VI1 ;
  RECT 2415.600 0.200 2416.400 1.000 ;
  LAYER VI2 ;
  RECT 2415.600 0.200 2416.400 1.000 ;
  LAYER VI3 ;
  RECT 2415.600 0.200 2416.400 1.000 ;
  LAYER VI1 ;
  RECT 2400.800 0.200 2401.600 1.000 ;
  LAYER VI2 ;
  RECT 2400.800 0.200 2401.600 1.000 ;
  LAYER VI3 ;
  RECT 2400.800 0.200 2401.600 1.000 ;
  LAYER VI1 ;
  RECT 2394.400 0.200 2395.200 1.000 ;
  LAYER VI2 ;
  RECT 2394.400 0.200 2395.200 1.000 ;
  LAYER VI3 ;
  RECT 2394.400 0.200 2395.200 1.000 ;
  LAYER VI1 ;
  RECT 2380.000 0.200 2380.800 1.000 ;
  LAYER VI2 ;
  RECT 2380.000 0.200 2380.800 1.000 ;
  LAYER VI3 ;
  RECT 2380.000 0.200 2380.800 1.000 ;
  LAYER VI1 ;
  RECT 2374.800 0.200 2375.600 1.000 ;
  LAYER VI2 ;
  RECT 2374.800 0.200 2375.600 1.000 ;
  LAYER VI3 ;
  RECT 2374.800 0.200 2375.600 1.000 ;
  LAYER VI1 ;
  RECT 2361.600 0.200 2362.400 1.000 ;
  LAYER VI2 ;
  RECT 2361.600 0.200 2362.400 1.000 ;
  LAYER VI3 ;
  RECT 2361.600 0.200 2362.400 1.000 ;
  LAYER VI1 ;
  RECT 2360.000 0.200 2360.800 1.000 ;
  LAYER VI2 ;
  RECT 2360.000 0.200 2360.800 1.000 ;
  LAYER VI3 ;
  RECT 2360.000 0.200 2360.800 1.000 ;
  LAYER VI1 ;
  RECT 2353.600 0.200 2354.400 1.000 ;
  LAYER VI2 ;
  RECT 2353.600 0.200 2354.400 1.000 ;
  LAYER VI3 ;
  RECT 2353.600 0.200 2354.400 1.000 ;
  LAYER VI1 ;
  RECT 2338.800 0.200 2339.600 1.000 ;
  LAYER VI2 ;
  RECT 2338.800 0.200 2339.600 1.000 ;
  LAYER VI3 ;
  RECT 2338.800 0.200 2339.600 1.000 ;
  LAYER VI1 ;
  RECT 2333.600 0.200 2334.400 1.000 ;
  LAYER VI2 ;
  RECT 2333.600 0.200 2334.400 1.000 ;
  LAYER VI3 ;
  RECT 2333.600 0.200 2334.400 1.000 ;
  LAYER VI1 ;
  RECT 2319.200 0.200 2320.000 1.000 ;
  LAYER VI2 ;
  RECT 2319.200 0.200 2320.000 1.000 ;
  LAYER VI3 ;
  RECT 2319.200 0.200 2320.000 1.000 ;
  LAYER VI1 ;
  RECT 2312.800 0.200 2313.600 1.000 ;
  LAYER VI2 ;
  RECT 2312.800 0.200 2313.600 1.000 ;
  LAYER VI3 ;
  RECT 2312.800 0.200 2313.600 1.000 ;
  LAYER VI1 ;
  RECT 2298.000 0.200 2298.800 1.000 ;
  LAYER VI2 ;
  RECT 2298.000 0.200 2298.800 1.000 ;
  LAYER VI3 ;
  RECT 2298.000 0.200 2298.800 1.000 ;
  LAYER VI1 ;
  RECT 2292.800 0.200 2293.600 1.000 ;
  LAYER VI2 ;
  RECT 2292.800 0.200 2293.600 1.000 ;
  LAYER VI3 ;
  RECT 2292.800 0.200 2293.600 1.000 ;
  LAYER VI1 ;
  RECT 2278.400 0.200 2279.200 1.000 ;
  LAYER VI2 ;
  RECT 2278.400 0.200 2279.200 1.000 ;
  LAYER VI3 ;
  RECT 2278.400 0.200 2279.200 1.000 ;
  LAYER VI1 ;
  RECT 2271.600 0.200 2272.400 1.000 ;
  LAYER VI2 ;
  RECT 2271.600 0.200 2272.400 1.000 ;
  LAYER VI3 ;
  RECT 2271.600 0.200 2272.400 1.000 ;
  LAYER VI1 ;
  RECT 2257.200 0.200 2258.000 1.000 ;
  LAYER VI2 ;
  RECT 2257.200 0.200 2258.000 1.000 ;
  LAYER VI3 ;
  RECT 2257.200 0.200 2258.000 1.000 ;
  LAYER VI1 ;
  RECT 2252.000 0.200 2252.800 1.000 ;
  LAYER VI2 ;
  RECT 2252.000 0.200 2252.800 1.000 ;
  LAYER VI3 ;
  RECT 2252.000 0.200 2252.800 1.000 ;
  LAYER VI1 ;
  RECT 2237.200 0.200 2238.000 1.000 ;
  LAYER VI2 ;
  RECT 2237.200 0.200 2238.000 1.000 ;
  LAYER VI3 ;
  RECT 2237.200 0.200 2238.000 1.000 ;
  LAYER VI1 ;
  RECT 2230.800 0.200 2231.600 1.000 ;
  LAYER VI2 ;
  RECT 2230.800 0.200 2231.600 1.000 ;
  LAYER VI3 ;
  RECT 2230.800 0.200 2231.600 1.000 ;
  LAYER VI1 ;
  RECT 2216.400 0.200 2217.200 1.000 ;
  LAYER VI2 ;
  RECT 2216.400 0.200 2217.200 1.000 ;
  LAYER VI3 ;
  RECT 2216.400 0.200 2217.200 1.000 ;
  LAYER VI1 ;
  RECT 2211.200 0.200 2212.000 1.000 ;
  LAYER VI2 ;
  RECT 2211.200 0.200 2212.000 1.000 ;
  LAYER VI3 ;
  RECT 2211.200 0.200 2212.000 1.000 ;
  LAYER VI1 ;
  RECT 2198.000 0.200 2198.800 1.000 ;
  LAYER VI2 ;
  RECT 2198.000 0.200 2198.800 1.000 ;
  LAYER VI3 ;
  RECT 2198.000 0.200 2198.800 1.000 ;
  LAYER VI1 ;
  RECT 2196.400 0.200 2197.200 1.000 ;
  LAYER VI2 ;
  RECT 2196.400 0.200 2197.200 1.000 ;
  LAYER VI3 ;
  RECT 2196.400 0.200 2197.200 1.000 ;
  LAYER VI1 ;
  RECT 2190.000 0.200 2190.800 1.000 ;
  LAYER VI2 ;
  RECT 2190.000 0.200 2190.800 1.000 ;
  LAYER VI3 ;
  RECT 2190.000 0.200 2190.800 1.000 ;
  LAYER VI1 ;
  RECT 2175.200 0.200 2176.000 1.000 ;
  LAYER VI2 ;
  RECT 2175.200 0.200 2176.000 1.000 ;
  LAYER VI3 ;
  RECT 2175.200 0.200 2176.000 1.000 ;
  LAYER VI1 ;
  RECT 2170.000 0.200 2170.800 1.000 ;
  LAYER VI2 ;
  RECT 2170.000 0.200 2170.800 1.000 ;
  LAYER VI3 ;
  RECT 2170.000 0.200 2170.800 1.000 ;
  LAYER VI1 ;
  RECT 2155.600 0.200 2156.400 1.000 ;
  LAYER VI2 ;
  RECT 2155.600 0.200 2156.400 1.000 ;
  LAYER VI3 ;
  RECT 2155.600 0.200 2156.400 1.000 ;
  LAYER VI1 ;
  RECT 2149.200 0.200 2150.000 1.000 ;
  LAYER VI2 ;
  RECT 2149.200 0.200 2150.000 1.000 ;
  LAYER VI3 ;
  RECT 2149.200 0.200 2150.000 1.000 ;
  LAYER VI1 ;
  RECT 2134.400 0.200 2135.200 1.000 ;
  LAYER VI2 ;
  RECT 2134.400 0.200 2135.200 1.000 ;
  LAYER VI3 ;
  RECT 2134.400 0.200 2135.200 1.000 ;
  LAYER VI1 ;
  RECT 2129.200 0.200 2130.000 1.000 ;
  LAYER VI2 ;
  RECT 2129.200 0.200 2130.000 1.000 ;
  LAYER VI3 ;
  RECT 2129.200 0.200 2130.000 1.000 ;
  LAYER VI1 ;
  RECT 2114.400 0.200 2115.200 1.000 ;
  LAYER VI2 ;
  RECT 2114.400 0.200 2115.200 1.000 ;
  LAYER VI3 ;
  RECT 2114.400 0.200 2115.200 1.000 ;
  LAYER VI1 ;
  RECT 2108.000 0.200 2108.800 1.000 ;
  LAYER VI2 ;
  RECT 2108.000 0.200 2108.800 1.000 ;
  LAYER VI3 ;
  RECT 2108.000 0.200 2108.800 1.000 ;
  LAYER VI1 ;
  RECT 2093.600 0.200 2094.400 1.000 ;
  LAYER VI2 ;
  RECT 2093.600 0.200 2094.400 1.000 ;
  LAYER VI3 ;
  RECT 2093.600 0.200 2094.400 1.000 ;
  LAYER VI1 ;
  RECT 2088.400 0.200 2089.200 1.000 ;
  LAYER VI2 ;
  RECT 2088.400 0.200 2089.200 1.000 ;
  LAYER VI3 ;
  RECT 2088.400 0.200 2089.200 1.000 ;
  LAYER VI1 ;
  RECT 2073.600 0.200 2074.400 1.000 ;
  LAYER VI2 ;
  RECT 2073.600 0.200 2074.400 1.000 ;
  LAYER VI3 ;
  RECT 2073.600 0.200 2074.400 1.000 ;
  LAYER VI1 ;
  RECT 2067.200 0.200 2068.000 1.000 ;
  LAYER VI2 ;
  RECT 2067.200 0.200 2068.000 1.000 ;
  LAYER VI3 ;
  RECT 2067.200 0.200 2068.000 1.000 ;
  LAYER VI1 ;
  RECT 2052.400 0.200 2053.200 1.000 ;
  LAYER VI2 ;
  RECT 2052.400 0.200 2053.200 1.000 ;
  LAYER VI3 ;
  RECT 2052.400 0.200 2053.200 1.000 ;
  LAYER VI1 ;
  RECT 2047.200 0.200 2048.000 1.000 ;
  LAYER VI2 ;
  RECT 2047.200 0.200 2048.000 1.000 ;
  LAYER VI3 ;
  RECT 2047.200 0.200 2048.000 1.000 ;
  LAYER VI1 ;
  RECT 2034.400 0.200 2035.200 1.000 ;
  LAYER VI2 ;
  RECT 2034.400 0.200 2035.200 1.000 ;
  LAYER VI3 ;
  RECT 2034.400 0.200 2035.200 1.000 ;
  LAYER VI1 ;
  RECT 2032.800 0.200 2033.600 1.000 ;
  LAYER VI2 ;
  RECT 2032.800 0.200 2033.600 1.000 ;
  LAYER VI3 ;
  RECT 2032.800 0.200 2033.600 1.000 ;
  LAYER VI1 ;
  RECT 2026.400 0.200 2027.200 1.000 ;
  LAYER VI2 ;
  RECT 2026.400 0.200 2027.200 1.000 ;
  LAYER VI3 ;
  RECT 2026.400 0.200 2027.200 1.000 ;
  LAYER VI1 ;
  RECT 2011.600 0.200 2012.400 1.000 ;
  LAYER VI2 ;
  RECT 2011.600 0.200 2012.400 1.000 ;
  LAYER VI3 ;
  RECT 2011.600 0.200 2012.400 1.000 ;
  LAYER VI1 ;
  RECT 2006.400 0.200 2007.200 1.000 ;
  LAYER VI2 ;
  RECT 2006.400 0.200 2007.200 1.000 ;
  LAYER VI3 ;
  RECT 2006.400 0.200 2007.200 1.000 ;
  LAYER VI1 ;
  RECT 1991.600 0.200 1992.400 1.000 ;
  LAYER VI2 ;
  RECT 1991.600 0.200 1992.400 1.000 ;
  LAYER VI3 ;
  RECT 1991.600 0.200 1992.400 1.000 ;
  LAYER VI1 ;
  RECT 1985.200 0.200 1986.000 1.000 ;
  LAYER VI2 ;
  RECT 1985.200 0.200 1986.000 1.000 ;
  LAYER VI3 ;
  RECT 1985.200 0.200 1986.000 1.000 ;
  LAYER VI1 ;
  RECT 1970.800 0.200 1971.600 1.000 ;
  LAYER VI2 ;
  RECT 1970.800 0.200 1971.600 1.000 ;
  LAYER VI3 ;
  RECT 1970.800 0.200 1971.600 1.000 ;
  LAYER VI1 ;
  RECT 1965.600 0.200 1966.400 1.000 ;
  LAYER VI2 ;
  RECT 1965.600 0.200 1966.400 1.000 ;
  LAYER VI3 ;
  RECT 1965.600 0.200 1966.400 1.000 ;
  LAYER VI1 ;
  RECT 1950.800 0.200 1951.600 1.000 ;
  LAYER VI2 ;
  RECT 1950.800 0.200 1951.600 1.000 ;
  LAYER VI3 ;
  RECT 1950.800 0.200 1951.600 1.000 ;
  LAYER VI1 ;
  RECT 1944.400 0.200 1945.200 1.000 ;
  LAYER VI2 ;
  RECT 1944.400 0.200 1945.200 1.000 ;
  LAYER VI3 ;
  RECT 1944.400 0.200 1945.200 1.000 ;
  LAYER VI1 ;
  RECT 1929.600 0.200 1930.400 1.000 ;
  LAYER VI2 ;
  RECT 1929.600 0.200 1930.400 1.000 ;
  LAYER VI3 ;
  RECT 1929.600 0.200 1930.400 1.000 ;
  LAYER VI1 ;
  RECT 1924.400 0.200 1925.200 1.000 ;
  LAYER VI2 ;
  RECT 1924.400 0.200 1925.200 1.000 ;
  LAYER VI3 ;
  RECT 1924.400 0.200 1925.200 1.000 ;
  LAYER VI1 ;
  RECT 1910.000 0.200 1910.800 1.000 ;
  LAYER VI2 ;
  RECT 1910.000 0.200 1910.800 1.000 ;
  LAYER VI3 ;
  RECT 1910.000 0.200 1910.800 1.000 ;
  LAYER VI1 ;
  RECT 1903.600 0.200 1904.400 1.000 ;
  LAYER VI2 ;
  RECT 1903.600 0.200 1904.400 1.000 ;
  LAYER VI3 ;
  RECT 1903.600 0.200 1904.400 1.000 ;
  LAYER VI1 ;
  RECT 1888.800 0.200 1889.600 1.000 ;
  LAYER VI2 ;
  RECT 1888.800 0.200 1889.600 1.000 ;
  LAYER VI3 ;
  RECT 1888.800 0.200 1889.600 1.000 ;
  LAYER VI1 ;
  RECT 1883.600 0.200 1884.400 1.000 ;
  LAYER VI2 ;
  RECT 1883.600 0.200 1884.400 1.000 ;
  LAYER VI3 ;
  RECT 1883.600 0.200 1884.400 1.000 ;
  LAYER VI1 ;
  RECT 1870.800 0.200 1871.600 1.000 ;
  LAYER VI2 ;
  RECT 1870.800 0.200 1871.600 1.000 ;
  LAYER VI3 ;
  RECT 1870.800 0.200 1871.600 1.000 ;
  LAYER VI1 ;
  RECT 1869.200 0.200 1870.000 1.000 ;
  LAYER VI2 ;
  RECT 1869.200 0.200 1870.000 1.000 ;
  LAYER VI3 ;
  RECT 1869.200 0.200 1870.000 1.000 ;
  LAYER VI1 ;
  RECT 1862.400 0.200 1863.200 1.000 ;
  LAYER VI2 ;
  RECT 1862.400 0.200 1863.200 1.000 ;
  LAYER VI3 ;
  RECT 1862.400 0.200 1863.200 1.000 ;
  LAYER VI1 ;
  RECT 1848.000 0.200 1848.800 1.000 ;
  LAYER VI2 ;
  RECT 1848.000 0.200 1848.800 1.000 ;
  LAYER VI3 ;
  RECT 1848.000 0.200 1848.800 1.000 ;
  LAYER VI1 ;
  RECT 1842.800 0.200 1843.600 1.000 ;
  LAYER VI2 ;
  RECT 1842.800 0.200 1843.600 1.000 ;
  LAYER VI3 ;
  RECT 1842.800 0.200 1843.600 1.000 ;
  LAYER VI1 ;
  RECT 1828.000 0.200 1828.800 1.000 ;
  LAYER VI2 ;
  RECT 1828.000 0.200 1828.800 1.000 ;
  LAYER VI3 ;
  RECT 1828.000 0.200 1828.800 1.000 ;
  LAYER VI1 ;
  RECT 1821.600 0.200 1822.400 1.000 ;
  LAYER VI2 ;
  RECT 1821.600 0.200 1822.400 1.000 ;
  LAYER VI3 ;
  RECT 1821.600 0.200 1822.400 1.000 ;
  LAYER VI1 ;
  RECT 1807.200 0.200 1808.000 1.000 ;
  LAYER VI2 ;
  RECT 1807.200 0.200 1808.000 1.000 ;
  LAYER VI3 ;
  RECT 1807.200 0.200 1808.000 1.000 ;
  LAYER VI1 ;
  RECT 1802.000 0.200 1802.800 1.000 ;
  LAYER VI2 ;
  RECT 1802.000 0.200 1802.800 1.000 ;
  LAYER VI3 ;
  RECT 1802.000 0.200 1802.800 1.000 ;
  LAYER VI1 ;
  RECT 1787.200 0.200 1788.000 1.000 ;
  LAYER VI2 ;
  RECT 1787.200 0.200 1788.000 1.000 ;
  LAYER VI3 ;
  RECT 1787.200 0.200 1788.000 1.000 ;
  LAYER VI1 ;
  RECT 1780.800 0.200 1781.600 1.000 ;
  LAYER VI2 ;
  RECT 1780.800 0.200 1781.600 1.000 ;
  LAYER VI3 ;
  RECT 1780.800 0.200 1781.600 1.000 ;
  LAYER VI1 ;
  RECT 1766.000 0.200 1766.800 1.000 ;
  LAYER VI2 ;
  RECT 1766.000 0.200 1766.800 1.000 ;
  LAYER VI3 ;
  RECT 1766.000 0.200 1766.800 1.000 ;
  LAYER VI1 ;
  RECT 1760.800 0.200 1761.600 1.000 ;
  LAYER VI2 ;
  RECT 1760.800 0.200 1761.600 1.000 ;
  LAYER VI3 ;
  RECT 1760.800 0.200 1761.600 1.000 ;
  LAYER VI1 ;
  RECT 1746.400 0.200 1747.200 1.000 ;
  LAYER VI2 ;
  RECT 1746.400 0.200 1747.200 1.000 ;
  LAYER VI3 ;
  RECT 1746.400 0.200 1747.200 1.000 ;
  LAYER VI1 ;
  RECT 1740.000 0.200 1740.800 1.000 ;
  LAYER VI2 ;
  RECT 1740.000 0.200 1740.800 1.000 ;
  LAYER VI3 ;
  RECT 1740.000 0.200 1740.800 1.000 ;
  LAYER VI1 ;
  RECT 1725.200 0.200 1726.000 1.000 ;
  LAYER VI2 ;
  RECT 1725.200 0.200 1726.000 1.000 ;
  LAYER VI3 ;
  RECT 1725.200 0.200 1726.000 1.000 ;
  LAYER VI1 ;
  RECT 1720.000 0.200 1720.800 1.000 ;
  LAYER VI2 ;
  RECT 1720.000 0.200 1720.800 1.000 ;
  LAYER VI3 ;
  RECT 1720.000 0.200 1720.800 1.000 ;
  LAYER VI1 ;
  RECT 1707.200 0.200 1708.000 1.000 ;
  LAYER VI2 ;
  RECT 1707.200 0.200 1708.000 1.000 ;
  LAYER VI3 ;
  RECT 1707.200 0.200 1708.000 1.000 ;
  LAYER VI1 ;
  RECT 1705.200 0.200 1706.000 1.000 ;
  LAYER VI2 ;
  RECT 1705.200 0.200 1706.000 1.000 ;
  LAYER VI3 ;
  RECT 1705.200 0.200 1706.000 1.000 ;
  LAYER VI1 ;
  RECT 1698.800 0.200 1699.600 1.000 ;
  LAYER VI2 ;
  RECT 1698.800 0.200 1699.600 1.000 ;
  LAYER VI3 ;
  RECT 1698.800 0.200 1699.600 1.000 ;
  LAYER VI1 ;
  RECT 1684.400 0.200 1685.200 1.000 ;
  LAYER VI2 ;
  RECT 1684.400 0.200 1685.200 1.000 ;
  LAYER VI3 ;
  RECT 1684.400 0.200 1685.200 1.000 ;
  LAYER VI1 ;
  RECT 1679.200 0.200 1680.000 1.000 ;
  LAYER VI2 ;
  RECT 1679.200 0.200 1680.000 1.000 ;
  LAYER VI3 ;
  RECT 1679.200 0.200 1680.000 1.000 ;
  LAYER VI1 ;
  RECT 1664.400 0.200 1665.200 1.000 ;
  LAYER VI2 ;
  RECT 1664.400 0.200 1665.200 1.000 ;
  LAYER VI3 ;
  RECT 1664.400 0.200 1665.200 1.000 ;
  LAYER VI1 ;
  RECT 1658.000 0.200 1658.800 1.000 ;
  LAYER VI2 ;
  RECT 1658.000 0.200 1658.800 1.000 ;
  LAYER VI3 ;
  RECT 1658.000 0.200 1658.800 1.000 ;
  LAYER VI1 ;
  RECT 1643.200 0.200 1644.000 1.000 ;
  LAYER VI2 ;
  RECT 1643.200 0.200 1644.000 1.000 ;
  LAYER VI3 ;
  RECT 1643.200 0.200 1644.000 1.000 ;
  LAYER VI1 ;
  RECT 1638.000 0.200 1638.800 1.000 ;
  LAYER VI2 ;
  RECT 1638.000 0.200 1638.800 1.000 ;
  LAYER VI3 ;
  RECT 1638.000 0.200 1638.800 1.000 ;
  LAYER VI1 ;
  RECT 1623.600 0.200 1624.400 1.000 ;
  LAYER VI2 ;
  RECT 1623.600 0.200 1624.400 1.000 ;
  LAYER VI3 ;
  RECT 1623.600 0.200 1624.400 1.000 ;
  LAYER VI1 ;
  RECT 1617.200 0.200 1618.000 1.000 ;
  LAYER VI2 ;
  RECT 1617.200 0.200 1618.000 1.000 ;
  LAYER VI3 ;
  RECT 1617.200 0.200 1618.000 1.000 ;
  LAYER VI1 ;
  RECT 1602.400 0.200 1603.200 1.000 ;
  LAYER VI2 ;
  RECT 1602.400 0.200 1603.200 1.000 ;
  LAYER VI3 ;
  RECT 1602.400 0.200 1603.200 1.000 ;
  LAYER VI1 ;
  RECT 1597.200 0.200 1598.000 1.000 ;
  LAYER VI2 ;
  RECT 1597.200 0.200 1598.000 1.000 ;
  LAYER VI3 ;
  RECT 1597.200 0.200 1598.000 1.000 ;
  LAYER VI1 ;
  RECT 1582.400 0.200 1583.200 1.000 ;
  LAYER VI2 ;
  RECT 1582.400 0.200 1583.200 1.000 ;
  LAYER VI3 ;
  RECT 1582.400 0.200 1583.200 1.000 ;
  LAYER VI1 ;
  RECT 1576.000 0.200 1576.800 1.000 ;
  LAYER VI2 ;
  RECT 1576.000 0.200 1576.800 1.000 ;
  LAYER VI3 ;
  RECT 1576.000 0.200 1576.800 1.000 ;
  LAYER VI1 ;
  RECT 1561.600 0.200 1562.400 1.000 ;
  LAYER VI2 ;
  RECT 1561.600 0.200 1562.400 1.000 ;
  LAYER VI3 ;
  RECT 1561.600 0.200 1562.400 1.000 ;
  LAYER VI1 ;
  RECT 1556.400 0.200 1557.200 1.000 ;
  LAYER VI2 ;
  RECT 1556.400 0.200 1557.200 1.000 ;
  LAYER VI3 ;
  RECT 1556.400 0.200 1557.200 1.000 ;
  LAYER VI1 ;
  RECT 1543.200 0.200 1544.000 1.000 ;
  LAYER VI2 ;
  RECT 1543.200 0.200 1544.000 1.000 ;
  LAYER VI3 ;
  RECT 1543.200 0.200 1544.000 1.000 ;
  LAYER VI1 ;
  RECT 1541.600 0.200 1542.400 1.000 ;
  LAYER VI2 ;
  RECT 1541.600 0.200 1542.400 1.000 ;
  LAYER VI3 ;
  RECT 1541.600 0.200 1542.400 1.000 ;
  LAYER VI1 ;
  RECT 1535.200 0.200 1536.000 1.000 ;
  LAYER VI2 ;
  RECT 1535.200 0.200 1536.000 1.000 ;
  LAYER VI3 ;
  RECT 1535.200 0.200 1536.000 1.000 ;
  LAYER VI1 ;
  RECT 1520.400 0.200 1521.200 1.000 ;
  LAYER VI2 ;
  RECT 1520.400 0.200 1521.200 1.000 ;
  LAYER VI3 ;
  RECT 1520.400 0.200 1521.200 1.000 ;
  LAYER VI1 ;
  RECT 1515.200 0.200 1516.000 1.000 ;
  LAYER VI2 ;
  RECT 1515.200 0.200 1516.000 1.000 ;
  LAYER VI3 ;
  RECT 1515.200 0.200 1516.000 1.000 ;
  LAYER VI1 ;
  RECT 1500.800 0.200 1501.600 1.000 ;
  LAYER VI2 ;
  RECT 1500.800 0.200 1501.600 1.000 ;
  LAYER VI3 ;
  RECT 1500.800 0.200 1501.600 1.000 ;
  LAYER VI1 ;
  RECT 1494.400 0.200 1495.200 1.000 ;
  LAYER VI2 ;
  RECT 1494.400 0.200 1495.200 1.000 ;
  LAYER VI3 ;
  RECT 1494.400 0.200 1495.200 1.000 ;
  LAYER VI1 ;
  RECT 1479.600 0.200 1480.400 1.000 ;
  LAYER VI2 ;
  RECT 1479.600 0.200 1480.400 1.000 ;
  LAYER VI3 ;
  RECT 1479.600 0.200 1480.400 1.000 ;
  LAYER VI1 ;
  RECT 1474.400 0.200 1475.200 1.000 ;
  LAYER VI2 ;
  RECT 1474.400 0.200 1475.200 1.000 ;
  LAYER VI3 ;
  RECT 1474.400 0.200 1475.200 1.000 ;
  LAYER VI1 ;
  RECT 1460.000 0.200 1460.800 1.000 ;
  LAYER VI2 ;
  RECT 1460.000 0.200 1460.800 1.000 ;
  LAYER VI3 ;
  RECT 1460.000 0.200 1460.800 1.000 ;
  LAYER VI1 ;
  RECT 1453.200 0.200 1454.000 1.000 ;
  LAYER VI2 ;
  RECT 1453.200 0.200 1454.000 1.000 ;
  LAYER VI3 ;
  RECT 1453.200 0.200 1454.000 1.000 ;
  LAYER VI1 ;
  RECT 1438.800 0.200 1439.600 1.000 ;
  LAYER VI2 ;
  RECT 1438.800 0.200 1439.600 1.000 ;
  LAYER VI3 ;
  RECT 1438.800 0.200 1439.600 1.000 ;
  LAYER VI1 ;
  RECT 1433.600 0.200 1434.400 1.000 ;
  LAYER VI2 ;
  RECT 1433.600 0.200 1434.400 1.000 ;
  LAYER VI3 ;
  RECT 1433.600 0.200 1434.400 1.000 ;
  LAYER VI1 ;
  RECT 1418.800 0.200 1419.600 1.000 ;
  LAYER VI2 ;
  RECT 1418.800 0.200 1419.600 1.000 ;
  LAYER VI3 ;
  RECT 1418.800 0.200 1419.600 1.000 ;
  LAYER VI1 ;
  RECT 1412.400 0.200 1413.200 1.000 ;
  LAYER VI2 ;
  RECT 1412.400 0.200 1413.200 1.000 ;
  LAYER VI3 ;
  RECT 1412.400 0.200 1413.200 1.000 ;
  LAYER VI1 ;
  RECT 1398.000 0.200 1398.800 1.000 ;
  LAYER VI2 ;
  RECT 1398.000 0.200 1398.800 1.000 ;
  LAYER VI3 ;
  RECT 1398.000 0.200 1398.800 1.000 ;
  LAYER VI1 ;
  RECT 1392.800 0.200 1393.600 1.000 ;
  LAYER VI2 ;
  RECT 1392.800 0.200 1393.600 1.000 ;
  LAYER VI3 ;
  RECT 1392.800 0.200 1393.600 1.000 ;
  LAYER VI1 ;
  RECT 1379.600 0.200 1380.400 1.000 ;
  LAYER VI2 ;
  RECT 1379.600 0.200 1380.400 1.000 ;
  LAYER VI3 ;
  RECT 1379.600 0.200 1380.400 1.000 ;
  LAYER VI1 ;
  RECT 1378.000 0.200 1378.800 1.000 ;
  LAYER VI2 ;
  RECT 1378.000 0.200 1378.800 1.000 ;
  LAYER VI3 ;
  RECT 1378.000 0.200 1378.800 1.000 ;
  LAYER VI1 ;
  RECT 1357.200 0.200 1358.000 1.000 ;
  LAYER VI2 ;
  RECT 1357.200 0.200 1358.000 1.000 ;
  LAYER VI3 ;
  RECT 1357.200 0.200 1358.000 1.000 ;
  LAYER VI1 ;
  RECT 1356.000 0.200 1356.800 1.000 ;
  LAYER VI2 ;
  RECT 1356.000 0.200 1356.800 1.000 ;
  LAYER VI3 ;
  RECT 1356.000 0.200 1356.800 1.000 ;
  LAYER VI1 ;
  RECT 1354.800 0.200 1355.600 1.000 ;
  LAYER VI2 ;
  RECT 1354.800 0.200 1355.600 1.000 ;
  LAYER VI3 ;
  RECT 1354.800 0.200 1355.600 1.000 ;
  LAYER VI1 ;
  RECT 1353.600 0.200 1354.400 1.000 ;
  LAYER VI2 ;
  RECT 1353.600 0.200 1354.400 1.000 ;
  LAYER VI3 ;
  RECT 1353.600 0.200 1354.400 1.000 ;
  LAYER VI1 ;
  RECT 1352.400 0.200 1353.200 1.000 ;
  LAYER VI2 ;
  RECT 1352.400 0.200 1353.200 1.000 ;
  LAYER VI3 ;
  RECT 1352.400 0.200 1353.200 1.000 ;
  LAYER VI1 ;
  RECT 1351.200 0.200 1352.000 1.000 ;
  LAYER VI2 ;
  RECT 1351.200 0.200 1352.000 1.000 ;
  LAYER VI3 ;
  RECT 1351.200 0.200 1352.000 1.000 ;
  LAYER VI1 ;
  RECT 1345.200 0.200 1346.000 1.000 ;
  LAYER VI2 ;
  RECT 1345.200 0.200 1346.000 1.000 ;
  LAYER VI3 ;
  RECT 1345.200 0.200 1346.000 1.000 ;
  LAYER VI1 ;
  RECT 1338.000 0.200 1338.800 1.000 ;
  LAYER VI2 ;
  RECT 1338.000 0.200 1338.800 1.000 ;
  LAYER VI3 ;
  RECT 1338.000 0.200 1338.800 1.000 ;
  LAYER VI1 ;
  RECT 1335.200 0.200 1336.000 1.000 ;
  LAYER VI2 ;
  RECT 1335.200 0.200 1336.000 1.000 ;
  LAYER VI3 ;
  RECT 1335.200 0.200 1336.000 1.000 ;
  LAYER VI1 ;
  RECT 1332.400 0.200 1333.200 1.000 ;
  LAYER VI2 ;
  RECT 1332.400 0.200 1333.200 1.000 ;
  LAYER VI3 ;
  RECT 1332.400 0.200 1333.200 1.000 ;
  LAYER VI1 ;
  RECT 1330.000 0.200 1330.800 1.000 ;
  LAYER VI2 ;
  RECT 1330.000 0.200 1330.800 1.000 ;
  LAYER VI3 ;
  RECT 1330.000 0.200 1330.800 1.000 ;
  LAYER VI1 ;
  RECT 1328.400 0.200 1329.200 1.000 ;
  LAYER VI2 ;
  RECT 1328.400 0.200 1329.200 1.000 ;
  LAYER VI3 ;
  RECT 1328.400 0.200 1329.200 1.000 ;
  LAYER VI1 ;
  RECT 1326.000 0.200 1326.800 1.000 ;
  LAYER VI2 ;
  RECT 1326.000 0.200 1326.800 1.000 ;
  LAYER VI3 ;
  RECT 1326.000 0.200 1326.800 1.000 ;
  LAYER VI1 ;
  RECT 1324.400 0.200 1325.200 1.000 ;
  LAYER VI2 ;
  RECT 1324.400 0.200 1325.200 1.000 ;
  LAYER VI3 ;
  RECT 1324.400 0.200 1325.200 1.000 ;
  LAYER VI1 ;
  RECT 1322.000 0.200 1322.800 1.000 ;
  LAYER VI2 ;
  RECT 1322.000 0.200 1322.800 1.000 ;
  LAYER VI3 ;
  RECT 1322.000 0.200 1322.800 1.000 ;
  LAYER VI1 ;
  RECT 1320.400 0.200 1321.200 1.000 ;
  LAYER VI2 ;
  RECT 1320.400 0.200 1321.200 1.000 ;
  LAYER VI3 ;
  RECT 1320.400 0.200 1321.200 1.000 ;
  LAYER VI1 ;
  RECT 1311.200 0.200 1312.000 1.000 ;
  LAYER VI2 ;
  RECT 1311.200 0.200 1312.000 1.000 ;
  LAYER VI3 ;
  RECT 1311.200 0.200 1312.000 1.000 ;
  LAYER VI1 ;
  RECT 1296.400 0.200 1297.200 1.000 ;
  LAYER VI2 ;
  RECT 1296.400 0.200 1297.200 1.000 ;
  LAYER VI3 ;
  RECT 1296.400 0.200 1297.200 1.000 ;
  LAYER VI1 ;
  RECT 1291.200 0.200 1292.000 1.000 ;
  LAYER VI2 ;
  RECT 1291.200 0.200 1292.000 1.000 ;
  LAYER VI3 ;
  RECT 1291.200 0.200 1292.000 1.000 ;
  LAYER VI1 ;
  RECT 1276.800 0.200 1277.600 1.000 ;
  LAYER VI2 ;
  RECT 1276.800 0.200 1277.600 1.000 ;
  LAYER VI3 ;
  RECT 1276.800 0.200 1277.600 1.000 ;
  LAYER VI1 ;
  RECT 1270.400 0.200 1271.200 1.000 ;
  LAYER VI2 ;
  RECT 1270.400 0.200 1271.200 1.000 ;
  LAYER VI3 ;
  RECT 1270.400 0.200 1271.200 1.000 ;
  LAYER VI1 ;
  RECT 1255.600 0.200 1256.400 1.000 ;
  LAYER VI2 ;
  RECT 1255.600 0.200 1256.400 1.000 ;
  LAYER VI3 ;
  RECT 1255.600 0.200 1256.400 1.000 ;
  LAYER VI1 ;
  RECT 1250.400 0.200 1251.200 1.000 ;
  LAYER VI2 ;
  RECT 1250.400 0.200 1251.200 1.000 ;
  LAYER VI3 ;
  RECT 1250.400 0.200 1251.200 1.000 ;
  LAYER VI1 ;
  RECT 1235.600 0.200 1236.400 1.000 ;
  LAYER VI2 ;
  RECT 1235.600 0.200 1236.400 1.000 ;
  LAYER VI3 ;
  RECT 1235.600 0.200 1236.400 1.000 ;
  LAYER VI1 ;
  RECT 1229.200 0.200 1230.000 1.000 ;
  LAYER VI2 ;
  RECT 1229.200 0.200 1230.000 1.000 ;
  LAYER VI3 ;
  RECT 1229.200 0.200 1230.000 1.000 ;
  LAYER VI1 ;
  RECT 1214.800 0.200 1215.600 1.000 ;
  LAYER VI2 ;
  RECT 1214.800 0.200 1215.600 1.000 ;
  LAYER VI3 ;
  RECT 1214.800 0.200 1215.600 1.000 ;
  LAYER VI1 ;
  RECT 1209.600 0.200 1210.400 1.000 ;
  LAYER VI2 ;
  RECT 1209.600 0.200 1210.400 1.000 ;
  LAYER VI3 ;
  RECT 1209.600 0.200 1210.400 1.000 ;
  LAYER VI1 ;
  RECT 1194.800 0.200 1195.600 1.000 ;
  LAYER VI2 ;
  RECT 1194.800 0.200 1195.600 1.000 ;
  LAYER VI3 ;
  RECT 1194.800 0.200 1195.600 1.000 ;
  LAYER VI1 ;
  RECT 1188.400 0.200 1189.200 1.000 ;
  LAYER VI2 ;
  RECT 1188.400 0.200 1189.200 1.000 ;
  LAYER VI3 ;
  RECT 1188.400 0.200 1189.200 1.000 ;
  LAYER VI1 ;
  RECT 1173.600 0.200 1174.400 1.000 ;
  LAYER VI2 ;
  RECT 1173.600 0.200 1174.400 1.000 ;
  LAYER VI3 ;
  RECT 1173.600 0.200 1174.400 1.000 ;
  LAYER VI1 ;
  RECT 1168.400 0.200 1169.200 1.000 ;
  LAYER VI2 ;
  RECT 1168.400 0.200 1169.200 1.000 ;
  LAYER VI3 ;
  RECT 1168.400 0.200 1169.200 1.000 ;
  LAYER VI1 ;
  RECT 1155.600 0.200 1156.400 1.000 ;
  LAYER VI2 ;
  RECT 1155.600 0.200 1156.400 1.000 ;
  LAYER VI3 ;
  RECT 1155.600 0.200 1156.400 1.000 ;
  LAYER VI1 ;
  RECT 1154.000 0.200 1154.800 1.000 ;
  LAYER VI2 ;
  RECT 1154.000 0.200 1154.800 1.000 ;
  LAYER VI3 ;
  RECT 1154.000 0.200 1154.800 1.000 ;
  LAYER VI1 ;
  RECT 1147.600 0.200 1148.400 1.000 ;
  LAYER VI2 ;
  RECT 1147.600 0.200 1148.400 1.000 ;
  LAYER VI3 ;
  RECT 1147.600 0.200 1148.400 1.000 ;
  LAYER VI1 ;
  RECT 1132.800 0.200 1133.600 1.000 ;
  LAYER VI2 ;
  RECT 1132.800 0.200 1133.600 1.000 ;
  LAYER VI3 ;
  RECT 1132.800 0.200 1133.600 1.000 ;
  LAYER VI1 ;
  RECT 1127.600 0.200 1128.400 1.000 ;
  LAYER VI2 ;
  RECT 1127.600 0.200 1128.400 1.000 ;
  LAYER VI3 ;
  RECT 1127.600 0.200 1128.400 1.000 ;
  LAYER VI1 ;
  RECT 1113.200 0.200 1114.000 1.000 ;
  LAYER VI2 ;
  RECT 1113.200 0.200 1114.000 1.000 ;
  LAYER VI3 ;
  RECT 1113.200 0.200 1114.000 1.000 ;
  LAYER VI1 ;
  RECT 1106.400 0.200 1107.200 1.000 ;
  LAYER VI2 ;
  RECT 1106.400 0.200 1107.200 1.000 ;
  LAYER VI3 ;
  RECT 1106.400 0.200 1107.200 1.000 ;
  LAYER VI1 ;
  RECT 1092.000 0.200 1092.800 1.000 ;
  LAYER VI2 ;
  RECT 1092.000 0.200 1092.800 1.000 ;
  LAYER VI3 ;
  RECT 1092.000 0.200 1092.800 1.000 ;
  LAYER VI1 ;
  RECT 1086.800 0.200 1087.600 1.000 ;
  LAYER VI2 ;
  RECT 1086.800 0.200 1087.600 1.000 ;
  LAYER VI3 ;
  RECT 1086.800 0.200 1087.600 1.000 ;
  LAYER VI1 ;
  RECT 1072.000 0.200 1072.800 1.000 ;
  LAYER VI2 ;
  RECT 1072.000 0.200 1072.800 1.000 ;
  LAYER VI3 ;
  RECT 1072.000 0.200 1072.800 1.000 ;
  LAYER VI1 ;
  RECT 1065.600 0.200 1066.400 1.000 ;
  LAYER VI2 ;
  RECT 1065.600 0.200 1066.400 1.000 ;
  LAYER VI3 ;
  RECT 1065.600 0.200 1066.400 1.000 ;
  LAYER VI1 ;
  RECT 1051.200 0.200 1052.000 1.000 ;
  LAYER VI2 ;
  RECT 1051.200 0.200 1052.000 1.000 ;
  LAYER VI3 ;
  RECT 1051.200 0.200 1052.000 1.000 ;
  LAYER VI1 ;
  RECT 1045.600 0.200 1046.400 1.000 ;
  LAYER VI2 ;
  RECT 1045.600 0.200 1046.400 1.000 ;
  LAYER VI3 ;
  RECT 1045.600 0.200 1046.400 1.000 ;
  LAYER VI1 ;
  RECT 1031.200 0.200 1032.000 1.000 ;
  LAYER VI2 ;
  RECT 1031.200 0.200 1032.000 1.000 ;
  LAYER VI3 ;
  RECT 1031.200 0.200 1032.000 1.000 ;
  LAYER VI1 ;
  RECT 1024.800 0.200 1025.600 1.000 ;
  LAYER VI2 ;
  RECT 1024.800 0.200 1025.600 1.000 ;
  LAYER VI3 ;
  RECT 1024.800 0.200 1025.600 1.000 ;
  LAYER VI1 ;
  RECT 1010.000 0.200 1010.800 1.000 ;
  LAYER VI2 ;
  RECT 1010.000 0.200 1010.800 1.000 ;
  LAYER VI3 ;
  RECT 1010.000 0.200 1010.800 1.000 ;
  LAYER VI1 ;
  RECT 1004.800 0.200 1005.600 1.000 ;
  LAYER VI2 ;
  RECT 1004.800 0.200 1005.600 1.000 ;
  LAYER VI3 ;
  RECT 1004.800 0.200 1005.600 1.000 ;
  LAYER VI1 ;
  RECT 992.000 0.200 992.800 1.000 ;
  LAYER VI2 ;
  RECT 992.000 0.200 992.800 1.000 ;
  LAYER VI3 ;
  RECT 992.000 0.200 992.800 1.000 ;
  LAYER VI1 ;
  RECT 990.400 0.200 991.200 1.000 ;
  LAYER VI2 ;
  RECT 990.400 0.200 991.200 1.000 ;
  LAYER VI3 ;
  RECT 990.400 0.200 991.200 1.000 ;
  LAYER VI1 ;
  RECT 983.600 0.200 984.400 1.000 ;
  LAYER VI2 ;
  RECT 983.600 0.200 984.400 1.000 ;
  LAYER VI3 ;
  RECT 983.600 0.200 984.400 1.000 ;
  LAYER VI1 ;
  RECT 969.200 0.200 970.000 1.000 ;
  LAYER VI2 ;
  RECT 969.200 0.200 970.000 1.000 ;
  LAYER VI3 ;
  RECT 969.200 0.200 970.000 1.000 ;
  LAYER VI1 ;
  RECT 964.000 0.200 964.800 1.000 ;
  LAYER VI2 ;
  RECT 964.000 0.200 964.800 1.000 ;
  LAYER VI3 ;
  RECT 964.000 0.200 964.800 1.000 ;
  LAYER VI1 ;
  RECT 949.200 0.200 950.000 1.000 ;
  LAYER VI2 ;
  RECT 949.200 0.200 950.000 1.000 ;
  LAYER VI3 ;
  RECT 949.200 0.200 950.000 1.000 ;
  LAYER VI1 ;
  RECT 942.800 0.200 943.600 1.000 ;
  LAYER VI2 ;
  RECT 942.800 0.200 943.600 1.000 ;
  LAYER VI3 ;
  RECT 942.800 0.200 943.600 1.000 ;
  LAYER VI1 ;
  RECT 928.400 0.200 929.200 1.000 ;
  LAYER VI2 ;
  RECT 928.400 0.200 929.200 1.000 ;
  LAYER VI3 ;
  RECT 928.400 0.200 929.200 1.000 ;
  LAYER VI1 ;
  RECT 923.200 0.200 924.000 1.000 ;
  LAYER VI2 ;
  RECT 923.200 0.200 924.000 1.000 ;
  LAYER VI3 ;
  RECT 923.200 0.200 924.000 1.000 ;
  LAYER VI1 ;
  RECT 908.400 0.200 909.200 1.000 ;
  LAYER VI2 ;
  RECT 908.400 0.200 909.200 1.000 ;
  LAYER VI3 ;
  RECT 908.400 0.200 909.200 1.000 ;
  LAYER VI1 ;
  RECT 902.000 0.200 902.800 1.000 ;
  LAYER VI2 ;
  RECT 902.000 0.200 902.800 1.000 ;
  LAYER VI3 ;
  RECT 902.000 0.200 902.800 1.000 ;
  LAYER VI1 ;
  RECT 887.200 0.200 888.000 1.000 ;
  LAYER VI2 ;
  RECT 887.200 0.200 888.000 1.000 ;
  LAYER VI3 ;
  RECT 887.200 0.200 888.000 1.000 ;
  LAYER VI1 ;
  RECT 882.000 0.200 882.800 1.000 ;
  LAYER VI2 ;
  RECT 882.000 0.200 882.800 1.000 ;
  LAYER VI3 ;
  RECT 882.000 0.200 882.800 1.000 ;
  LAYER VI1 ;
  RECT 867.600 0.200 868.400 1.000 ;
  LAYER VI2 ;
  RECT 867.600 0.200 868.400 1.000 ;
  LAYER VI3 ;
  RECT 867.600 0.200 868.400 1.000 ;
  LAYER VI1 ;
  RECT 861.200 0.200 862.000 1.000 ;
  LAYER VI2 ;
  RECT 861.200 0.200 862.000 1.000 ;
  LAYER VI3 ;
  RECT 861.200 0.200 862.000 1.000 ;
  LAYER VI1 ;
  RECT 846.400 0.200 847.200 1.000 ;
  LAYER VI2 ;
  RECT 846.400 0.200 847.200 1.000 ;
  LAYER VI3 ;
  RECT 846.400 0.200 847.200 1.000 ;
  LAYER VI1 ;
  RECT 841.200 0.200 842.000 1.000 ;
  LAYER VI2 ;
  RECT 841.200 0.200 842.000 1.000 ;
  LAYER VI3 ;
  RECT 841.200 0.200 842.000 1.000 ;
  LAYER VI1 ;
  RECT 828.400 0.200 829.200 1.000 ;
  LAYER VI2 ;
  RECT 828.400 0.200 829.200 1.000 ;
  LAYER VI3 ;
  RECT 828.400 0.200 829.200 1.000 ;
  LAYER VI1 ;
  RECT 826.400 0.200 827.200 1.000 ;
  LAYER VI2 ;
  RECT 826.400 0.200 827.200 1.000 ;
  LAYER VI3 ;
  RECT 826.400 0.200 827.200 1.000 ;
  LAYER VI1 ;
  RECT 820.000 0.200 820.800 1.000 ;
  LAYER VI2 ;
  RECT 820.000 0.200 820.800 1.000 ;
  LAYER VI3 ;
  RECT 820.000 0.200 820.800 1.000 ;
  LAYER VI1 ;
  RECT 805.600 0.200 806.400 1.000 ;
  LAYER VI2 ;
  RECT 805.600 0.200 806.400 1.000 ;
  LAYER VI3 ;
  RECT 805.600 0.200 806.400 1.000 ;
  LAYER VI1 ;
  RECT 800.400 0.200 801.200 1.000 ;
  LAYER VI2 ;
  RECT 800.400 0.200 801.200 1.000 ;
  LAYER VI3 ;
  RECT 800.400 0.200 801.200 1.000 ;
  LAYER VI1 ;
  RECT 785.600 0.200 786.400 1.000 ;
  LAYER VI2 ;
  RECT 785.600 0.200 786.400 1.000 ;
  LAYER VI3 ;
  RECT 785.600 0.200 786.400 1.000 ;
  LAYER VI1 ;
  RECT 779.200 0.200 780.000 1.000 ;
  LAYER VI2 ;
  RECT 779.200 0.200 780.000 1.000 ;
  LAYER VI3 ;
  RECT 779.200 0.200 780.000 1.000 ;
  LAYER VI1 ;
  RECT 764.400 0.200 765.200 1.000 ;
  LAYER VI2 ;
  RECT 764.400 0.200 765.200 1.000 ;
  LAYER VI3 ;
  RECT 764.400 0.200 765.200 1.000 ;
  LAYER VI1 ;
  RECT 759.200 0.200 760.000 1.000 ;
  LAYER VI2 ;
  RECT 759.200 0.200 760.000 1.000 ;
  LAYER VI3 ;
  RECT 759.200 0.200 760.000 1.000 ;
  LAYER VI1 ;
  RECT 744.800 0.200 745.600 1.000 ;
  LAYER VI2 ;
  RECT 744.800 0.200 745.600 1.000 ;
  LAYER VI3 ;
  RECT 744.800 0.200 745.600 1.000 ;
  LAYER VI1 ;
  RECT 738.400 0.200 739.200 1.000 ;
  LAYER VI2 ;
  RECT 738.400 0.200 739.200 1.000 ;
  LAYER VI3 ;
  RECT 738.400 0.200 739.200 1.000 ;
  LAYER VI1 ;
  RECT 723.600 0.200 724.400 1.000 ;
  LAYER VI2 ;
  RECT 723.600 0.200 724.400 1.000 ;
  LAYER VI3 ;
  RECT 723.600 0.200 724.400 1.000 ;
  LAYER VI1 ;
  RECT 718.400 0.200 719.200 1.000 ;
  LAYER VI2 ;
  RECT 718.400 0.200 719.200 1.000 ;
  LAYER VI3 ;
  RECT 718.400 0.200 719.200 1.000 ;
  LAYER VI1 ;
  RECT 704.000 0.200 704.800 1.000 ;
  LAYER VI2 ;
  RECT 704.000 0.200 704.800 1.000 ;
  LAYER VI3 ;
  RECT 704.000 0.200 704.800 1.000 ;
  LAYER VI1 ;
  RECT 697.200 0.200 698.000 1.000 ;
  LAYER VI2 ;
  RECT 697.200 0.200 698.000 1.000 ;
  LAYER VI3 ;
  RECT 697.200 0.200 698.000 1.000 ;
  LAYER VI1 ;
  RECT 682.800 0.200 683.600 1.000 ;
  LAYER VI2 ;
  RECT 682.800 0.200 683.600 1.000 ;
  LAYER VI3 ;
  RECT 682.800 0.200 683.600 1.000 ;
  LAYER VI1 ;
  RECT 677.600 0.200 678.400 1.000 ;
  LAYER VI2 ;
  RECT 677.600 0.200 678.400 1.000 ;
  LAYER VI3 ;
  RECT 677.600 0.200 678.400 1.000 ;
  LAYER VI1 ;
  RECT 664.800 0.200 665.600 1.000 ;
  LAYER VI2 ;
  RECT 664.800 0.200 665.600 1.000 ;
  LAYER VI3 ;
  RECT 664.800 0.200 665.600 1.000 ;
  LAYER VI1 ;
  RECT 662.800 0.200 663.600 1.000 ;
  LAYER VI2 ;
  RECT 662.800 0.200 663.600 1.000 ;
  LAYER VI3 ;
  RECT 662.800 0.200 663.600 1.000 ;
  LAYER VI1 ;
  RECT 656.400 0.200 657.200 1.000 ;
  LAYER VI2 ;
  RECT 656.400 0.200 657.200 1.000 ;
  LAYER VI3 ;
  RECT 656.400 0.200 657.200 1.000 ;
  LAYER VI1 ;
  RECT 642.000 0.200 642.800 1.000 ;
  LAYER VI2 ;
  RECT 642.000 0.200 642.800 1.000 ;
  LAYER VI3 ;
  RECT 642.000 0.200 642.800 1.000 ;
  LAYER VI1 ;
  RECT 636.400 0.200 637.200 1.000 ;
  LAYER VI2 ;
  RECT 636.400 0.200 637.200 1.000 ;
  LAYER VI3 ;
  RECT 636.400 0.200 637.200 1.000 ;
  LAYER VI1 ;
  RECT 622.000 0.200 622.800 1.000 ;
  LAYER VI2 ;
  RECT 622.000 0.200 622.800 1.000 ;
  LAYER VI3 ;
  RECT 622.000 0.200 622.800 1.000 ;
  LAYER VI1 ;
  RECT 615.600 0.200 616.400 1.000 ;
  LAYER VI2 ;
  RECT 615.600 0.200 616.400 1.000 ;
  LAYER VI3 ;
  RECT 615.600 0.200 616.400 1.000 ;
  LAYER VI1 ;
  RECT 600.800 0.200 601.600 1.000 ;
  LAYER VI2 ;
  RECT 600.800 0.200 601.600 1.000 ;
  LAYER VI3 ;
  RECT 600.800 0.200 601.600 1.000 ;
  LAYER VI1 ;
  RECT 595.600 0.200 596.400 1.000 ;
  LAYER VI2 ;
  RECT 595.600 0.200 596.400 1.000 ;
  LAYER VI3 ;
  RECT 595.600 0.200 596.400 1.000 ;
  LAYER VI1 ;
  RECT 581.200 0.200 582.000 1.000 ;
  LAYER VI2 ;
  RECT 581.200 0.200 582.000 1.000 ;
  LAYER VI3 ;
  RECT 581.200 0.200 582.000 1.000 ;
  LAYER VI1 ;
  RECT 574.400 0.200 575.200 1.000 ;
  LAYER VI2 ;
  RECT 574.400 0.200 575.200 1.000 ;
  LAYER VI3 ;
  RECT 574.400 0.200 575.200 1.000 ;
  LAYER VI1 ;
  RECT 560.000 0.200 560.800 1.000 ;
  LAYER VI2 ;
  RECT 560.000 0.200 560.800 1.000 ;
  LAYER VI3 ;
  RECT 560.000 0.200 560.800 1.000 ;
  LAYER VI1 ;
  RECT 554.800 0.200 555.600 1.000 ;
  LAYER VI2 ;
  RECT 554.800 0.200 555.600 1.000 ;
  LAYER VI3 ;
  RECT 554.800 0.200 555.600 1.000 ;
  LAYER VI1 ;
  RECT 540.000 0.200 540.800 1.000 ;
  LAYER VI2 ;
  RECT 540.000 0.200 540.800 1.000 ;
  LAYER VI3 ;
  RECT 540.000 0.200 540.800 1.000 ;
  LAYER VI1 ;
  RECT 533.600 0.200 534.400 1.000 ;
  LAYER VI2 ;
  RECT 533.600 0.200 534.400 1.000 ;
  LAYER VI3 ;
  RECT 533.600 0.200 534.400 1.000 ;
  LAYER VI1 ;
  RECT 519.200 0.200 520.000 1.000 ;
  LAYER VI2 ;
  RECT 519.200 0.200 520.000 1.000 ;
  LAYER VI3 ;
  RECT 519.200 0.200 520.000 1.000 ;
  LAYER VI1 ;
  RECT 514.000 0.200 514.800 1.000 ;
  LAYER VI2 ;
  RECT 514.000 0.200 514.800 1.000 ;
  LAYER VI3 ;
  RECT 514.000 0.200 514.800 1.000 ;
  LAYER VI1 ;
  RECT 500.800 0.200 501.600 1.000 ;
  LAYER VI2 ;
  RECT 500.800 0.200 501.600 1.000 ;
  LAYER VI3 ;
  RECT 500.800 0.200 501.600 1.000 ;
  LAYER VI1 ;
  RECT 499.200 0.200 500.000 1.000 ;
  LAYER VI2 ;
  RECT 499.200 0.200 500.000 1.000 ;
  LAYER VI3 ;
  RECT 499.200 0.200 500.000 1.000 ;
  LAYER VI1 ;
  RECT 492.800 0.200 493.600 1.000 ;
  LAYER VI2 ;
  RECT 492.800 0.200 493.600 1.000 ;
  LAYER VI3 ;
  RECT 492.800 0.200 493.600 1.000 ;
  LAYER VI1 ;
  RECT 478.000 0.200 478.800 1.000 ;
  LAYER VI2 ;
  RECT 478.000 0.200 478.800 1.000 ;
  LAYER VI3 ;
  RECT 478.000 0.200 478.800 1.000 ;
  LAYER VI1 ;
  RECT 472.800 0.200 473.600 1.000 ;
  LAYER VI2 ;
  RECT 472.800 0.200 473.600 1.000 ;
  LAYER VI3 ;
  RECT 472.800 0.200 473.600 1.000 ;
  LAYER VI1 ;
  RECT 458.400 0.200 459.200 1.000 ;
  LAYER VI2 ;
  RECT 458.400 0.200 459.200 1.000 ;
  LAYER VI3 ;
  RECT 458.400 0.200 459.200 1.000 ;
  LAYER VI1 ;
  RECT 452.000 0.200 452.800 1.000 ;
  LAYER VI2 ;
  RECT 452.000 0.200 452.800 1.000 ;
  LAYER VI3 ;
  RECT 452.000 0.200 452.800 1.000 ;
  LAYER VI1 ;
  RECT 437.200 0.200 438.000 1.000 ;
  LAYER VI2 ;
  RECT 437.200 0.200 438.000 1.000 ;
  LAYER VI3 ;
  RECT 437.200 0.200 438.000 1.000 ;
  LAYER VI1 ;
  RECT 432.000 0.200 432.800 1.000 ;
  LAYER VI2 ;
  RECT 432.000 0.200 432.800 1.000 ;
  LAYER VI3 ;
  RECT 432.000 0.200 432.800 1.000 ;
  LAYER VI1 ;
  RECT 417.200 0.200 418.000 1.000 ;
  LAYER VI2 ;
  RECT 417.200 0.200 418.000 1.000 ;
  LAYER VI3 ;
  RECT 417.200 0.200 418.000 1.000 ;
  LAYER VI1 ;
  RECT 410.800 0.200 411.600 1.000 ;
  LAYER VI2 ;
  RECT 410.800 0.200 411.600 1.000 ;
  LAYER VI3 ;
  RECT 410.800 0.200 411.600 1.000 ;
  LAYER VI1 ;
  RECT 396.400 0.200 397.200 1.000 ;
  LAYER VI2 ;
  RECT 396.400 0.200 397.200 1.000 ;
  LAYER VI3 ;
  RECT 396.400 0.200 397.200 1.000 ;
  LAYER VI1 ;
  RECT 391.200 0.200 392.000 1.000 ;
  LAYER VI2 ;
  RECT 391.200 0.200 392.000 1.000 ;
  LAYER VI3 ;
  RECT 391.200 0.200 392.000 1.000 ;
  LAYER VI1 ;
  RECT 376.400 0.200 377.200 1.000 ;
  LAYER VI2 ;
  RECT 376.400 0.200 377.200 1.000 ;
  LAYER VI3 ;
  RECT 376.400 0.200 377.200 1.000 ;
  LAYER VI1 ;
  RECT 370.000 0.200 370.800 1.000 ;
  LAYER VI2 ;
  RECT 370.000 0.200 370.800 1.000 ;
  LAYER VI3 ;
  RECT 370.000 0.200 370.800 1.000 ;
  LAYER VI1 ;
  RECT 355.200 0.200 356.000 1.000 ;
  LAYER VI2 ;
  RECT 355.200 0.200 356.000 1.000 ;
  LAYER VI3 ;
  RECT 355.200 0.200 356.000 1.000 ;
  LAYER VI1 ;
  RECT 350.000 0.200 350.800 1.000 ;
  LAYER VI2 ;
  RECT 350.000 0.200 350.800 1.000 ;
  LAYER VI3 ;
  RECT 350.000 0.200 350.800 1.000 ;
  LAYER VI1 ;
  RECT 337.200 0.200 338.000 1.000 ;
  LAYER VI2 ;
  RECT 337.200 0.200 338.000 1.000 ;
  LAYER VI3 ;
  RECT 337.200 0.200 338.000 1.000 ;
  LAYER VI1 ;
  RECT 335.600 0.200 336.400 1.000 ;
  LAYER VI2 ;
  RECT 335.600 0.200 336.400 1.000 ;
  LAYER VI3 ;
  RECT 335.600 0.200 336.400 1.000 ;
  LAYER VI1 ;
  RECT 329.200 0.200 330.000 1.000 ;
  LAYER VI2 ;
  RECT 329.200 0.200 330.000 1.000 ;
  LAYER VI3 ;
  RECT 329.200 0.200 330.000 1.000 ;
  LAYER VI1 ;
  RECT 314.400 0.200 315.200 1.000 ;
  LAYER VI2 ;
  RECT 314.400 0.200 315.200 1.000 ;
  LAYER VI3 ;
  RECT 314.400 0.200 315.200 1.000 ;
  LAYER VI1 ;
  RECT 309.200 0.200 310.000 1.000 ;
  LAYER VI2 ;
  RECT 309.200 0.200 310.000 1.000 ;
  LAYER VI3 ;
  RECT 309.200 0.200 310.000 1.000 ;
  LAYER VI1 ;
  RECT 294.800 0.200 295.600 1.000 ;
  LAYER VI2 ;
  RECT 294.800 0.200 295.600 1.000 ;
  LAYER VI3 ;
  RECT 294.800 0.200 295.600 1.000 ;
  LAYER VI1 ;
  RECT 288.000 0.200 288.800 1.000 ;
  LAYER VI2 ;
  RECT 288.000 0.200 288.800 1.000 ;
  LAYER VI3 ;
  RECT 288.000 0.200 288.800 1.000 ;
  LAYER VI1 ;
  RECT 273.600 0.200 274.400 1.000 ;
  LAYER VI2 ;
  RECT 273.600 0.200 274.400 1.000 ;
  LAYER VI3 ;
  RECT 273.600 0.200 274.400 1.000 ;
  LAYER VI1 ;
  RECT 268.400 0.200 269.200 1.000 ;
  LAYER VI2 ;
  RECT 268.400 0.200 269.200 1.000 ;
  LAYER VI3 ;
  RECT 268.400 0.200 269.200 1.000 ;
  LAYER VI1 ;
  RECT 253.600 0.200 254.400 1.000 ;
  LAYER VI2 ;
  RECT 253.600 0.200 254.400 1.000 ;
  LAYER VI3 ;
  RECT 253.600 0.200 254.400 1.000 ;
  LAYER VI1 ;
  RECT 247.200 0.200 248.000 1.000 ;
  LAYER VI2 ;
  RECT 247.200 0.200 248.000 1.000 ;
  LAYER VI3 ;
  RECT 247.200 0.200 248.000 1.000 ;
  LAYER VI1 ;
  RECT 232.800 0.200 233.600 1.000 ;
  LAYER VI2 ;
  RECT 232.800 0.200 233.600 1.000 ;
  LAYER VI3 ;
  RECT 232.800 0.200 233.600 1.000 ;
  LAYER VI1 ;
  RECT 227.200 0.200 228.000 1.000 ;
  LAYER VI2 ;
  RECT 227.200 0.200 228.000 1.000 ;
  LAYER VI3 ;
  RECT 227.200 0.200 228.000 1.000 ;
  LAYER VI1 ;
  RECT 212.800 0.200 213.600 1.000 ;
  LAYER VI2 ;
  RECT 212.800 0.200 213.600 1.000 ;
  LAYER VI3 ;
  RECT 212.800 0.200 213.600 1.000 ;
  LAYER VI1 ;
  RECT 206.400 0.200 207.200 1.000 ;
  LAYER VI2 ;
  RECT 206.400 0.200 207.200 1.000 ;
  LAYER VI3 ;
  RECT 206.400 0.200 207.200 1.000 ;
  LAYER VI1 ;
  RECT 191.600 0.200 192.400 1.000 ;
  LAYER VI2 ;
  RECT 191.600 0.200 192.400 1.000 ;
  LAYER VI3 ;
  RECT 191.600 0.200 192.400 1.000 ;
  LAYER VI1 ;
  RECT 186.400 0.200 187.200 1.000 ;
  LAYER VI2 ;
  RECT 186.400 0.200 187.200 1.000 ;
  LAYER VI3 ;
  RECT 186.400 0.200 187.200 1.000 ;
  LAYER VI1 ;
  RECT 173.600 0.200 174.400 1.000 ;
  LAYER VI2 ;
  RECT 173.600 0.200 174.400 1.000 ;
  LAYER VI3 ;
  RECT 173.600 0.200 174.400 1.000 ;
  LAYER VI1 ;
  RECT 172.000 0.200 172.800 1.000 ;
  LAYER VI2 ;
  RECT 172.000 0.200 172.800 1.000 ;
  LAYER VI3 ;
  RECT 172.000 0.200 172.800 1.000 ;
  LAYER VI1 ;
  RECT 165.200 0.200 166.000 1.000 ;
  LAYER VI2 ;
  RECT 165.200 0.200 166.000 1.000 ;
  LAYER VI3 ;
  RECT 165.200 0.200 166.000 1.000 ;
  LAYER VI1 ;
  RECT 150.800 0.200 151.600 1.000 ;
  LAYER VI2 ;
  RECT 150.800 0.200 151.600 1.000 ;
  LAYER VI3 ;
  RECT 150.800 0.200 151.600 1.000 ;
  LAYER VI1 ;
  RECT 145.600 0.200 146.400 1.000 ;
  LAYER VI2 ;
  RECT 145.600 0.200 146.400 1.000 ;
  LAYER VI3 ;
  RECT 145.600 0.200 146.400 1.000 ;
  LAYER VI1 ;
  RECT 130.800 0.200 131.600 1.000 ;
  LAYER VI2 ;
  RECT 130.800 0.200 131.600 1.000 ;
  LAYER VI3 ;
  RECT 130.800 0.200 131.600 1.000 ;
  LAYER VI1 ;
  RECT 124.400 0.200 125.200 1.000 ;
  LAYER VI2 ;
  RECT 124.400 0.200 125.200 1.000 ;
  LAYER VI3 ;
  RECT 124.400 0.200 125.200 1.000 ;
  LAYER VI1 ;
  RECT 110.000 0.200 110.800 1.000 ;
  LAYER VI2 ;
  RECT 110.000 0.200 110.800 1.000 ;
  LAYER VI3 ;
  RECT 110.000 0.200 110.800 1.000 ;
  LAYER VI1 ;
  RECT 104.800 0.200 105.600 1.000 ;
  LAYER VI2 ;
  RECT 104.800 0.200 105.600 1.000 ;
  LAYER VI3 ;
  RECT 104.800 0.200 105.600 1.000 ;
  LAYER VI1 ;
  RECT 90.000 0.200 90.800 1.000 ;
  LAYER VI2 ;
  RECT 90.000 0.200 90.800 1.000 ;
  LAYER VI3 ;
  RECT 90.000 0.200 90.800 1.000 ;
  LAYER VI1 ;
  RECT 83.600 0.200 84.400 1.000 ;
  LAYER VI2 ;
  RECT 83.600 0.200 84.400 1.000 ;
  LAYER VI3 ;
  RECT 83.600 0.200 84.400 1.000 ;
  LAYER VI1 ;
  RECT 68.800 0.200 69.600 1.000 ;
  LAYER VI2 ;
  RECT 68.800 0.200 69.600 1.000 ;
  LAYER VI3 ;
  RECT 68.800 0.200 69.600 1.000 ;
  LAYER VI1 ;
  RECT 63.600 0.200 64.400 1.000 ;
  LAYER VI2 ;
  RECT 63.600 0.200 64.400 1.000 ;
  LAYER VI3 ;
  RECT 63.600 0.200 64.400 1.000 ;
  LAYER VI1 ;
  RECT 49.200 0.200 50.000 1.000 ;
  LAYER VI2 ;
  RECT 49.200 0.200 50.000 1.000 ;
  LAYER VI3 ;
  RECT 49.200 0.200 50.000 1.000 ;
  LAYER VI1 ;
  RECT 42.800 0.200 43.600 1.000 ;
  LAYER VI2 ;
  RECT 42.800 0.200 43.600 1.000 ;
  LAYER VI3 ;
  RECT 42.800 0.200 43.600 1.000 ;
  LAYER VI1 ;
  RECT 28.000 0.200 28.800 1.000 ;
  LAYER VI2 ;
  RECT 28.000 0.200 28.800 1.000 ;
  LAYER VI3 ;
  RECT 28.000 0.200 28.800 1.000 ;
  LAYER VI1 ;
  RECT 22.800 0.200 23.600 1.000 ;
  LAYER VI2 ;
  RECT 22.800 0.200 23.600 1.000 ;
  LAYER VI3 ;
  RECT 22.800 0.200 23.600 1.000 ;
  LAYER VI1 ;
  RECT 10.000 0.200 10.800 1.000 ;
  LAYER VI2 ;
  RECT 10.000 0.200 10.800 1.000 ;
  LAYER VI3 ;
  RECT 10.000 0.200 10.800 1.000 ;
  LAYER VI1 ;
  RECT 8.000 0.200 8.800 1.000 ;
  LAYER VI2 ;
  RECT 8.000 0.200 8.800 1.000 ;
  LAYER VI3 ;
  RECT 8.000 0.200 8.800 1.000 ;
  LAYER VI3 ;
  RECT 2687.800 9.570 2688.660 11.170 ;
  LAYER VI3 ;
  RECT 2688.260 10.770 2688.460 10.970 ;
  LAYER VI3 ;
  RECT 2688.260 10.370 2688.460 10.570 ;
  LAYER VI3 ;
  RECT 2688.260 9.970 2688.460 10.170 ;
  LAYER VI3 ;
  RECT 2688.260 9.570 2688.460 9.770 ;
  LAYER VI3 ;
  RECT 2687.860 10.770 2688.060 10.970 ;
  LAYER VI3 ;
  RECT 2687.860 10.370 2688.060 10.570 ;
  LAYER VI3 ;
  RECT 2687.860 9.970 2688.060 10.170 ;
  LAYER VI3 ;
  RECT 2687.860 9.570 2688.060 9.770 ;
  LAYER VI2 ;
  RECT 2687.800 9.570 2688.660 11.170 ;
  LAYER VI2 ;
  RECT 2688.260 10.770 2688.460 10.970 ;
  LAYER VI2 ;
  RECT 2688.260 10.370 2688.460 10.570 ;
  LAYER VI2 ;
  RECT 2688.260 9.970 2688.460 10.170 ;
  LAYER VI2 ;
  RECT 2688.260 9.570 2688.460 9.770 ;
  LAYER VI2 ;
  RECT 2687.860 10.770 2688.060 10.970 ;
  LAYER VI2 ;
  RECT 2687.860 10.370 2688.060 10.570 ;
  LAYER VI2 ;
  RECT 2687.860 9.970 2688.060 10.170 ;
  LAYER VI2 ;
  RECT 2687.860 9.570 2688.060 9.770 ;
  LAYER VI3 ;
  RECT 2687.800 14.200 2688.660 15.200 ;
  LAYER VI3 ;
  RECT 2688.260 14.600 2688.460 14.800 ;
  LAYER VI3 ;
  RECT 2688.260 14.200 2688.460 14.400 ;
  LAYER VI3 ;
  RECT 2687.860 14.600 2688.060 14.800 ;
  LAYER VI3 ;
  RECT 2687.860 14.200 2688.060 14.400 ;
  LAYER VI2 ;
  RECT 2687.800 14.200 2688.660 15.200 ;
  LAYER VI2 ;
  RECT 2688.260 14.600 2688.460 14.800 ;
  LAYER VI2 ;
  RECT 2688.260 14.200 2688.460 14.400 ;
  LAYER VI2 ;
  RECT 2687.860 14.600 2688.060 14.800 ;
  LAYER VI2 ;
  RECT 2687.860 14.200 2688.060 14.400 ;
  LAYER VI3 ;
  RECT 2687.800 18.730 2688.660 19.730 ;
  LAYER VI3 ;
  RECT 2688.260 19.130 2688.460 19.330 ;
  LAYER VI3 ;
  RECT 2688.260 18.730 2688.460 18.930 ;
  LAYER VI3 ;
  RECT 2687.860 19.130 2688.060 19.330 ;
  LAYER VI3 ;
  RECT 2687.860 18.730 2688.060 18.930 ;
  LAYER VI2 ;
  RECT 2687.800 18.730 2688.660 19.730 ;
  LAYER VI2 ;
  RECT 2688.260 19.130 2688.460 19.330 ;
  LAYER VI2 ;
  RECT 2688.260 18.730 2688.460 18.930 ;
  LAYER VI2 ;
  RECT 2687.860 19.130 2688.060 19.330 ;
  LAYER VI2 ;
  RECT 2687.860 18.730 2688.060 18.930 ;
  LAYER VI3 ;
  RECT 2687.800 21.230 2688.660 22.070 ;
  LAYER VI3 ;
  RECT 2688.200 21.690 2688.400 21.890 ;
  LAYER VI3 ;
  RECT 2688.200 21.290 2688.400 21.490 ;
  LAYER VI3 ;
  RECT 2687.800 21.690 2688.000 21.890 ;
  LAYER VI3 ;
  RECT 2687.800 21.290 2688.000 21.490 ;
  LAYER VI2 ;
  RECT 2687.800 21.230 2688.660 22.070 ;
  LAYER VI2 ;
  RECT 2688.200 21.690 2688.400 21.890 ;
  LAYER VI2 ;
  RECT 2688.200 21.290 2688.400 21.490 ;
  LAYER VI2 ;
  RECT 2687.800 21.690 2688.000 21.890 ;
  LAYER VI2 ;
  RECT 2687.800 21.290 2688.000 21.490 ;
  LAYER VI3 ;
  RECT 2687.800 24.170 2688.660 25.170 ;
  LAYER VI3 ;
  RECT 2688.260 24.570 2688.460 24.770 ;
  LAYER VI3 ;
  RECT 2688.260 24.170 2688.460 24.370 ;
  LAYER VI3 ;
  RECT 2687.860 24.570 2688.060 24.770 ;
  LAYER VI3 ;
  RECT 2687.860 24.170 2688.060 24.370 ;
  LAYER VI2 ;
  RECT 2687.800 24.170 2688.660 25.170 ;
  LAYER VI2 ;
  RECT 2688.260 24.570 2688.460 24.770 ;
  LAYER VI2 ;
  RECT 2688.260 24.170 2688.460 24.370 ;
  LAYER VI2 ;
  RECT 2687.860 24.570 2688.060 24.770 ;
  LAYER VI2 ;
  RECT 2687.860 24.170 2688.060 24.370 ;
  LAYER VI3 ;
  RECT 2687.800 36.320 2688.660 37.320 ;
  LAYER VI3 ;
  RECT 2688.260 36.720 2688.460 36.920 ;
  LAYER VI3 ;
  RECT 2688.260 36.320 2688.460 36.520 ;
  LAYER VI3 ;
  RECT 2687.860 36.720 2688.060 36.920 ;
  LAYER VI3 ;
  RECT 2687.860 36.320 2688.060 36.520 ;
  LAYER VI2 ;
  RECT 2687.800 36.320 2688.660 37.320 ;
  LAYER VI2 ;
  RECT 2688.260 36.720 2688.460 36.920 ;
  LAYER VI2 ;
  RECT 2688.260 36.320 2688.460 36.520 ;
  LAYER VI2 ;
  RECT 2687.860 36.720 2688.060 36.920 ;
  LAYER VI2 ;
  RECT 2687.860 36.320 2688.060 36.520 ;
  LAYER VI3 ;
  RECT 2687.800 39.480 2688.660 40.080 ;
  LAYER VI3 ;
  RECT 2688.200 39.540 2688.400 39.740 ;
  LAYER VI3 ;
  RECT 2687.800 39.540 2688.000 39.740 ;
  LAYER VI2 ;
  RECT 2687.800 39.480 2688.660 40.080 ;
  LAYER VI2 ;
  RECT 2688.200 39.540 2688.400 39.740 ;
  LAYER VI2 ;
  RECT 2687.800 39.540 2688.000 39.740 ;
  LAYER VI3 ;
  RECT 2687.800 45.560 2688.660 46.160 ;
  LAYER VI3 ;
  RECT 2688.200 45.620 2688.400 45.820 ;
  LAYER VI3 ;
  RECT 2687.800 45.620 2688.000 45.820 ;
  LAYER VI2 ;
  RECT 2687.800 45.560 2688.660 46.160 ;
  LAYER VI2 ;
  RECT 2688.200 45.620 2688.400 45.820 ;
  LAYER VI2 ;
  RECT 2687.800 45.620 2688.000 45.820 ;
  LAYER VI3 ;
  RECT 2687.800 57.100 2688.660 61.420 ;
  LAYER VI3 ;
  RECT 2688.260 61.100 2688.460 61.300 ;
  LAYER VI3 ;
  RECT 2688.260 60.700 2688.460 60.900 ;
  LAYER VI3 ;
  RECT 2688.260 60.300 2688.460 60.500 ;
  LAYER VI3 ;
  RECT 2688.260 59.900 2688.460 60.100 ;
  LAYER VI3 ;
  RECT 2688.260 59.500 2688.460 59.700 ;
  LAYER VI3 ;
  RECT 2688.260 59.100 2688.460 59.300 ;
  LAYER VI3 ;
  RECT 2688.260 58.700 2688.460 58.900 ;
  LAYER VI3 ;
  RECT 2688.260 58.300 2688.460 58.500 ;
  LAYER VI3 ;
  RECT 2688.260 57.900 2688.460 58.100 ;
  LAYER VI3 ;
  RECT 2688.260 57.500 2688.460 57.700 ;
  LAYER VI3 ;
  RECT 2688.260 57.100 2688.460 57.300 ;
  LAYER VI3 ;
  RECT 2687.860 61.100 2688.060 61.300 ;
  LAYER VI3 ;
  RECT 2687.860 60.700 2688.060 60.900 ;
  LAYER VI3 ;
  RECT 2687.860 60.300 2688.060 60.500 ;
  LAYER VI3 ;
  RECT 2687.860 59.900 2688.060 60.100 ;
  LAYER VI3 ;
  RECT 2687.860 59.500 2688.060 59.700 ;
  LAYER VI3 ;
  RECT 2687.860 59.100 2688.060 59.300 ;
  LAYER VI3 ;
  RECT 2687.860 58.700 2688.060 58.900 ;
  LAYER VI3 ;
  RECT 2687.860 58.300 2688.060 58.500 ;
  LAYER VI3 ;
  RECT 2687.860 57.900 2688.060 58.100 ;
  LAYER VI3 ;
  RECT 2687.860 57.500 2688.060 57.700 ;
  LAYER VI3 ;
  RECT 2687.860 57.100 2688.060 57.300 ;
  LAYER VI2 ;
  RECT 2687.800 57.100 2688.660 61.420 ;
  LAYER VI2 ;
  RECT 2688.260 61.100 2688.460 61.300 ;
  LAYER VI2 ;
  RECT 2688.260 60.700 2688.460 60.900 ;
  LAYER VI2 ;
  RECT 2688.260 60.300 2688.460 60.500 ;
  LAYER VI2 ;
  RECT 2688.260 59.900 2688.460 60.100 ;
  LAYER VI2 ;
  RECT 2688.260 59.500 2688.460 59.700 ;
  LAYER VI2 ;
  RECT 2688.260 59.100 2688.460 59.300 ;
  LAYER VI2 ;
  RECT 2688.260 58.700 2688.460 58.900 ;
  LAYER VI2 ;
  RECT 2688.260 58.300 2688.460 58.500 ;
  LAYER VI2 ;
  RECT 2688.260 57.900 2688.460 58.100 ;
  LAYER VI2 ;
  RECT 2688.260 57.500 2688.460 57.700 ;
  LAYER VI2 ;
  RECT 2688.260 57.100 2688.460 57.300 ;
  LAYER VI2 ;
  RECT 2687.860 61.100 2688.060 61.300 ;
  LAYER VI2 ;
  RECT 2687.860 60.700 2688.060 60.900 ;
  LAYER VI2 ;
  RECT 2687.860 60.300 2688.060 60.500 ;
  LAYER VI2 ;
  RECT 2687.860 59.900 2688.060 60.100 ;
  LAYER VI2 ;
  RECT 2687.860 59.500 2688.060 59.700 ;
  LAYER VI2 ;
  RECT 2687.860 59.100 2688.060 59.300 ;
  LAYER VI2 ;
  RECT 2687.860 58.700 2688.060 58.900 ;
  LAYER VI2 ;
  RECT 2687.860 58.300 2688.060 58.500 ;
  LAYER VI2 ;
  RECT 2687.860 57.900 2688.060 58.100 ;
  LAYER VI2 ;
  RECT 2687.860 57.500 2688.060 57.700 ;
  LAYER VI2 ;
  RECT 2687.860 57.100 2688.060 57.300 ;
  LAYER VI3 ;
  RECT 2686.380 5.880 2687.520 6.740 ;
  LAYER VI3 ;
  RECT 2687.180 6.340 2687.380 6.540 ;
  LAYER VI3 ;
  RECT 2687.180 5.940 2687.380 6.140 ;
  LAYER VI3 ;
  RECT 2686.780 6.340 2686.980 6.540 ;
  LAYER VI3 ;
  RECT 2686.780 5.940 2686.980 6.140 ;
  LAYER VI3 ;
  RECT 2686.380 6.340 2686.580 6.540 ;
  LAYER VI3 ;
  RECT 2686.380 5.940 2686.580 6.140 ;
  LAYER VI3 ;
  RECT 1378.180 5.880 1386.180 6.740 ;
  LAYER VI3 ;
  RECT 1385.780 6.340 1385.980 6.540 ;
  LAYER VI3 ;
  RECT 1385.780 5.940 1385.980 6.140 ;
  LAYER VI3 ;
  RECT 1385.380 6.340 1385.580 6.540 ;
  LAYER VI3 ;
  RECT 1385.380 5.940 1385.580 6.140 ;
  LAYER VI3 ;
  RECT 1384.980 6.340 1385.180 6.540 ;
  LAYER VI3 ;
  RECT 1384.980 5.940 1385.180 6.140 ;
  LAYER VI3 ;
  RECT 1384.580 6.340 1384.780 6.540 ;
  LAYER VI3 ;
  RECT 1384.580 5.940 1384.780 6.140 ;
  LAYER VI3 ;
  RECT 1384.180 6.340 1384.380 6.540 ;
  LAYER VI3 ;
  RECT 1384.180 5.940 1384.380 6.140 ;
  LAYER VI3 ;
  RECT 1383.780 6.340 1383.980 6.540 ;
  LAYER VI3 ;
  RECT 1383.780 5.940 1383.980 6.140 ;
  LAYER VI3 ;
  RECT 1383.380 6.340 1383.580 6.540 ;
  LAYER VI3 ;
  RECT 1383.380 5.940 1383.580 6.140 ;
  LAYER VI3 ;
  RECT 1382.980 6.340 1383.180 6.540 ;
  LAYER VI3 ;
  RECT 1382.980 5.940 1383.180 6.140 ;
  LAYER VI3 ;
  RECT 1382.580 6.340 1382.780 6.540 ;
  LAYER VI3 ;
  RECT 1382.580 5.940 1382.780 6.140 ;
  LAYER VI3 ;
  RECT 1382.180 6.340 1382.380 6.540 ;
  LAYER VI3 ;
  RECT 1382.180 5.940 1382.380 6.140 ;
  LAYER VI3 ;
  RECT 1381.780 6.340 1381.980 6.540 ;
  LAYER VI3 ;
  RECT 1381.780 5.940 1381.980 6.140 ;
  LAYER VI3 ;
  RECT 1381.380 6.340 1381.580 6.540 ;
  LAYER VI3 ;
  RECT 1381.380 5.940 1381.580 6.140 ;
  LAYER VI3 ;
  RECT 1380.980 6.340 1381.180 6.540 ;
  LAYER VI3 ;
  RECT 1380.980 5.940 1381.180 6.140 ;
  LAYER VI3 ;
  RECT 1380.580 6.340 1380.780 6.540 ;
  LAYER VI3 ;
  RECT 1380.580 5.940 1380.780 6.140 ;
  LAYER VI3 ;
  RECT 1380.180 6.340 1380.380 6.540 ;
  LAYER VI3 ;
  RECT 1380.180 5.940 1380.380 6.140 ;
  LAYER VI3 ;
  RECT 1379.780 6.340 1379.980 6.540 ;
  LAYER VI3 ;
  RECT 1379.780 5.940 1379.980 6.140 ;
  LAYER VI3 ;
  RECT 1379.380 6.340 1379.580 6.540 ;
  LAYER VI3 ;
  RECT 1379.380 5.940 1379.580 6.140 ;
  LAYER VI3 ;
  RECT 1378.980 6.340 1379.180 6.540 ;
  LAYER VI3 ;
  RECT 1378.980 5.940 1379.180 6.140 ;
  LAYER VI3 ;
  RECT 1378.580 6.340 1378.780 6.540 ;
  LAYER VI3 ;
  RECT 1378.580 5.940 1378.780 6.140 ;
  LAYER VI3 ;
  RECT 1378.180 6.340 1378.380 6.540 ;
  LAYER VI3 ;
  RECT 1378.180 5.940 1378.380 6.140 ;
  LAYER VI3 ;
  RECT 1398.020 5.880 1406.020 6.740 ;
  LAYER VI3 ;
  RECT 1405.620 6.340 1405.820 6.540 ;
  LAYER VI3 ;
  RECT 1405.620 5.940 1405.820 6.140 ;
  LAYER VI3 ;
  RECT 1405.220 6.340 1405.420 6.540 ;
  LAYER VI3 ;
  RECT 1405.220 5.940 1405.420 6.140 ;
  LAYER VI3 ;
  RECT 1404.820 6.340 1405.020 6.540 ;
  LAYER VI3 ;
  RECT 1404.820 5.940 1405.020 6.140 ;
  LAYER VI3 ;
  RECT 1404.420 6.340 1404.620 6.540 ;
  LAYER VI3 ;
  RECT 1404.420 5.940 1404.620 6.140 ;
  LAYER VI3 ;
  RECT 1404.020 6.340 1404.220 6.540 ;
  LAYER VI3 ;
  RECT 1404.020 5.940 1404.220 6.140 ;
  LAYER VI3 ;
  RECT 1403.620 6.340 1403.820 6.540 ;
  LAYER VI3 ;
  RECT 1403.620 5.940 1403.820 6.140 ;
  LAYER VI3 ;
  RECT 1403.220 6.340 1403.420 6.540 ;
  LAYER VI3 ;
  RECT 1403.220 5.940 1403.420 6.140 ;
  LAYER VI3 ;
  RECT 1402.820 6.340 1403.020 6.540 ;
  LAYER VI3 ;
  RECT 1402.820 5.940 1403.020 6.140 ;
  LAYER VI3 ;
  RECT 1402.420 6.340 1402.620 6.540 ;
  LAYER VI3 ;
  RECT 1402.420 5.940 1402.620 6.140 ;
  LAYER VI3 ;
  RECT 1402.020 6.340 1402.220 6.540 ;
  LAYER VI3 ;
  RECT 1402.020 5.940 1402.220 6.140 ;
  LAYER VI3 ;
  RECT 1401.620 6.340 1401.820 6.540 ;
  LAYER VI3 ;
  RECT 1401.620 5.940 1401.820 6.140 ;
  LAYER VI3 ;
  RECT 1401.220 6.340 1401.420 6.540 ;
  LAYER VI3 ;
  RECT 1401.220 5.940 1401.420 6.140 ;
  LAYER VI3 ;
  RECT 1400.820 6.340 1401.020 6.540 ;
  LAYER VI3 ;
  RECT 1400.820 5.940 1401.020 6.140 ;
  LAYER VI3 ;
  RECT 1400.420 6.340 1400.620 6.540 ;
  LAYER VI3 ;
  RECT 1400.420 5.940 1400.620 6.140 ;
  LAYER VI3 ;
  RECT 1400.020 6.340 1400.220 6.540 ;
  LAYER VI3 ;
  RECT 1400.020 5.940 1400.220 6.140 ;
  LAYER VI3 ;
  RECT 1399.620 6.340 1399.820 6.540 ;
  LAYER VI3 ;
  RECT 1399.620 5.940 1399.820 6.140 ;
  LAYER VI3 ;
  RECT 1399.220 6.340 1399.420 6.540 ;
  LAYER VI3 ;
  RECT 1399.220 5.940 1399.420 6.140 ;
  LAYER VI3 ;
  RECT 1398.820 6.340 1399.020 6.540 ;
  LAYER VI3 ;
  RECT 1398.820 5.940 1399.020 6.140 ;
  LAYER VI3 ;
  RECT 1398.420 6.340 1398.620 6.540 ;
  LAYER VI3 ;
  RECT 1398.420 5.940 1398.620 6.140 ;
  LAYER VI3 ;
  RECT 1398.020 6.340 1398.220 6.540 ;
  LAYER VI3 ;
  RECT 1398.020 5.940 1398.220 6.140 ;
  LAYER VI3 ;
  RECT 1419.100 5.880 1427.100 6.740 ;
  LAYER VI3 ;
  RECT 1426.700 6.340 1426.900 6.540 ;
  LAYER VI3 ;
  RECT 1426.700 5.940 1426.900 6.140 ;
  LAYER VI3 ;
  RECT 1426.300 6.340 1426.500 6.540 ;
  LAYER VI3 ;
  RECT 1426.300 5.940 1426.500 6.140 ;
  LAYER VI3 ;
  RECT 1425.900 6.340 1426.100 6.540 ;
  LAYER VI3 ;
  RECT 1425.900 5.940 1426.100 6.140 ;
  LAYER VI3 ;
  RECT 1425.500 6.340 1425.700 6.540 ;
  LAYER VI3 ;
  RECT 1425.500 5.940 1425.700 6.140 ;
  LAYER VI3 ;
  RECT 1425.100 6.340 1425.300 6.540 ;
  LAYER VI3 ;
  RECT 1425.100 5.940 1425.300 6.140 ;
  LAYER VI3 ;
  RECT 1424.700 6.340 1424.900 6.540 ;
  LAYER VI3 ;
  RECT 1424.700 5.940 1424.900 6.140 ;
  LAYER VI3 ;
  RECT 1424.300 6.340 1424.500 6.540 ;
  LAYER VI3 ;
  RECT 1424.300 5.940 1424.500 6.140 ;
  LAYER VI3 ;
  RECT 1423.900 6.340 1424.100 6.540 ;
  LAYER VI3 ;
  RECT 1423.900 5.940 1424.100 6.140 ;
  LAYER VI3 ;
  RECT 1423.500 6.340 1423.700 6.540 ;
  LAYER VI3 ;
  RECT 1423.500 5.940 1423.700 6.140 ;
  LAYER VI3 ;
  RECT 1423.100 6.340 1423.300 6.540 ;
  LAYER VI3 ;
  RECT 1423.100 5.940 1423.300 6.140 ;
  LAYER VI3 ;
  RECT 1422.700 6.340 1422.900 6.540 ;
  LAYER VI3 ;
  RECT 1422.700 5.940 1422.900 6.140 ;
  LAYER VI3 ;
  RECT 1422.300 6.340 1422.500 6.540 ;
  LAYER VI3 ;
  RECT 1422.300 5.940 1422.500 6.140 ;
  LAYER VI3 ;
  RECT 1421.900 6.340 1422.100 6.540 ;
  LAYER VI3 ;
  RECT 1421.900 5.940 1422.100 6.140 ;
  LAYER VI3 ;
  RECT 1421.500 6.340 1421.700 6.540 ;
  LAYER VI3 ;
  RECT 1421.500 5.940 1421.700 6.140 ;
  LAYER VI3 ;
  RECT 1421.100 6.340 1421.300 6.540 ;
  LAYER VI3 ;
  RECT 1421.100 5.940 1421.300 6.140 ;
  LAYER VI3 ;
  RECT 1420.700 6.340 1420.900 6.540 ;
  LAYER VI3 ;
  RECT 1420.700 5.940 1420.900 6.140 ;
  LAYER VI3 ;
  RECT 1420.300 6.340 1420.500 6.540 ;
  LAYER VI3 ;
  RECT 1420.300 5.940 1420.500 6.140 ;
  LAYER VI3 ;
  RECT 1419.900 6.340 1420.100 6.540 ;
  LAYER VI3 ;
  RECT 1419.900 5.940 1420.100 6.140 ;
  LAYER VI3 ;
  RECT 1419.500 6.340 1419.700 6.540 ;
  LAYER VI3 ;
  RECT 1419.500 5.940 1419.700 6.140 ;
  LAYER VI3 ;
  RECT 1419.100 6.340 1419.300 6.540 ;
  LAYER VI3 ;
  RECT 1419.100 5.940 1419.300 6.140 ;
  LAYER VI3 ;
  RECT 1438.940 5.880 1446.940 6.740 ;
  LAYER VI3 ;
  RECT 1446.540 6.340 1446.740 6.540 ;
  LAYER VI3 ;
  RECT 1446.540 5.940 1446.740 6.140 ;
  LAYER VI3 ;
  RECT 1446.140 6.340 1446.340 6.540 ;
  LAYER VI3 ;
  RECT 1446.140 5.940 1446.340 6.140 ;
  LAYER VI3 ;
  RECT 1445.740 6.340 1445.940 6.540 ;
  LAYER VI3 ;
  RECT 1445.740 5.940 1445.940 6.140 ;
  LAYER VI3 ;
  RECT 1445.340 6.340 1445.540 6.540 ;
  LAYER VI3 ;
  RECT 1445.340 5.940 1445.540 6.140 ;
  LAYER VI3 ;
  RECT 1444.940 6.340 1445.140 6.540 ;
  LAYER VI3 ;
  RECT 1444.940 5.940 1445.140 6.140 ;
  LAYER VI3 ;
  RECT 1444.540 6.340 1444.740 6.540 ;
  LAYER VI3 ;
  RECT 1444.540 5.940 1444.740 6.140 ;
  LAYER VI3 ;
  RECT 1444.140 6.340 1444.340 6.540 ;
  LAYER VI3 ;
  RECT 1444.140 5.940 1444.340 6.140 ;
  LAYER VI3 ;
  RECT 1443.740 6.340 1443.940 6.540 ;
  LAYER VI3 ;
  RECT 1443.740 5.940 1443.940 6.140 ;
  LAYER VI3 ;
  RECT 1443.340 6.340 1443.540 6.540 ;
  LAYER VI3 ;
  RECT 1443.340 5.940 1443.540 6.140 ;
  LAYER VI3 ;
  RECT 1442.940 6.340 1443.140 6.540 ;
  LAYER VI3 ;
  RECT 1442.940 5.940 1443.140 6.140 ;
  LAYER VI3 ;
  RECT 1442.540 6.340 1442.740 6.540 ;
  LAYER VI3 ;
  RECT 1442.540 5.940 1442.740 6.140 ;
  LAYER VI3 ;
  RECT 1442.140 6.340 1442.340 6.540 ;
  LAYER VI3 ;
  RECT 1442.140 5.940 1442.340 6.140 ;
  LAYER VI3 ;
  RECT 1441.740 6.340 1441.940 6.540 ;
  LAYER VI3 ;
  RECT 1441.740 5.940 1441.940 6.140 ;
  LAYER VI3 ;
  RECT 1441.340 6.340 1441.540 6.540 ;
  LAYER VI3 ;
  RECT 1441.340 5.940 1441.540 6.140 ;
  LAYER VI3 ;
  RECT 1440.940 6.340 1441.140 6.540 ;
  LAYER VI3 ;
  RECT 1440.940 5.940 1441.140 6.140 ;
  LAYER VI3 ;
  RECT 1440.540 6.340 1440.740 6.540 ;
  LAYER VI3 ;
  RECT 1440.540 5.940 1440.740 6.140 ;
  LAYER VI3 ;
  RECT 1440.140 6.340 1440.340 6.540 ;
  LAYER VI3 ;
  RECT 1440.140 5.940 1440.340 6.140 ;
  LAYER VI3 ;
  RECT 1439.740 6.340 1439.940 6.540 ;
  LAYER VI3 ;
  RECT 1439.740 5.940 1439.940 6.140 ;
  LAYER VI3 ;
  RECT 1439.340 6.340 1439.540 6.540 ;
  LAYER VI3 ;
  RECT 1439.340 5.940 1439.540 6.140 ;
  LAYER VI3 ;
  RECT 1438.940 6.340 1439.140 6.540 ;
  LAYER VI3 ;
  RECT 1438.940 5.940 1439.140 6.140 ;
  LAYER VI3 ;
  RECT 1460.020 5.880 1468.020 6.740 ;
  LAYER VI3 ;
  RECT 1467.620 6.340 1467.820 6.540 ;
  LAYER VI3 ;
  RECT 1467.620 5.940 1467.820 6.140 ;
  LAYER VI3 ;
  RECT 1467.220 6.340 1467.420 6.540 ;
  LAYER VI3 ;
  RECT 1467.220 5.940 1467.420 6.140 ;
  LAYER VI3 ;
  RECT 1466.820 6.340 1467.020 6.540 ;
  LAYER VI3 ;
  RECT 1466.820 5.940 1467.020 6.140 ;
  LAYER VI3 ;
  RECT 1466.420 6.340 1466.620 6.540 ;
  LAYER VI3 ;
  RECT 1466.420 5.940 1466.620 6.140 ;
  LAYER VI3 ;
  RECT 1466.020 6.340 1466.220 6.540 ;
  LAYER VI3 ;
  RECT 1466.020 5.940 1466.220 6.140 ;
  LAYER VI3 ;
  RECT 1465.620 6.340 1465.820 6.540 ;
  LAYER VI3 ;
  RECT 1465.620 5.940 1465.820 6.140 ;
  LAYER VI3 ;
  RECT 1465.220 6.340 1465.420 6.540 ;
  LAYER VI3 ;
  RECT 1465.220 5.940 1465.420 6.140 ;
  LAYER VI3 ;
  RECT 1464.820 6.340 1465.020 6.540 ;
  LAYER VI3 ;
  RECT 1464.820 5.940 1465.020 6.140 ;
  LAYER VI3 ;
  RECT 1464.420 6.340 1464.620 6.540 ;
  LAYER VI3 ;
  RECT 1464.420 5.940 1464.620 6.140 ;
  LAYER VI3 ;
  RECT 1464.020 6.340 1464.220 6.540 ;
  LAYER VI3 ;
  RECT 1464.020 5.940 1464.220 6.140 ;
  LAYER VI3 ;
  RECT 1463.620 6.340 1463.820 6.540 ;
  LAYER VI3 ;
  RECT 1463.620 5.940 1463.820 6.140 ;
  LAYER VI3 ;
  RECT 1463.220 6.340 1463.420 6.540 ;
  LAYER VI3 ;
  RECT 1463.220 5.940 1463.420 6.140 ;
  LAYER VI3 ;
  RECT 1462.820 6.340 1463.020 6.540 ;
  LAYER VI3 ;
  RECT 1462.820 5.940 1463.020 6.140 ;
  LAYER VI3 ;
  RECT 1462.420 6.340 1462.620 6.540 ;
  LAYER VI3 ;
  RECT 1462.420 5.940 1462.620 6.140 ;
  LAYER VI3 ;
  RECT 1462.020 6.340 1462.220 6.540 ;
  LAYER VI3 ;
  RECT 1462.020 5.940 1462.220 6.140 ;
  LAYER VI3 ;
  RECT 1461.620 6.340 1461.820 6.540 ;
  LAYER VI3 ;
  RECT 1461.620 5.940 1461.820 6.140 ;
  LAYER VI3 ;
  RECT 1461.220 6.340 1461.420 6.540 ;
  LAYER VI3 ;
  RECT 1461.220 5.940 1461.420 6.140 ;
  LAYER VI3 ;
  RECT 1460.820 6.340 1461.020 6.540 ;
  LAYER VI3 ;
  RECT 1460.820 5.940 1461.020 6.140 ;
  LAYER VI3 ;
  RECT 1460.420 6.340 1460.620 6.540 ;
  LAYER VI3 ;
  RECT 1460.420 5.940 1460.620 6.140 ;
  LAYER VI3 ;
  RECT 1460.020 6.340 1460.220 6.540 ;
  LAYER VI3 ;
  RECT 1460.020 5.940 1460.220 6.140 ;
  LAYER VI3 ;
  RECT 1479.860 5.880 1487.860 6.740 ;
  LAYER VI3 ;
  RECT 1487.460 6.340 1487.660 6.540 ;
  LAYER VI3 ;
  RECT 1487.460 5.940 1487.660 6.140 ;
  LAYER VI3 ;
  RECT 1487.060 6.340 1487.260 6.540 ;
  LAYER VI3 ;
  RECT 1487.060 5.940 1487.260 6.140 ;
  LAYER VI3 ;
  RECT 1486.660 6.340 1486.860 6.540 ;
  LAYER VI3 ;
  RECT 1486.660 5.940 1486.860 6.140 ;
  LAYER VI3 ;
  RECT 1486.260 6.340 1486.460 6.540 ;
  LAYER VI3 ;
  RECT 1486.260 5.940 1486.460 6.140 ;
  LAYER VI3 ;
  RECT 1485.860 6.340 1486.060 6.540 ;
  LAYER VI3 ;
  RECT 1485.860 5.940 1486.060 6.140 ;
  LAYER VI3 ;
  RECT 1485.460 6.340 1485.660 6.540 ;
  LAYER VI3 ;
  RECT 1485.460 5.940 1485.660 6.140 ;
  LAYER VI3 ;
  RECT 1485.060 6.340 1485.260 6.540 ;
  LAYER VI3 ;
  RECT 1485.060 5.940 1485.260 6.140 ;
  LAYER VI3 ;
  RECT 1484.660 6.340 1484.860 6.540 ;
  LAYER VI3 ;
  RECT 1484.660 5.940 1484.860 6.140 ;
  LAYER VI3 ;
  RECT 1484.260 6.340 1484.460 6.540 ;
  LAYER VI3 ;
  RECT 1484.260 5.940 1484.460 6.140 ;
  LAYER VI3 ;
  RECT 1483.860 6.340 1484.060 6.540 ;
  LAYER VI3 ;
  RECT 1483.860 5.940 1484.060 6.140 ;
  LAYER VI3 ;
  RECT 1483.460 6.340 1483.660 6.540 ;
  LAYER VI3 ;
  RECT 1483.460 5.940 1483.660 6.140 ;
  LAYER VI3 ;
  RECT 1483.060 6.340 1483.260 6.540 ;
  LAYER VI3 ;
  RECT 1483.060 5.940 1483.260 6.140 ;
  LAYER VI3 ;
  RECT 1482.660 6.340 1482.860 6.540 ;
  LAYER VI3 ;
  RECT 1482.660 5.940 1482.860 6.140 ;
  LAYER VI3 ;
  RECT 1482.260 6.340 1482.460 6.540 ;
  LAYER VI3 ;
  RECT 1482.260 5.940 1482.460 6.140 ;
  LAYER VI3 ;
  RECT 1481.860 6.340 1482.060 6.540 ;
  LAYER VI3 ;
  RECT 1481.860 5.940 1482.060 6.140 ;
  LAYER VI3 ;
  RECT 1481.460 6.340 1481.660 6.540 ;
  LAYER VI3 ;
  RECT 1481.460 5.940 1481.660 6.140 ;
  LAYER VI3 ;
  RECT 1481.060 6.340 1481.260 6.540 ;
  LAYER VI3 ;
  RECT 1481.060 5.940 1481.260 6.140 ;
  LAYER VI3 ;
  RECT 1480.660 6.340 1480.860 6.540 ;
  LAYER VI3 ;
  RECT 1480.660 5.940 1480.860 6.140 ;
  LAYER VI3 ;
  RECT 1480.260 6.340 1480.460 6.540 ;
  LAYER VI3 ;
  RECT 1480.260 5.940 1480.460 6.140 ;
  LAYER VI3 ;
  RECT 1479.860 6.340 1480.060 6.540 ;
  LAYER VI3 ;
  RECT 1479.860 5.940 1480.060 6.140 ;
  LAYER VI3 ;
  RECT 1500.940 5.880 1508.940 6.740 ;
  LAYER VI3 ;
  RECT 1508.540 6.340 1508.740 6.540 ;
  LAYER VI3 ;
  RECT 1508.540 5.940 1508.740 6.140 ;
  LAYER VI3 ;
  RECT 1508.140 6.340 1508.340 6.540 ;
  LAYER VI3 ;
  RECT 1508.140 5.940 1508.340 6.140 ;
  LAYER VI3 ;
  RECT 1507.740 6.340 1507.940 6.540 ;
  LAYER VI3 ;
  RECT 1507.740 5.940 1507.940 6.140 ;
  LAYER VI3 ;
  RECT 1507.340 6.340 1507.540 6.540 ;
  LAYER VI3 ;
  RECT 1507.340 5.940 1507.540 6.140 ;
  LAYER VI3 ;
  RECT 1506.940 6.340 1507.140 6.540 ;
  LAYER VI3 ;
  RECT 1506.940 5.940 1507.140 6.140 ;
  LAYER VI3 ;
  RECT 1506.540 6.340 1506.740 6.540 ;
  LAYER VI3 ;
  RECT 1506.540 5.940 1506.740 6.140 ;
  LAYER VI3 ;
  RECT 1506.140 6.340 1506.340 6.540 ;
  LAYER VI3 ;
  RECT 1506.140 5.940 1506.340 6.140 ;
  LAYER VI3 ;
  RECT 1505.740 6.340 1505.940 6.540 ;
  LAYER VI3 ;
  RECT 1505.740 5.940 1505.940 6.140 ;
  LAYER VI3 ;
  RECT 1505.340 6.340 1505.540 6.540 ;
  LAYER VI3 ;
  RECT 1505.340 5.940 1505.540 6.140 ;
  LAYER VI3 ;
  RECT 1504.940 6.340 1505.140 6.540 ;
  LAYER VI3 ;
  RECT 1504.940 5.940 1505.140 6.140 ;
  LAYER VI3 ;
  RECT 1504.540 6.340 1504.740 6.540 ;
  LAYER VI3 ;
  RECT 1504.540 5.940 1504.740 6.140 ;
  LAYER VI3 ;
  RECT 1504.140 6.340 1504.340 6.540 ;
  LAYER VI3 ;
  RECT 1504.140 5.940 1504.340 6.140 ;
  LAYER VI3 ;
  RECT 1503.740 6.340 1503.940 6.540 ;
  LAYER VI3 ;
  RECT 1503.740 5.940 1503.940 6.140 ;
  LAYER VI3 ;
  RECT 1503.340 6.340 1503.540 6.540 ;
  LAYER VI3 ;
  RECT 1503.340 5.940 1503.540 6.140 ;
  LAYER VI3 ;
  RECT 1502.940 6.340 1503.140 6.540 ;
  LAYER VI3 ;
  RECT 1502.940 5.940 1503.140 6.140 ;
  LAYER VI3 ;
  RECT 1502.540 6.340 1502.740 6.540 ;
  LAYER VI3 ;
  RECT 1502.540 5.940 1502.740 6.140 ;
  LAYER VI3 ;
  RECT 1502.140 6.340 1502.340 6.540 ;
  LAYER VI3 ;
  RECT 1502.140 5.940 1502.340 6.140 ;
  LAYER VI3 ;
  RECT 1501.740 6.340 1501.940 6.540 ;
  LAYER VI3 ;
  RECT 1501.740 5.940 1501.940 6.140 ;
  LAYER VI3 ;
  RECT 1501.340 6.340 1501.540 6.540 ;
  LAYER VI3 ;
  RECT 1501.340 5.940 1501.540 6.140 ;
  LAYER VI3 ;
  RECT 1500.940 6.340 1501.140 6.540 ;
  LAYER VI3 ;
  RECT 1500.940 5.940 1501.140 6.140 ;
  LAYER VI3 ;
  RECT 1520.780 5.880 1528.780 6.740 ;
  LAYER VI3 ;
  RECT 1528.380 6.340 1528.580 6.540 ;
  LAYER VI3 ;
  RECT 1528.380 5.940 1528.580 6.140 ;
  LAYER VI3 ;
  RECT 1527.980 6.340 1528.180 6.540 ;
  LAYER VI3 ;
  RECT 1527.980 5.940 1528.180 6.140 ;
  LAYER VI3 ;
  RECT 1527.580 6.340 1527.780 6.540 ;
  LAYER VI3 ;
  RECT 1527.580 5.940 1527.780 6.140 ;
  LAYER VI3 ;
  RECT 1527.180 6.340 1527.380 6.540 ;
  LAYER VI3 ;
  RECT 1527.180 5.940 1527.380 6.140 ;
  LAYER VI3 ;
  RECT 1526.780 6.340 1526.980 6.540 ;
  LAYER VI3 ;
  RECT 1526.780 5.940 1526.980 6.140 ;
  LAYER VI3 ;
  RECT 1526.380 6.340 1526.580 6.540 ;
  LAYER VI3 ;
  RECT 1526.380 5.940 1526.580 6.140 ;
  LAYER VI3 ;
  RECT 1525.980 6.340 1526.180 6.540 ;
  LAYER VI3 ;
  RECT 1525.980 5.940 1526.180 6.140 ;
  LAYER VI3 ;
  RECT 1525.580 6.340 1525.780 6.540 ;
  LAYER VI3 ;
  RECT 1525.580 5.940 1525.780 6.140 ;
  LAYER VI3 ;
  RECT 1525.180 6.340 1525.380 6.540 ;
  LAYER VI3 ;
  RECT 1525.180 5.940 1525.380 6.140 ;
  LAYER VI3 ;
  RECT 1524.780 6.340 1524.980 6.540 ;
  LAYER VI3 ;
  RECT 1524.780 5.940 1524.980 6.140 ;
  LAYER VI3 ;
  RECT 1524.380 6.340 1524.580 6.540 ;
  LAYER VI3 ;
  RECT 1524.380 5.940 1524.580 6.140 ;
  LAYER VI3 ;
  RECT 1523.980 6.340 1524.180 6.540 ;
  LAYER VI3 ;
  RECT 1523.980 5.940 1524.180 6.140 ;
  LAYER VI3 ;
  RECT 1523.580 6.340 1523.780 6.540 ;
  LAYER VI3 ;
  RECT 1523.580 5.940 1523.780 6.140 ;
  LAYER VI3 ;
  RECT 1523.180 6.340 1523.380 6.540 ;
  LAYER VI3 ;
  RECT 1523.180 5.940 1523.380 6.140 ;
  LAYER VI3 ;
  RECT 1522.780 6.340 1522.980 6.540 ;
  LAYER VI3 ;
  RECT 1522.780 5.940 1522.980 6.140 ;
  LAYER VI3 ;
  RECT 1522.380 6.340 1522.580 6.540 ;
  LAYER VI3 ;
  RECT 1522.380 5.940 1522.580 6.140 ;
  LAYER VI3 ;
  RECT 1521.980 6.340 1522.180 6.540 ;
  LAYER VI3 ;
  RECT 1521.980 5.940 1522.180 6.140 ;
  LAYER VI3 ;
  RECT 1521.580 6.340 1521.780 6.540 ;
  LAYER VI3 ;
  RECT 1521.580 5.940 1521.780 6.140 ;
  LAYER VI3 ;
  RECT 1521.180 6.340 1521.380 6.540 ;
  LAYER VI3 ;
  RECT 1521.180 5.940 1521.380 6.140 ;
  LAYER VI3 ;
  RECT 1520.780 6.340 1520.980 6.540 ;
  LAYER VI3 ;
  RECT 1520.780 5.940 1520.980 6.140 ;
  LAYER VI3 ;
  RECT 1541.860 5.880 1549.860 6.740 ;
  LAYER VI3 ;
  RECT 1549.460 6.340 1549.660 6.540 ;
  LAYER VI3 ;
  RECT 1549.460 5.940 1549.660 6.140 ;
  LAYER VI3 ;
  RECT 1549.060 6.340 1549.260 6.540 ;
  LAYER VI3 ;
  RECT 1549.060 5.940 1549.260 6.140 ;
  LAYER VI3 ;
  RECT 1548.660 6.340 1548.860 6.540 ;
  LAYER VI3 ;
  RECT 1548.660 5.940 1548.860 6.140 ;
  LAYER VI3 ;
  RECT 1548.260 6.340 1548.460 6.540 ;
  LAYER VI3 ;
  RECT 1548.260 5.940 1548.460 6.140 ;
  LAYER VI3 ;
  RECT 1547.860 6.340 1548.060 6.540 ;
  LAYER VI3 ;
  RECT 1547.860 5.940 1548.060 6.140 ;
  LAYER VI3 ;
  RECT 1547.460 6.340 1547.660 6.540 ;
  LAYER VI3 ;
  RECT 1547.460 5.940 1547.660 6.140 ;
  LAYER VI3 ;
  RECT 1547.060 6.340 1547.260 6.540 ;
  LAYER VI3 ;
  RECT 1547.060 5.940 1547.260 6.140 ;
  LAYER VI3 ;
  RECT 1546.660 6.340 1546.860 6.540 ;
  LAYER VI3 ;
  RECT 1546.660 5.940 1546.860 6.140 ;
  LAYER VI3 ;
  RECT 1546.260 6.340 1546.460 6.540 ;
  LAYER VI3 ;
  RECT 1546.260 5.940 1546.460 6.140 ;
  LAYER VI3 ;
  RECT 1545.860 6.340 1546.060 6.540 ;
  LAYER VI3 ;
  RECT 1545.860 5.940 1546.060 6.140 ;
  LAYER VI3 ;
  RECT 1545.460 6.340 1545.660 6.540 ;
  LAYER VI3 ;
  RECT 1545.460 5.940 1545.660 6.140 ;
  LAYER VI3 ;
  RECT 1545.060 6.340 1545.260 6.540 ;
  LAYER VI3 ;
  RECT 1545.060 5.940 1545.260 6.140 ;
  LAYER VI3 ;
  RECT 1544.660 6.340 1544.860 6.540 ;
  LAYER VI3 ;
  RECT 1544.660 5.940 1544.860 6.140 ;
  LAYER VI3 ;
  RECT 1544.260 6.340 1544.460 6.540 ;
  LAYER VI3 ;
  RECT 1544.260 5.940 1544.460 6.140 ;
  LAYER VI3 ;
  RECT 1543.860 6.340 1544.060 6.540 ;
  LAYER VI3 ;
  RECT 1543.860 5.940 1544.060 6.140 ;
  LAYER VI3 ;
  RECT 1543.460 6.340 1543.660 6.540 ;
  LAYER VI3 ;
  RECT 1543.460 5.940 1543.660 6.140 ;
  LAYER VI3 ;
  RECT 1543.060 6.340 1543.260 6.540 ;
  LAYER VI3 ;
  RECT 1543.060 5.940 1543.260 6.140 ;
  LAYER VI3 ;
  RECT 1542.660 6.340 1542.860 6.540 ;
  LAYER VI3 ;
  RECT 1542.660 5.940 1542.860 6.140 ;
  LAYER VI3 ;
  RECT 1542.260 6.340 1542.460 6.540 ;
  LAYER VI3 ;
  RECT 1542.260 5.940 1542.460 6.140 ;
  LAYER VI3 ;
  RECT 1541.860 6.340 1542.060 6.540 ;
  LAYER VI3 ;
  RECT 1541.860 5.940 1542.060 6.140 ;
  LAYER VI3 ;
  RECT 1561.700 5.880 1569.700 6.740 ;
  LAYER VI3 ;
  RECT 1569.300 6.340 1569.500 6.540 ;
  LAYER VI3 ;
  RECT 1569.300 5.940 1569.500 6.140 ;
  LAYER VI3 ;
  RECT 1568.900 6.340 1569.100 6.540 ;
  LAYER VI3 ;
  RECT 1568.900 5.940 1569.100 6.140 ;
  LAYER VI3 ;
  RECT 1568.500 6.340 1568.700 6.540 ;
  LAYER VI3 ;
  RECT 1568.500 5.940 1568.700 6.140 ;
  LAYER VI3 ;
  RECT 1568.100 6.340 1568.300 6.540 ;
  LAYER VI3 ;
  RECT 1568.100 5.940 1568.300 6.140 ;
  LAYER VI3 ;
  RECT 1567.700 6.340 1567.900 6.540 ;
  LAYER VI3 ;
  RECT 1567.700 5.940 1567.900 6.140 ;
  LAYER VI3 ;
  RECT 1567.300 6.340 1567.500 6.540 ;
  LAYER VI3 ;
  RECT 1567.300 5.940 1567.500 6.140 ;
  LAYER VI3 ;
  RECT 1566.900 6.340 1567.100 6.540 ;
  LAYER VI3 ;
  RECT 1566.900 5.940 1567.100 6.140 ;
  LAYER VI3 ;
  RECT 1566.500 6.340 1566.700 6.540 ;
  LAYER VI3 ;
  RECT 1566.500 5.940 1566.700 6.140 ;
  LAYER VI3 ;
  RECT 1566.100 6.340 1566.300 6.540 ;
  LAYER VI3 ;
  RECT 1566.100 5.940 1566.300 6.140 ;
  LAYER VI3 ;
  RECT 1565.700 6.340 1565.900 6.540 ;
  LAYER VI3 ;
  RECT 1565.700 5.940 1565.900 6.140 ;
  LAYER VI3 ;
  RECT 1565.300 6.340 1565.500 6.540 ;
  LAYER VI3 ;
  RECT 1565.300 5.940 1565.500 6.140 ;
  LAYER VI3 ;
  RECT 1564.900 6.340 1565.100 6.540 ;
  LAYER VI3 ;
  RECT 1564.900 5.940 1565.100 6.140 ;
  LAYER VI3 ;
  RECT 1564.500 6.340 1564.700 6.540 ;
  LAYER VI3 ;
  RECT 1564.500 5.940 1564.700 6.140 ;
  LAYER VI3 ;
  RECT 1564.100 6.340 1564.300 6.540 ;
  LAYER VI3 ;
  RECT 1564.100 5.940 1564.300 6.140 ;
  LAYER VI3 ;
  RECT 1563.700 6.340 1563.900 6.540 ;
  LAYER VI3 ;
  RECT 1563.700 5.940 1563.900 6.140 ;
  LAYER VI3 ;
  RECT 1563.300 6.340 1563.500 6.540 ;
  LAYER VI3 ;
  RECT 1563.300 5.940 1563.500 6.140 ;
  LAYER VI3 ;
  RECT 1562.900 6.340 1563.100 6.540 ;
  LAYER VI3 ;
  RECT 1562.900 5.940 1563.100 6.140 ;
  LAYER VI3 ;
  RECT 1562.500 6.340 1562.700 6.540 ;
  LAYER VI3 ;
  RECT 1562.500 5.940 1562.700 6.140 ;
  LAYER VI3 ;
  RECT 1562.100 6.340 1562.300 6.540 ;
  LAYER VI3 ;
  RECT 1562.100 5.940 1562.300 6.140 ;
  LAYER VI3 ;
  RECT 1561.700 6.340 1561.900 6.540 ;
  LAYER VI3 ;
  RECT 1561.700 5.940 1561.900 6.140 ;
  LAYER VI3 ;
  RECT 1582.780 5.880 1590.780 6.740 ;
  LAYER VI3 ;
  RECT 1590.380 6.340 1590.580 6.540 ;
  LAYER VI3 ;
  RECT 1590.380 5.940 1590.580 6.140 ;
  LAYER VI3 ;
  RECT 1589.980 6.340 1590.180 6.540 ;
  LAYER VI3 ;
  RECT 1589.980 5.940 1590.180 6.140 ;
  LAYER VI3 ;
  RECT 1589.580 6.340 1589.780 6.540 ;
  LAYER VI3 ;
  RECT 1589.580 5.940 1589.780 6.140 ;
  LAYER VI3 ;
  RECT 1589.180 6.340 1589.380 6.540 ;
  LAYER VI3 ;
  RECT 1589.180 5.940 1589.380 6.140 ;
  LAYER VI3 ;
  RECT 1588.780 6.340 1588.980 6.540 ;
  LAYER VI3 ;
  RECT 1588.780 5.940 1588.980 6.140 ;
  LAYER VI3 ;
  RECT 1588.380 6.340 1588.580 6.540 ;
  LAYER VI3 ;
  RECT 1588.380 5.940 1588.580 6.140 ;
  LAYER VI3 ;
  RECT 1587.980 6.340 1588.180 6.540 ;
  LAYER VI3 ;
  RECT 1587.980 5.940 1588.180 6.140 ;
  LAYER VI3 ;
  RECT 1587.580 6.340 1587.780 6.540 ;
  LAYER VI3 ;
  RECT 1587.580 5.940 1587.780 6.140 ;
  LAYER VI3 ;
  RECT 1587.180 6.340 1587.380 6.540 ;
  LAYER VI3 ;
  RECT 1587.180 5.940 1587.380 6.140 ;
  LAYER VI3 ;
  RECT 1586.780 6.340 1586.980 6.540 ;
  LAYER VI3 ;
  RECT 1586.780 5.940 1586.980 6.140 ;
  LAYER VI3 ;
  RECT 1586.380 6.340 1586.580 6.540 ;
  LAYER VI3 ;
  RECT 1586.380 5.940 1586.580 6.140 ;
  LAYER VI3 ;
  RECT 1585.980 6.340 1586.180 6.540 ;
  LAYER VI3 ;
  RECT 1585.980 5.940 1586.180 6.140 ;
  LAYER VI3 ;
  RECT 1585.580 6.340 1585.780 6.540 ;
  LAYER VI3 ;
  RECT 1585.580 5.940 1585.780 6.140 ;
  LAYER VI3 ;
  RECT 1585.180 6.340 1585.380 6.540 ;
  LAYER VI3 ;
  RECT 1585.180 5.940 1585.380 6.140 ;
  LAYER VI3 ;
  RECT 1584.780 6.340 1584.980 6.540 ;
  LAYER VI3 ;
  RECT 1584.780 5.940 1584.980 6.140 ;
  LAYER VI3 ;
  RECT 1584.380 6.340 1584.580 6.540 ;
  LAYER VI3 ;
  RECT 1584.380 5.940 1584.580 6.140 ;
  LAYER VI3 ;
  RECT 1583.980 6.340 1584.180 6.540 ;
  LAYER VI3 ;
  RECT 1583.980 5.940 1584.180 6.140 ;
  LAYER VI3 ;
  RECT 1583.580 6.340 1583.780 6.540 ;
  LAYER VI3 ;
  RECT 1583.580 5.940 1583.780 6.140 ;
  LAYER VI3 ;
  RECT 1583.180 6.340 1583.380 6.540 ;
  LAYER VI3 ;
  RECT 1583.180 5.940 1583.380 6.140 ;
  LAYER VI3 ;
  RECT 1582.780 6.340 1582.980 6.540 ;
  LAYER VI3 ;
  RECT 1582.780 5.940 1582.980 6.140 ;
  LAYER VI3 ;
  RECT 1602.620 5.880 1610.620 6.740 ;
  LAYER VI3 ;
  RECT 1610.220 6.340 1610.420 6.540 ;
  LAYER VI3 ;
  RECT 1610.220 5.940 1610.420 6.140 ;
  LAYER VI3 ;
  RECT 1609.820 6.340 1610.020 6.540 ;
  LAYER VI3 ;
  RECT 1609.820 5.940 1610.020 6.140 ;
  LAYER VI3 ;
  RECT 1609.420 6.340 1609.620 6.540 ;
  LAYER VI3 ;
  RECT 1609.420 5.940 1609.620 6.140 ;
  LAYER VI3 ;
  RECT 1609.020 6.340 1609.220 6.540 ;
  LAYER VI3 ;
  RECT 1609.020 5.940 1609.220 6.140 ;
  LAYER VI3 ;
  RECT 1608.620 6.340 1608.820 6.540 ;
  LAYER VI3 ;
  RECT 1608.620 5.940 1608.820 6.140 ;
  LAYER VI3 ;
  RECT 1608.220 6.340 1608.420 6.540 ;
  LAYER VI3 ;
  RECT 1608.220 5.940 1608.420 6.140 ;
  LAYER VI3 ;
  RECT 1607.820 6.340 1608.020 6.540 ;
  LAYER VI3 ;
  RECT 1607.820 5.940 1608.020 6.140 ;
  LAYER VI3 ;
  RECT 1607.420 6.340 1607.620 6.540 ;
  LAYER VI3 ;
  RECT 1607.420 5.940 1607.620 6.140 ;
  LAYER VI3 ;
  RECT 1607.020 6.340 1607.220 6.540 ;
  LAYER VI3 ;
  RECT 1607.020 5.940 1607.220 6.140 ;
  LAYER VI3 ;
  RECT 1606.620 6.340 1606.820 6.540 ;
  LAYER VI3 ;
  RECT 1606.620 5.940 1606.820 6.140 ;
  LAYER VI3 ;
  RECT 1606.220 6.340 1606.420 6.540 ;
  LAYER VI3 ;
  RECT 1606.220 5.940 1606.420 6.140 ;
  LAYER VI3 ;
  RECT 1605.820 6.340 1606.020 6.540 ;
  LAYER VI3 ;
  RECT 1605.820 5.940 1606.020 6.140 ;
  LAYER VI3 ;
  RECT 1605.420 6.340 1605.620 6.540 ;
  LAYER VI3 ;
  RECT 1605.420 5.940 1605.620 6.140 ;
  LAYER VI3 ;
  RECT 1605.020 6.340 1605.220 6.540 ;
  LAYER VI3 ;
  RECT 1605.020 5.940 1605.220 6.140 ;
  LAYER VI3 ;
  RECT 1604.620 6.340 1604.820 6.540 ;
  LAYER VI3 ;
  RECT 1604.620 5.940 1604.820 6.140 ;
  LAYER VI3 ;
  RECT 1604.220 6.340 1604.420 6.540 ;
  LAYER VI3 ;
  RECT 1604.220 5.940 1604.420 6.140 ;
  LAYER VI3 ;
  RECT 1603.820 6.340 1604.020 6.540 ;
  LAYER VI3 ;
  RECT 1603.820 5.940 1604.020 6.140 ;
  LAYER VI3 ;
  RECT 1603.420 6.340 1603.620 6.540 ;
  LAYER VI3 ;
  RECT 1603.420 5.940 1603.620 6.140 ;
  LAYER VI3 ;
  RECT 1603.020 6.340 1603.220 6.540 ;
  LAYER VI3 ;
  RECT 1603.020 5.940 1603.220 6.140 ;
  LAYER VI3 ;
  RECT 1602.620 6.340 1602.820 6.540 ;
  LAYER VI3 ;
  RECT 1602.620 5.940 1602.820 6.140 ;
  LAYER VI3 ;
  RECT 1623.700 5.880 1631.700 6.740 ;
  LAYER VI3 ;
  RECT 1631.300 6.340 1631.500 6.540 ;
  LAYER VI3 ;
  RECT 1631.300 5.940 1631.500 6.140 ;
  LAYER VI3 ;
  RECT 1630.900 6.340 1631.100 6.540 ;
  LAYER VI3 ;
  RECT 1630.900 5.940 1631.100 6.140 ;
  LAYER VI3 ;
  RECT 1630.500 6.340 1630.700 6.540 ;
  LAYER VI3 ;
  RECT 1630.500 5.940 1630.700 6.140 ;
  LAYER VI3 ;
  RECT 1630.100 6.340 1630.300 6.540 ;
  LAYER VI3 ;
  RECT 1630.100 5.940 1630.300 6.140 ;
  LAYER VI3 ;
  RECT 1629.700 6.340 1629.900 6.540 ;
  LAYER VI3 ;
  RECT 1629.700 5.940 1629.900 6.140 ;
  LAYER VI3 ;
  RECT 1629.300 6.340 1629.500 6.540 ;
  LAYER VI3 ;
  RECT 1629.300 5.940 1629.500 6.140 ;
  LAYER VI3 ;
  RECT 1628.900 6.340 1629.100 6.540 ;
  LAYER VI3 ;
  RECT 1628.900 5.940 1629.100 6.140 ;
  LAYER VI3 ;
  RECT 1628.500 6.340 1628.700 6.540 ;
  LAYER VI3 ;
  RECT 1628.500 5.940 1628.700 6.140 ;
  LAYER VI3 ;
  RECT 1628.100 6.340 1628.300 6.540 ;
  LAYER VI3 ;
  RECT 1628.100 5.940 1628.300 6.140 ;
  LAYER VI3 ;
  RECT 1627.700 6.340 1627.900 6.540 ;
  LAYER VI3 ;
  RECT 1627.700 5.940 1627.900 6.140 ;
  LAYER VI3 ;
  RECT 1627.300 6.340 1627.500 6.540 ;
  LAYER VI3 ;
  RECT 1627.300 5.940 1627.500 6.140 ;
  LAYER VI3 ;
  RECT 1626.900 6.340 1627.100 6.540 ;
  LAYER VI3 ;
  RECT 1626.900 5.940 1627.100 6.140 ;
  LAYER VI3 ;
  RECT 1626.500 6.340 1626.700 6.540 ;
  LAYER VI3 ;
  RECT 1626.500 5.940 1626.700 6.140 ;
  LAYER VI3 ;
  RECT 1626.100 6.340 1626.300 6.540 ;
  LAYER VI3 ;
  RECT 1626.100 5.940 1626.300 6.140 ;
  LAYER VI3 ;
  RECT 1625.700 6.340 1625.900 6.540 ;
  LAYER VI3 ;
  RECT 1625.700 5.940 1625.900 6.140 ;
  LAYER VI3 ;
  RECT 1625.300 6.340 1625.500 6.540 ;
  LAYER VI3 ;
  RECT 1625.300 5.940 1625.500 6.140 ;
  LAYER VI3 ;
  RECT 1624.900 6.340 1625.100 6.540 ;
  LAYER VI3 ;
  RECT 1624.900 5.940 1625.100 6.140 ;
  LAYER VI3 ;
  RECT 1624.500 6.340 1624.700 6.540 ;
  LAYER VI3 ;
  RECT 1624.500 5.940 1624.700 6.140 ;
  LAYER VI3 ;
  RECT 1624.100 6.340 1624.300 6.540 ;
  LAYER VI3 ;
  RECT 1624.100 5.940 1624.300 6.140 ;
  LAYER VI3 ;
  RECT 1623.700 6.340 1623.900 6.540 ;
  LAYER VI3 ;
  RECT 1623.700 5.940 1623.900 6.140 ;
  LAYER VI3 ;
  RECT 1643.540 5.880 1651.540 6.740 ;
  LAYER VI3 ;
  RECT 1651.140 6.340 1651.340 6.540 ;
  LAYER VI3 ;
  RECT 1651.140 5.940 1651.340 6.140 ;
  LAYER VI3 ;
  RECT 1650.740 6.340 1650.940 6.540 ;
  LAYER VI3 ;
  RECT 1650.740 5.940 1650.940 6.140 ;
  LAYER VI3 ;
  RECT 1650.340 6.340 1650.540 6.540 ;
  LAYER VI3 ;
  RECT 1650.340 5.940 1650.540 6.140 ;
  LAYER VI3 ;
  RECT 1649.940 6.340 1650.140 6.540 ;
  LAYER VI3 ;
  RECT 1649.940 5.940 1650.140 6.140 ;
  LAYER VI3 ;
  RECT 1649.540 6.340 1649.740 6.540 ;
  LAYER VI3 ;
  RECT 1649.540 5.940 1649.740 6.140 ;
  LAYER VI3 ;
  RECT 1649.140 6.340 1649.340 6.540 ;
  LAYER VI3 ;
  RECT 1649.140 5.940 1649.340 6.140 ;
  LAYER VI3 ;
  RECT 1648.740 6.340 1648.940 6.540 ;
  LAYER VI3 ;
  RECT 1648.740 5.940 1648.940 6.140 ;
  LAYER VI3 ;
  RECT 1648.340 6.340 1648.540 6.540 ;
  LAYER VI3 ;
  RECT 1648.340 5.940 1648.540 6.140 ;
  LAYER VI3 ;
  RECT 1647.940 6.340 1648.140 6.540 ;
  LAYER VI3 ;
  RECT 1647.940 5.940 1648.140 6.140 ;
  LAYER VI3 ;
  RECT 1647.540 6.340 1647.740 6.540 ;
  LAYER VI3 ;
  RECT 1647.540 5.940 1647.740 6.140 ;
  LAYER VI3 ;
  RECT 1647.140 6.340 1647.340 6.540 ;
  LAYER VI3 ;
  RECT 1647.140 5.940 1647.340 6.140 ;
  LAYER VI3 ;
  RECT 1646.740 6.340 1646.940 6.540 ;
  LAYER VI3 ;
  RECT 1646.740 5.940 1646.940 6.140 ;
  LAYER VI3 ;
  RECT 1646.340 6.340 1646.540 6.540 ;
  LAYER VI3 ;
  RECT 1646.340 5.940 1646.540 6.140 ;
  LAYER VI3 ;
  RECT 1645.940 6.340 1646.140 6.540 ;
  LAYER VI3 ;
  RECT 1645.940 5.940 1646.140 6.140 ;
  LAYER VI3 ;
  RECT 1645.540 6.340 1645.740 6.540 ;
  LAYER VI3 ;
  RECT 1645.540 5.940 1645.740 6.140 ;
  LAYER VI3 ;
  RECT 1645.140 6.340 1645.340 6.540 ;
  LAYER VI3 ;
  RECT 1645.140 5.940 1645.340 6.140 ;
  LAYER VI3 ;
  RECT 1644.740 6.340 1644.940 6.540 ;
  LAYER VI3 ;
  RECT 1644.740 5.940 1644.940 6.140 ;
  LAYER VI3 ;
  RECT 1644.340 6.340 1644.540 6.540 ;
  LAYER VI3 ;
  RECT 1644.340 5.940 1644.540 6.140 ;
  LAYER VI3 ;
  RECT 1643.940 6.340 1644.140 6.540 ;
  LAYER VI3 ;
  RECT 1643.940 5.940 1644.140 6.140 ;
  LAYER VI3 ;
  RECT 1643.540 6.340 1643.740 6.540 ;
  LAYER VI3 ;
  RECT 1643.540 5.940 1643.740 6.140 ;
  LAYER VI3 ;
  RECT 1664.620 5.880 1672.620 6.740 ;
  LAYER VI3 ;
  RECT 1672.220 6.340 1672.420 6.540 ;
  LAYER VI3 ;
  RECT 1672.220 5.940 1672.420 6.140 ;
  LAYER VI3 ;
  RECT 1671.820 6.340 1672.020 6.540 ;
  LAYER VI3 ;
  RECT 1671.820 5.940 1672.020 6.140 ;
  LAYER VI3 ;
  RECT 1671.420 6.340 1671.620 6.540 ;
  LAYER VI3 ;
  RECT 1671.420 5.940 1671.620 6.140 ;
  LAYER VI3 ;
  RECT 1671.020 6.340 1671.220 6.540 ;
  LAYER VI3 ;
  RECT 1671.020 5.940 1671.220 6.140 ;
  LAYER VI3 ;
  RECT 1670.620 6.340 1670.820 6.540 ;
  LAYER VI3 ;
  RECT 1670.620 5.940 1670.820 6.140 ;
  LAYER VI3 ;
  RECT 1670.220 6.340 1670.420 6.540 ;
  LAYER VI3 ;
  RECT 1670.220 5.940 1670.420 6.140 ;
  LAYER VI3 ;
  RECT 1669.820 6.340 1670.020 6.540 ;
  LAYER VI3 ;
  RECT 1669.820 5.940 1670.020 6.140 ;
  LAYER VI3 ;
  RECT 1669.420 6.340 1669.620 6.540 ;
  LAYER VI3 ;
  RECT 1669.420 5.940 1669.620 6.140 ;
  LAYER VI3 ;
  RECT 1669.020 6.340 1669.220 6.540 ;
  LAYER VI3 ;
  RECT 1669.020 5.940 1669.220 6.140 ;
  LAYER VI3 ;
  RECT 1668.620 6.340 1668.820 6.540 ;
  LAYER VI3 ;
  RECT 1668.620 5.940 1668.820 6.140 ;
  LAYER VI3 ;
  RECT 1668.220 6.340 1668.420 6.540 ;
  LAYER VI3 ;
  RECT 1668.220 5.940 1668.420 6.140 ;
  LAYER VI3 ;
  RECT 1667.820 6.340 1668.020 6.540 ;
  LAYER VI3 ;
  RECT 1667.820 5.940 1668.020 6.140 ;
  LAYER VI3 ;
  RECT 1667.420 6.340 1667.620 6.540 ;
  LAYER VI3 ;
  RECT 1667.420 5.940 1667.620 6.140 ;
  LAYER VI3 ;
  RECT 1667.020 6.340 1667.220 6.540 ;
  LAYER VI3 ;
  RECT 1667.020 5.940 1667.220 6.140 ;
  LAYER VI3 ;
  RECT 1666.620 6.340 1666.820 6.540 ;
  LAYER VI3 ;
  RECT 1666.620 5.940 1666.820 6.140 ;
  LAYER VI3 ;
  RECT 1666.220 6.340 1666.420 6.540 ;
  LAYER VI3 ;
  RECT 1666.220 5.940 1666.420 6.140 ;
  LAYER VI3 ;
  RECT 1665.820 6.340 1666.020 6.540 ;
  LAYER VI3 ;
  RECT 1665.820 5.940 1666.020 6.140 ;
  LAYER VI3 ;
  RECT 1665.420 6.340 1665.620 6.540 ;
  LAYER VI3 ;
  RECT 1665.420 5.940 1665.620 6.140 ;
  LAYER VI3 ;
  RECT 1665.020 6.340 1665.220 6.540 ;
  LAYER VI3 ;
  RECT 1665.020 5.940 1665.220 6.140 ;
  LAYER VI3 ;
  RECT 1664.620 6.340 1664.820 6.540 ;
  LAYER VI3 ;
  RECT 1664.620 5.940 1664.820 6.140 ;
  LAYER VI3 ;
  RECT 1684.460 5.880 1692.460 6.740 ;
  LAYER VI3 ;
  RECT 1692.060 6.340 1692.260 6.540 ;
  LAYER VI3 ;
  RECT 1692.060 5.940 1692.260 6.140 ;
  LAYER VI3 ;
  RECT 1691.660 6.340 1691.860 6.540 ;
  LAYER VI3 ;
  RECT 1691.660 5.940 1691.860 6.140 ;
  LAYER VI3 ;
  RECT 1691.260 6.340 1691.460 6.540 ;
  LAYER VI3 ;
  RECT 1691.260 5.940 1691.460 6.140 ;
  LAYER VI3 ;
  RECT 1690.860 6.340 1691.060 6.540 ;
  LAYER VI3 ;
  RECT 1690.860 5.940 1691.060 6.140 ;
  LAYER VI3 ;
  RECT 1690.460 6.340 1690.660 6.540 ;
  LAYER VI3 ;
  RECT 1690.460 5.940 1690.660 6.140 ;
  LAYER VI3 ;
  RECT 1690.060 6.340 1690.260 6.540 ;
  LAYER VI3 ;
  RECT 1690.060 5.940 1690.260 6.140 ;
  LAYER VI3 ;
  RECT 1689.660 6.340 1689.860 6.540 ;
  LAYER VI3 ;
  RECT 1689.660 5.940 1689.860 6.140 ;
  LAYER VI3 ;
  RECT 1689.260 6.340 1689.460 6.540 ;
  LAYER VI3 ;
  RECT 1689.260 5.940 1689.460 6.140 ;
  LAYER VI3 ;
  RECT 1688.860 6.340 1689.060 6.540 ;
  LAYER VI3 ;
  RECT 1688.860 5.940 1689.060 6.140 ;
  LAYER VI3 ;
  RECT 1688.460 6.340 1688.660 6.540 ;
  LAYER VI3 ;
  RECT 1688.460 5.940 1688.660 6.140 ;
  LAYER VI3 ;
  RECT 1688.060 6.340 1688.260 6.540 ;
  LAYER VI3 ;
  RECT 1688.060 5.940 1688.260 6.140 ;
  LAYER VI3 ;
  RECT 1687.660 6.340 1687.860 6.540 ;
  LAYER VI3 ;
  RECT 1687.660 5.940 1687.860 6.140 ;
  LAYER VI3 ;
  RECT 1687.260 6.340 1687.460 6.540 ;
  LAYER VI3 ;
  RECT 1687.260 5.940 1687.460 6.140 ;
  LAYER VI3 ;
  RECT 1686.860 6.340 1687.060 6.540 ;
  LAYER VI3 ;
  RECT 1686.860 5.940 1687.060 6.140 ;
  LAYER VI3 ;
  RECT 1686.460 6.340 1686.660 6.540 ;
  LAYER VI3 ;
  RECT 1686.460 5.940 1686.660 6.140 ;
  LAYER VI3 ;
  RECT 1686.060 6.340 1686.260 6.540 ;
  LAYER VI3 ;
  RECT 1686.060 5.940 1686.260 6.140 ;
  LAYER VI3 ;
  RECT 1685.660 6.340 1685.860 6.540 ;
  LAYER VI3 ;
  RECT 1685.660 5.940 1685.860 6.140 ;
  LAYER VI3 ;
  RECT 1685.260 6.340 1685.460 6.540 ;
  LAYER VI3 ;
  RECT 1685.260 5.940 1685.460 6.140 ;
  LAYER VI3 ;
  RECT 1684.860 6.340 1685.060 6.540 ;
  LAYER VI3 ;
  RECT 1684.860 5.940 1685.060 6.140 ;
  LAYER VI3 ;
  RECT 1684.460 6.340 1684.660 6.540 ;
  LAYER VI3 ;
  RECT 1684.460 5.940 1684.660 6.140 ;
  LAYER VI3 ;
  RECT 1705.540 5.880 1713.540 6.740 ;
  LAYER VI3 ;
  RECT 1713.140 6.340 1713.340 6.540 ;
  LAYER VI3 ;
  RECT 1713.140 5.940 1713.340 6.140 ;
  LAYER VI3 ;
  RECT 1712.740 6.340 1712.940 6.540 ;
  LAYER VI3 ;
  RECT 1712.740 5.940 1712.940 6.140 ;
  LAYER VI3 ;
  RECT 1712.340 6.340 1712.540 6.540 ;
  LAYER VI3 ;
  RECT 1712.340 5.940 1712.540 6.140 ;
  LAYER VI3 ;
  RECT 1711.940 6.340 1712.140 6.540 ;
  LAYER VI3 ;
  RECT 1711.940 5.940 1712.140 6.140 ;
  LAYER VI3 ;
  RECT 1711.540 6.340 1711.740 6.540 ;
  LAYER VI3 ;
  RECT 1711.540 5.940 1711.740 6.140 ;
  LAYER VI3 ;
  RECT 1711.140 6.340 1711.340 6.540 ;
  LAYER VI3 ;
  RECT 1711.140 5.940 1711.340 6.140 ;
  LAYER VI3 ;
  RECT 1710.740 6.340 1710.940 6.540 ;
  LAYER VI3 ;
  RECT 1710.740 5.940 1710.940 6.140 ;
  LAYER VI3 ;
  RECT 1710.340 6.340 1710.540 6.540 ;
  LAYER VI3 ;
  RECT 1710.340 5.940 1710.540 6.140 ;
  LAYER VI3 ;
  RECT 1709.940 6.340 1710.140 6.540 ;
  LAYER VI3 ;
  RECT 1709.940 5.940 1710.140 6.140 ;
  LAYER VI3 ;
  RECT 1709.540 6.340 1709.740 6.540 ;
  LAYER VI3 ;
  RECT 1709.540 5.940 1709.740 6.140 ;
  LAYER VI3 ;
  RECT 1709.140 6.340 1709.340 6.540 ;
  LAYER VI3 ;
  RECT 1709.140 5.940 1709.340 6.140 ;
  LAYER VI3 ;
  RECT 1708.740 6.340 1708.940 6.540 ;
  LAYER VI3 ;
  RECT 1708.740 5.940 1708.940 6.140 ;
  LAYER VI3 ;
  RECT 1708.340 6.340 1708.540 6.540 ;
  LAYER VI3 ;
  RECT 1708.340 5.940 1708.540 6.140 ;
  LAYER VI3 ;
  RECT 1707.940 6.340 1708.140 6.540 ;
  LAYER VI3 ;
  RECT 1707.940 5.940 1708.140 6.140 ;
  LAYER VI3 ;
  RECT 1707.540 6.340 1707.740 6.540 ;
  LAYER VI3 ;
  RECT 1707.540 5.940 1707.740 6.140 ;
  LAYER VI3 ;
  RECT 1707.140 6.340 1707.340 6.540 ;
  LAYER VI3 ;
  RECT 1707.140 5.940 1707.340 6.140 ;
  LAYER VI3 ;
  RECT 1706.740 6.340 1706.940 6.540 ;
  LAYER VI3 ;
  RECT 1706.740 5.940 1706.940 6.140 ;
  LAYER VI3 ;
  RECT 1706.340 6.340 1706.540 6.540 ;
  LAYER VI3 ;
  RECT 1706.340 5.940 1706.540 6.140 ;
  LAYER VI3 ;
  RECT 1705.940 6.340 1706.140 6.540 ;
  LAYER VI3 ;
  RECT 1705.940 5.940 1706.140 6.140 ;
  LAYER VI3 ;
  RECT 1705.540 6.340 1705.740 6.540 ;
  LAYER VI3 ;
  RECT 1705.540 5.940 1705.740 6.140 ;
  LAYER VI3 ;
  RECT 1725.380 5.880 1733.380 6.740 ;
  LAYER VI3 ;
  RECT 1732.980 6.340 1733.180 6.540 ;
  LAYER VI3 ;
  RECT 1732.980 5.940 1733.180 6.140 ;
  LAYER VI3 ;
  RECT 1732.580 6.340 1732.780 6.540 ;
  LAYER VI3 ;
  RECT 1732.580 5.940 1732.780 6.140 ;
  LAYER VI3 ;
  RECT 1732.180 6.340 1732.380 6.540 ;
  LAYER VI3 ;
  RECT 1732.180 5.940 1732.380 6.140 ;
  LAYER VI3 ;
  RECT 1731.780 6.340 1731.980 6.540 ;
  LAYER VI3 ;
  RECT 1731.780 5.940 1731.980 6.140 ;
  LAYER VI3 ;
  RECT 1731.380 6.340 1731.580 6.540 ;
  LAYER VI3 ;
  RECT 1731.380 5.940 1731.580 6.140 ;
  LAYER VI3 ;
  RECT 1730.980 6.340 1731.180 6.540 ;
  LAYER VI3 ;
  RECT 1730.980 5.940 1731.180 6.140 ;
  LAYER VI3 ;
  RECT 1730.580 6.340 1730.780 6.540 ;
  LAYER VI3 ;
  RECT 1730.580 5.940 1730.780 6.140 ;
  LAYER VI3 ;
  RECT 1730.180 6.340 1730.380 6.540 ;
  LAYER VI3 ;
  RECT 1730.180 5.940 1730.380 6.140 ;
  LAYER VI3 ;
  RECT 1729.780 6.340 1729.980 6.540 ;
  LAYER VI3 ;
  RECT 1729.780 5.940 1729.980 6.140 ;
  LAYER VI3 ;
  RECT 1729.380 6.340 1729.580 6.540 ;
  LAYER VI3 ;
  RECT 1729.380 5.940 1729.580 6.140 ;
  LAYER VI3 ;
  RECT 1728.980 6.340 1729.180 6.540 ;
  LAYER VI3 ;
  RECT 1728.980 5.940 1729.180 6.140 ;
  LAYER VI3 ;
  RECT 1728.580 6.340 1728.780 6.540 ;
  LAYER VI3 ;
  RECT 1728.580 5.940 1728.780 6.140 ;
  LAYER VI3 ;
  RECT 1728.180 6.340 1728.380 6.540 ;
  LAYER VI3 ;
  RECT 1728.180 5.940 1728.380 6.140 ;
  LAYER VI3 ;
  RECT 1727.780 6.340 1727.980 6.540 ;
  LAYER VI3 ;
  RECT 1727.780 5.940 1727.980 6.140 ;
  LAYER VI3 ;
  RECT 1727.380 6.340 1727.580 6.540 ;
  LAYER VI3 ;
  RECT 1727.380 5.940 1727.580 6.140 ;
  LAYER VI3 ;
  RECT 1726.980 6.340 1727.180 6.540 ;
  LAYER VI3 ;
  RECT 1726.980 5.940 1727.180 6.140 ;
  LAYER VI3 ;
  RECT 1726.580 6.340 1726.780 6.540 ;
  LAYER VI3 ;
  RECT 1726.580 5.940 1726.780 6.140 ;
  LAYER VI3 ;
  RECT 1726.180 6.340 1726.380 6.540 ;
  LAYER VI3 ;
  RECT 1726.180 5.940 1726.380 6.140 ;
  LAYER VI3 ;
  RECT 1725.780 6.340 1725.980 6.540 ;
  LAYER VI3 ;
  RECT 1725.780 5.940 1725.980 6.140 ;
  LAYER VI3 ;
  RECT 1725.380 6.340 1725.580 6.540 ;
  LAYER VI3 ;
  RECT 1725.380 5.940 1725.580 6.140 ;
  LAYER VI3 ;
  RECT 1746.460 5.880 1754.460 6.740 ;
  LAYER VI3 ;
  RECT 1754.060 6.340 1754.260 6.540 ;
  LAYER VI3 ;
  RECT 1754.060 5.940 1754.260 6.140 ;
  LAYER VI3 ;
  RECT 1753.660 6.340 1753.860 6.540 ;
  LAYER VI3 ;
  RECT 1753.660 5.940 1753.860 6.140 ;
  LAYER VI3 ;
  RECT 1753.260 6.340 1753.460 6.540 ;
  LAYER VI3 ;
  RECT 1753.260 5.940 1753.460 6.140 ;
  LAYER VI3 ;
  RECT 1752.860 6.340 1753.060 6.540 ;
  LAYER VI3 ;
  RECT 1752.860 5.940 1753.060 6.140 ;
  LAYER VI3 ;
  RECT 1752.460 6.340 1752.660 6.540 ;
  LAYER VI3 ;
  RECT 1752.460 5.940 1752.660 6.140 ;
  LAYER VI3 ;
  RECT 1752.060 6.340 1752.260 6.540 ;
  LAYER VI3 ;
  RECT 1752.060 5.940 1752.260 6.140 ;
  LAYER VI3 ;
  RECT 1751.660 6.340 1751.860 6.540 ;
  LAYER VI3 ;
  RECT 1751.660 5.940 1751.860 6.140 ;
  LAYER VI3 ;
  RECT 1751.260 6.340 1751.460 6.540 ;
  LAYER VI3 ;
  RECT 1751.260 5.940 1751.460 6.140 ;
  LAYER VI3 ;
  RECT 1750.860 6.340 1751.060 6.540 ;
  LAYER VI3 ;
  RECT 1750.860 5.940 1751.060 6.140 ;
  LAYER VI3 ;
  RECT 1750.460 6.340 1750.660 6.540 ;
  LAYER VI3 ;
  RECT 1750.460 5.940 1750.660 6.140 ;
  LAYER VI3 ;
  RECT 1750.060 6.340 1750.260 6.540 ;
  LAYER VI3 ;
  RECT 1750.060 5.940 1750.260 6.140 ;
  LAYER VI3 ;
  RECT 1749.660 6.340 1749.860 6.540 ;
  LAYER VI3 ;
  RECT 1749.660 5.940 1749.860 6.140 ;
  LAYER VI3 ;
  RECT 1749.260 6.340 1749.460 6.540 ;
  LAYER VI3 ;
  RECT 1749.260 5.940 1749.460 6.140 ;
  LAYER VI3 ;
  RECT 1748.860 6.340 1749.060 6.540 ;
  LAYER VI3 ;
  RECT 1748.860 5.940 1749.060 6.140 ;
  LAYER VI3 ;
  RECT 1748.460 6.340 1748.660 6.540 ;
  LAYER VI3 ;
  RECT 1748.460 5.940 1748.660 6.140 ;
  LAYER VI3 ;
  RECT 1748.060 6.340 1748.260 6.540 ;
  LAYER VI3 ;
  RECT 1748.060 5.940 1748.260 6.140 ;
  LAYER VI3 ;
  RECT 1747.660 6.340 1747.860 6.540 ;
  LAYER VI3 ;
  RECT 1747.660 5.940 1747.860 6.140 ;
  LAYER VI3 ;
  RECT 1747.260 6.340 1747.460 6.540 ;
  LAYER VI3 ;
  RECT 1747.260 5.940 1747.460 6.140 ;
  LAYER VI3 ;
  RECT 1746.860 6.340 1747.060 6.540 ;
  LAYER VI3 ;
  RECT 1746.860 5.940 1747.060 6.140 ;
  LAYER VI3 ;
  RECT 1746.460 6.340 1746.660 6.540 ;
  LAYER VI3 ;
  RECT 1746.460 5.940 1746.660 6.140 ;
  LAYER VI3 ;
  RECT 1766.300 5.880 1774.300 6.740 ;
  LAYER VI3 ;
  RECT 1773.900 6.340 1774.100 6.540 ;
  LAYER VI3 ;
  RECT 1773.900 5.940 1774.100 6.140 ;
  LAYER VI3 ;
  RECT 1773.500 6.340 1773.700 6.540 ;
  LAYER VI3 ;
  RECT 1773.500 5.940 1773.700 6.140 ;
  LAYER VI3 ;
  RECT 1773.100 6.340 1773.300 6.540 ;
  LAYER VI3 ;
  RECT 1773.100 5.940 1773.300 6.140 ;
  LAYER VI3 ;
  RECT 1772.700 6.340 1772.900 6.540 ;
  LAYER VI3 ;
  RECT 1772.700 5.940 1772.900 6.140 ;
  LAYER VI3 ;
  RECT 1772.300 6.340 1772.500 6.540 ;
  LAYER VI3 ;
  RECT 1772.300 5.940 1772.500 6.140 ;
  LAYER VI3 ;
  RECT 1771.900 6.340 1772.100 6.540 ;
  LAYER VI3 ;
  RECT 1771.900 5.940 1772.100 6.140 ;
  LAYER VI3 ;
  RECT 1771.500 6.340 1771.700 6.540 ;
  LAYER VI3 ;
  RECT 1771.500 5.940 1771.700 6.140 ;
  LAYER VI3 ;
  RECT 1771.100 6.340 1771.300 6.540 ;
  LAYER VI3 ;
  RECT 1771.100 5.940 1771.300 6.140 ;
  LAYER VI3 ;
  RECT 1770.700 6.340 1770.900 6.540 ;
  LAYER VI3 ;
  RECT 1770.700 5.940 1770.900 6.140 ;
  LAYER VI3 ;
  RECT 1770.300 6.340 1770.500 6.540 ;
  LAYER VI3 ;
  RECT 1770.300 5.940 1770.500 6.140 ;
  LAYER VI3 ;
  RECT 1769.900 6.340 1770.100 6.540 ;
  LAYER VI3 ;
  RECT 1769.900 5.940 1770.100 6.140 ;
  LAYER VI3 ;
  RECT 1769.500 6.340 1769.700 6.540 ;
  LAYER VI3 ;
  RECT 1769.500 5.940 1769.700 6.140 ;
  LAYER VI3 ;
  RECT 1769.100 6.340 1769.300 6.540 ;
  LAYER VI3 ;
  RECT 1769.100 5.940 1769.300 6.140 ;
  LAYER VI3 ;
  RECT 1768.700 6.340 1768.900 6.540 ;
  LAYER VI3 ;
  RECT 1768.700 5.940 1768.900 6.140 ;
  LAYER VI3 ;
  RECT 1768.300 6.340 1768.500 6.540 ;
  LAYER VI3 ;
  RECT 1768.300 5.940 1768.500 6.140 ;
  LAYER VI3 ;
  RECT 1767.900 6.340 1768.100 6.540 ;
  LAYER VI3 ;
  RECT 1767.900 5.940 1768.100 6.140 ;
  LAYER VI3 ;
  RECT 1767.500 6.340 1767.700 6.540 ;
  LAYER VI3 ;
  RECT 1767.500 5.940 1767.700 6.140 ;
  LAYER VI3 ;
  RECT 1767.100 6.340 1767.300 6.540 ;
  LAYER VI3 ;
  RECT 1767.100 5.940 1767.300 6.140 ;
  LAYER VI3 ;
  RECT 1766.700 6.340 1766.900 6.540 ;
  LAYER VI3 ;
  RECT 1766.700 5.940 1766.900 6.140 ;
  LAYER VI3 ;
  RECT 1766.300 6.340 1766.500 6.540 ;
  LAYER VI3 ;
  RECT 1766.300 5.940 1766.500 6.140 ;
  LAYER VI3 ;
  RECT 1787.380 5.880 1795.380 6.740 ;
  LAYER VI3 ;
  RECT 1794.980 6.340 1795.180 6.540 ;
  LAYER VI3 ;
  RECT 1794.980 5.940 1795.180 6.140 ;
  LAYER VI3 ;
  RECT 1794.580 6.340 1794.780 6.540 ;
  LAYER VI3 ;
  RECT 1794.580 5.940 1794.780 6.140 ;
  LAYER VI3 ;
  RECT 1794.180 6.340 1794.380 6.540 ;
  LAYER VI3 ;
  RECT 1794.180 5.940 1794.380 6.140 ;
  LAYER VI3 ;
  RECT 1793.780 6.340 1793.980 6.540 ;
  LAYER VI3 ;
  RECT 1793.780 5.940 1793.980 6.140 ;
  LAYER VI3 ;
  RECT 1793.380 6.340 1793.580 6.540 ;
  LAYER VI3 ;
  RECT 1793.380 5.940 1793.580 6.140 ;
  LAYER VI3 ;
  RECT 1792.980 6.340 1793.180 6.540 ;
  LAYER VI3 ;
  RECT 1792.980 5.940 1793.180 6.140 ;
  LAYER VI3 ;
  RECT 1792.580 6.340 1792.780 6.540 ;
  LAYER VI3 ;
  RECT 1792.580 5.940 1792.780 6.140 ;
  LAYER VI3 ;
  RECT 1792.180 6.340 1792.380 6.540 ;
  LAYER VI3 ;
  RECT 1792.180 5.940 1792.380 6.140 ;
  LAYER VI3 ;
  RECT 1791.780 6.340 1791.980 6.540 ;
  LAYER VI3 ;
  RECT 1791.780 5.940 1791.980 6.140 ;
  LAYER VI3 ;
  RECT 1791.380 6.340 1791.580 6.540 ;
  LAYER VI3 ;
  RECT 1791.380 5.940 1791.580 6.140 ;
  LAYER VI3 ;
  RECT 1790.980 6.340 1791.180 6.540 ;
  LAYER VI3 ;
  RECT 1790.980 5.940 1791.180 6.140 ;
  LAYER VI3 ;
  RECT 1790.580 6.340 1790.780 6.540 ;
  LAYER VI3 ;
  RECT 1790.580 5.940 1790.780 6.140 ;
  LAYER VI3 ;
  RECT 1790.180 6.340 1790.380 6.540 ;
  LAYER VI3 ;
  RECT 1790.180 5.940 1790.380 6.140 ;
  LAYER VI3 ;
  RECT 1789.780 6.340 1789.980 6.540 ;
  LAYER VI3 ;
  RECT 1789.780 5.940 1789.980 6.140 ;
  LAYER VI3 ;
  RECT 1789.380 6.340 1789.580 6.540 ;
  LAYER VI3 ;
  RECT 1789.380 5.940 1789.580 6.140 ;
  LAYER VI3 ;
  RECT 1788.980 6.340 1789.180 6.540 ;
  LAYER VI3 ;
  RECT 1788.980 5.940 1789.180 6.140 ;
  LAYER VI3 ;
  RECT 1788.580 6.340 1788.780 6.540 ;
  LAYER VI3 ;
  RECT 1788.580 5.940 1788.780 6.140 ;
  LAYER VI3 ;
  RECT 1788.180 6.340 1788.380 6.540 ;
  LAYER VI3 ;
  RECT 1788.180 5.940 1788.380 6.140 ;
  LAYER VI3 ;
  RECT 1787.780 6.340 1787.980 6.540 ;
  LAYER VI3 ;
  RECT 1787.780 5.940 1787.980 6.140 ;
  LAYER VI3 ;
  RECT 1787.380 6.340 1787.580 6.540 ;
  LAYER VI3 ;
  RECT 1787.380 5.940 1787.580 6.140 ;
  LAYER VI3 ;
  RECT 1807.220 5.880 1815.220 6.740 ;
  LAYER VI3 ;
  RECT 1814.820 6.340 1815.020 6.540 ;
  LAYER VI3 ;
  RECT 1814.820 5.940 1815.020 6.140 ;
  LAYER VI3 ;
  RECT 1814.420 6.340 1814.620 6.540 ;
  LAYER VI3 ;
  RECT 1814.420 5.940 1814.620 6.140 ;
  LAYER VI3 ;
  RECT 1814.020 6.340 1814.220 6.540 ;
  LAYER VI3 ;
  RECT 1814.020 5.940 1814.220 6.140 ;
  LAYER VI3 ;
  RECT 1813.620 6.340 1813.820 6.540 ;
  LAYER VI3 ;
  RECT 1813.620 5.940 1813.820 6.140 ;
  LAYER VI3 ;
  RECT 1813.220 6.340 1813.420 6.540 ;
  LAYER VI3 ;
  RECT 1813.220 5.940 1813.420 6.140 ;
  LAYER VI3 ;
  RECT 1812.820 6.340 1813.020 6.540 ;
  LAYER VI3 ;
  RECT 1812.820 5.940 1813.020 6.140 ;
  LAYER VI3 ;
  RECT 1812.420 6.340 1812.620 6.540 ;
  LAYER VI3 ;
  RECT 1812.420 5.940 1812.620 6.140 ;
  LAYER VI3 ;
  RECT 1812.020 6.340 1812.220 6.540 ;
  LAYER VI3 ;
  RECT 1812.020 5.940 1812.220 6.140 ;
  LAYER VI3 ;
  RECT 1811.620 6.340 1811.820 6.540 ;
  LAYER VI3 ;
  RECT 1811.620 5.940 1811.820 6.140 ;
  LAYER VI3 ;
  RECT 1811.220 6.340 1811.420 6.540 ;
  LAYER VI3 ;
  RECT 1811.220 5.940 1811.420 6.140 ;
  LAYER VI3 ;
  RECT 1810.820 6.340 1811.020 6.540 ;
  LAYER VI3 ;
  RECT 1810.820 5.940 1811.020 6.140 ;
  LAYER VI3 ;
  RECT 1810.420 6.340 1810.620 6.540 ;
  LAYER VI3 ;
  RECT 1810.420 5.940 1810.620 6.140 ;
  LAYER VI3 ;
  RECT 1810.020 6.340 1810.220 6.540 ;
  LAYER VI3 ;
  RECT 1810.020 5.940 1810.220 6.140 ;
  LAYER VI3 ;
  RECT 1809.620 6.340 1809.820 6.540 ;
  LAYER VI3 ;
  RECT 1809.620 5.940 1809.820 6.140 ;
  LAYER VI3 ;
  RECT 1809.220 6.340 1809.420 6.540 ;
  LAYER VI3 ;
  RECT 1809.220 5.940 1809.420 6.140 ;
  LAYER VI3 ;
  RECT 1808.820 6.340 1809.020 6.540 ;
  LAYER VI3 ;
  RECT 1808.820 5.940 1809.020 6.140 ;
  LAYER VI3 ;
  RECT 1808.420 6.340 1808.620 6.540 ;
  LAYER VI3 ;
  RECT 1808.420 5.940 1808.620 6.140 ;
  LAYER VI3 ;
  RECT 1808.020 6.340 1808.220 6.540 ;
  LAYER VI3 ;
  RECT 1808.020 5.940 1808.220 6.140 ;
  LAYER VI3 ;
  RECT 1807.620 6.340 1807.820 6.540 ;
  LAYER VI3 ;
  RECT 1807.620 5.940 1807.820 6.140 ;
  LAYER VI3 ;
  RECT 1807.220 6.340 1807.420 6.540 ;
  LAYER VI3 ;
  RECT 1807.220 5.940 1807.420 6.140 ;
  LAYER VI3 ;
  RECT 1828.300 5.880 1836.300 6.740 ;
  LAYER VI3 ;
  RECT 1835.900 6.340 1836.100 6.540 ;
  LAYER VI3 ;
  RECT 1835.900 5.940 1836.100 6.140 ;
  LAYER VI3 ;
  RECT 1835.500 6.340 1835.700 6.540 ;
  LAYER VI3 ;
  RECT 1835.500 5.940 1835.700 6.140 ;
  LAYER VI3 ;
  RECT 1835.100 6.340 1835.300 6.540 ;
  LAYER VI3 ;
  RECT 1835.100 5.940 1835.300 6.140 ;
  LAYER VI3 ;
  RECT 1834.700 6.340 1834.900 6.540 ;
  LAYER VI3 ;
  RECT 1834.700 5.940 1834.900 6.140 ;
  LAYER VI3 ;
  RECT 1834.300 6.340 1834.500 6.540 ;
  LAYER VI3 ;
  RECT 1834.300 5.940 1834.500 6.140 ;
  LAYER VI3 ;
  RECT 1833.900 6.340 1834.100 6.540 ;
  LAYER VI3 ;
  RECT 1833.900 5.940 1834.100 6.140 ;
  LAYER VI3 ;
  RECT 1833.500 6.340 1833.700 6.540 ;
  LAYER VI3 ;
  RECT 1833.500 5.940 1833.700 6.140 ;
  LAYER VI3 ;
  RECT 1833.100 6.340 1833.300 6.540 ;
  LAYER VI3 ;
  RECT 1833.100 5.940 1833.300 6.140 ;
  LAYER VI3 ;
  RECT 1832.700 6.340 1832.900 6.540 ;
  LAYER VI3 ;
  RECT 1832.700 5.940 1832.900 6.140 ;
  LAYER VI3 ;
  RECT 1832.300 6.340 1832.500 6.540 ;
  LAYER VI3 ;
  RECT 1832.300 5.940 1832.500 6.140 ;
  LAYER VI3 ;
  RECT 1831.900 6.340 1832.100 6.540 ;
  LAYER VI3 ;
  RECT 1831.900 5.940 1832.100 6.140 ;
  LAYER VI3 ;
  RECT 1831.500 6.340 1831.700 6.540 ;
  LAYER VI3 ;
  RECT 1831.500 5.940 1831.700 6.140 ;
  LAYER VI3 ;
  RECT 1831.100 6.340 1831.300 6.540 ;
  LAYER VI3 ;
  RECT 1831.100 5.940 1831.300 6.140 ;
  LAYER VI3 ;
  RECT 1830.700 6.340 1830.900 6.540 ;
  LAYER VI3 ;
  RECT 1830.700 5.940 1830.900 6.140 ;
  LAYER VI3 ;
  RECT 1830.300 6.340 1830.500 6.540 ;
  LAYER VI3 ;
  RECT 1830.300 5.940 1830.500 6.140 ;
  LAYER VI3 ;
  RECT 1829.900 6.340 1830.100 6.540 ;
  LAYER VI3 ;
  RECT 1829.900 5.940 1830.100 6.140 ;
  LAYER VI3 ;
  RECT 1829.500 6.340 1829.700 6.540 ;
  LAYER VI3 ;
  RECT 1829.500 5.940 1829.700 6.140 ;
  LAYER VI3 ;
  RECT 1829.100 6.340 1829.300 6.540 ;
  LAYER VI3 ;
  RECT 1829.100 5.940 1829.300 6.140 ;
  LAYER VI3 ;
  RECT 1828.700 6.340 1828.900 6.540 ;
  LAYER VI3 ;
  RECT 1828.700 5.940 1828.900 6.140 ;
  LAYER VI3 ;
  RECT 1828.300 6.340 1828.500 6.540 ;
  LAYER VI3 ;
  RECT 1828.300 5.940 1828.500 6.140 ;
  LAYER VI3 ;
  RECT 1848.140 5.880 1856.140 6.740 ;
  LAYER VI3 ;
  RECT 1855.740 6.340 1855.940 6.540 ;
  LAYER VI3 ;
  RECT 1855.740 5.940 1855.940 6.140 ;
  LAYER VI3 ;
  RECT 1855.340 6.340 1855.540 6.540 ;
  LAYER VI3 ;
  RECT 1855.340 5.940 1855.540 6.140 ;
  LAYER VI3 ;
  RECT 1854.940 6.340 1855.140 6.540 ;
  LAYER VI3 ;
  RECT 1854.940 5.940 1855.140 6.140 ;
  LAYER VI3 ;
  RECT 1854.540 6.340 1854.740 6.540 ;
  LAYER VI3 ;
  RECT 1854.540 5.940 1854.740 6.140 ;
  LAYER VI3 ;
  RECT 1854.140 6.340 1854.340 6.540 ;
  LAYER VI3 ;
  RECT 1854.140 5.940 1854.340 6.140 ;
  LAYER VI3 ;
  RECT 1853.740 6.340 1853.940 6.540 ;
  LAYER VI3 ;
  RECT 1853.740 5.940 1853.940 6.140 ;
  LAYER VI3 ;
  RECT 1853.340 6.340 1853.540 6.540 ;
  LAYER VI3 ;
  RECT 1853.340 5.940 1853.540 6.140 ;
  LAYER VI3 ;
  RECT 1852.940 6.340 1853.140 6.540 ;
  LAYER VI3 ;
  RECT 1852.940 5.940 1853.140 6.140 ;
  LAYER VI3 ;
  RECT 1852.540 6.340 1852.740 6.540 ;
  LAYER VI3 ;
  RECT 1852.540 5.940 1852.740 6.140 ;
  LAYER VI3 ;
  RECT 1852.140 6.340 1852.340 6.540 ;
  LAYER VI3 ;
  RECT 1852.140 5.940 1852.340 6.140 ;
  LAYER VI3 ;
  RECT 1851.740 6.340 1851.940 6.540 ;
  LAYER VI3 ;
  RECT 1851.740 5.940 1851.940 6.140 ;
  LAYER VI3 ;
  RECT 1851.340 6.340 1851.540 6.540 ;
  LAYER VI3 ;
  RECT 1851.340 5.940 1851.540 6.140 ;
  LAYER VI3 ;
  RECT 1850.940 6.340 1851.140 6.540 ;
  LAYER VI3 ;
  RECT 1850.940 5.940 1851.140 6.140 ;
  LAYER VI3 ;
  RECT 1850.540 6.340 1850.740 6.540 ;
  LAYER VI3 ;
  RECT 1850.540 5.940 1850.740 6.140 ;
  LAYER VI3 ;
  RECT 1850.140 6.340 1850.340 6.540 ;
  LAYER VI3 ;
  RECT 1850.140 5.940 1850.340 6.140 ;
  LAYER VI3 ;
  RECT 1849.740 6.340 1849.940 6.540 ;
  LAYER VI3 ;
  RECT 1849.740 5.940 1849.940 6.140 ;
  LAYER VI3 ;
  RECT 1849.340 6.340 1849.540 6.540 ;
  LAYER VI3 ;
  RECT 1849.340 5.940 1849.540 6.140 ;
  LAYER VI3 ;
  RECT 1848.940 6.340 1849.140 6.540 ;
  LAYER VI3 ;
  RECT 1848.940 5.940 1849.140 6.140 ;
  LAYER VI3 ;
  RECT 1848.540 6.340 1848.740 6.540 ;
  LAYER VI3 ;
  RECT 1848.540 5.940 1848.740 6.140 ;
  LAYER VI3 ;
  RECT 1848.140 6.340 1848.340 6.540 ;
  LAYER VI3 ;
  RECT 1848.140 5.940 1848.340 6.140 ;
  LAYER VI3 ;
  RECT 1869.220 5.880 1877.220 6.740 ;
  LAYER VI3 ;
  RECT 1876.820 6.340 1877.020 6.540 ;
  LAYER VI3 ;
  RECT 1876.820 5.940 1877.020 6.140 ;
  LAYER VI3 ;
  RECT 1876.420 6.340 1876.620 6.540 ;
  LAYER VI3 ;
  RECT 1876.420 5.940 1876.620 6.140 ;
  LAYER VI3 ;
  RECT 1876.020 6.340 1876.220 6.540 ;
  LAYER VI3 ;
  RECT 1876.020 5.940 1876.220 6.140 ;
  LAYER VI3 ;
  RECT 1875.620 6.340 1875.820 6.540 ;
  LAYER VI3 ;
  RECT 1875.620 5.940 1875.820 6.140 ;
  LAYER VI3 ;
  RECT 1875.220 6.340 1875.420 6.540 ;
  LAYER VI3 ;
  RECT 1875.220 5.940 1875.420 6.140 ;
  LAYER VI3 ;
  RECT 1874.820 6.340 1875.020 6.540 ;
  LAYER VI3 ;
  RECT 1874.820 5.940 1875.020 6.140 ;
  LAYER VI3 ;
  RECT 1874.420 6.340 1874.620 6.540 ;
  LAYER VI3 ;
  RECT 1874.420 5.940 1874.620 6.140 ;
  LAYER VI3 ;
  RECT 1874.020 6.340 1874.220 6.540 ;
  LAYER VI3 ;
  RECT 1874.020 5.940 1874.220 6.140 ;
  LAYER VI3 ;
  RECT 1873.620 6.340 1873.820 6.540 ;
  LAYER VI3 ;
  RECT 1873.620 5.940 1873.820 6.140 ;
  LAYER VI3 ;
  RECT 1873.220 6.340 1873.420 6.540 ;
  LAYER VI3 ;
  RECT 1873.220 5.940 1873.420 6.140 ;
  LAYER VI3 ;
  RECT 1872.820 6.340 1873.020 6.540 ;
  LAYER VI3 ;
  RECT 1872.820 5.940 1873.020 6.140 ;
  LAYER VI3 ;
  RECT 1872.420 6.340 1872.620 6.540 ;
  LAYER VI3 ;
  RECT 1872.420 5.940 1872.620 6.140 ;
  LAYER VI3 ;
  RECT 1872.020 6.340 1872.220 6.540 ;
  LAYER VI3 ;
  RECT 1872.020 5.940 1872.220 6.140 ;
  LAYER VI3 ;
  RECT 1871.620 6.340 1871.820 6.540 ;
  LAYER VI3 ;
  RECT 1871.620 5.940 1871.820 6.140 ;
  LAYER VI3 ;
  RECT 1871.220 6.340 1871.420 6.540 ;
  LAYER VI3 ;
  RECT 1871.220 5.940 1871.420 6.140 ;
  LAYER VI3 ;
  RECT 1870.820 6.340 1871.020 6.540 ;
  LAYER VI3 ;
  RECT 1870.820 5.940 1871.020 6.140 ;
  LAYER VI3 ;
  RECT 1870.420 6.340 1870.620 6.540 ;
  LAYER VI3 ;
  RECT 1870.420 5.940 1870.620 6.140 ;
  LAYER VI3 ;
  RECT 1870.020 6.340 1870.220 6.540 ;
  LAYER VI3 ;
  RECT 1870.020 5.940 1870.220 6.140 ;
  LAYER VI3 ;
  RECT 1869.620 6.340 1869.820 6.540 ;
  LAYER VI3 ;
  RECT 1869.620 5.940 1869.820 6.140 ;
  LAYER VI3 ;
  RECT 1869.220 6.340 1869.420 6.540 ;
  LAYER VI3 ;
  RECT 1869.220 5.940 1869.420 6.140 ;
  LAYER VI3 ;
  RECT 1889.060 5.880 1897.060 6.740 ;
  LAYER VI3 ;
  RECT 1896.660 6.340 1896.860 6.540 ;
  LAYER VI3 ;
  RECT 1896.660 5.940 1896.860 6.140 ;
  LAYER VI3 ;
  RECT 1896.260 6.340 1896.460 6.540 ;
  LAYER VI3 ;
  RECT 1896.260 5.940 1896.460 6.140 ;
  LAYER VI3 ;
  RECT 1895.860 6.340 1896.060 6.540 ;
  LAYER VI3 ;
  RECT 1895.860 5.940 1896.060 6.140 ;
  LAYER VI3 ;
  RECT 1895.460 6.340 1895.660 6.540 ;
  LAYER VI3 ;
  RECT 1895.460 5.940 1895.660 6.140 ;
  LAYER VI3 ;
  RECT 1895.060 6.340 1895.260 6.540 ;
  LAYER VI3 ;
  RECT 1895.060 5.940 1895.260 6.140 ;
  LAYER VI3 ;
  RECT 1894.660 6.340 1894.860 6.540 ;
  LAYER VI3 ;
  RECT 1894.660 5.940 1894.860 6.140 ;
  LAYER VI3 ;
  RECT 1894.260 6.340 1894.460 6.540 ;
  LAYER VI3 ;
  RECT 1894.260 5.940 1894.460 6.140 ;
  LAYER VI3 ;
  RECT 1893.860 6.340 1894.060 6.540 ;
  LAYER VI3 ;
  RECT 1893.860 5.940 1894.060 6.140 ;
  LAYER VI3 ;
  RECT 1893.460 6.340 1893.660 6.540 ;
  LAYER VI3 ;
  RECT 1893.460 5.940 1893.660 6.140 ;
  LAYER VI3 ;
  RECT 1893.060 6.340 1893.260 6.540 ;
  LAYER VI3 ;
  RECT 1893.060 5.940 1893.260 6.140 ;
  LAYER VI3 ;
  RECT 1892.660 6.340 1892.860 6.540 ;
  LAYER VI3 ;
  RECT 1892.660 5.940 1892.860 6.140 ;
  LAYER VI3 ;
  RECT 1892.260 6.340 1892.460 6.540 ;
  LAYER VI3 ;
  RECT 1892.260 5.940 1892.460 6.140 ;
  LAYER VI3 ;
  RECT 1891.860 6.340 1892.060 6.540 ;
  LAYER VI3 ;
  RECT 1891.860 5.940 1892.060 6.140 ;
  LAYER VI3 ;
  RECT 1891.460 6.340 1891.660 6.540 ;
  LAYER VI3 ;
  RECT 1891.460 5.940 1891.660 6.140 ;
  LAYER VI3 ;
  RECT 1891.060 6.340 1891.260 6.540 ;
  LAYER VI3 ;
  RECT 1891.060 5.940 1891.260 6.140 ;
  LAYER VI3 ;
  RECT 1890.660 6.340 1890.860 6.540 ;
  LAYER VI3 ;
  RECT 1890.660 5.940 1890.860 6.140 ;
  LAYER VI3 ;
  RECT 1890.260 6.340 1890.460 6.540 ;
  LAYER VI3 ;
  RECT 1890.260 5.940 1890.460 6.140 ;
  LAYER VI3 ;
  RECT 1889.860 6.340 1890.060 6.540 ;
  LAYER VI3 ;
  RECT 1889.860 5.940 1890.060 6.140 ;
  LAYER VI3 ;
  RECT 1889.460 6.340 1889.660 6.540 ;
  LAYER VI3 ;
  RECT 1889.460 5.940 1889.660 6.140 ;
  LAYER VI3 ;
  RECT 1889.060 6.340 1889.260 6.540 ;
  LAYER VI3 ;
  RECT 1889.060 5.940 1889.260 6.140 ;
  LAYER VI3 ;
  RECT 1910.140 5.880 1918.140 6.740 ;
  LAYER VI3 ;
  RECT 1917.740 6.340 1917.940 6.540 ;
  LAYER VI3 ;
  RECT 1917.740 5.940 1917.940 6.140 ;
  LAYER VI3 ;
  RECT 1917.340 6.340 1917.540 6.540 ;
  LAYER VI3 ;
  RECT 1917.340 5.940 1917.540 6.140 ;
  LAYER VI3 ;
  RECT 1916.940 6.340 1917.140 6.540 ;
  LAYER VI3 ;
  RECT 1916.940 5.940 1917.140 6.140 ;
  LAYER VI3 ;
  RECT 1916.540 6.340 1916.740 6.540 ;
  LAYER VI3 ;
  RECT 1916.540 5.940 1916.740 6.140 ;
  LAYER VI3 ;
  RECT 1916.140 6.340 1916.340 6.540 ;
  LAYER VI3 ;
  RECT 1916.140 5.940 1916.340 6.140 ;
  LAYER VI3 ;
  RECT 1915.740 6.340 1915.940 6.540 ;
  LAYER VI3 ;
  RECT 1915.740 5.940 1915.940 6.140 ;
  LAYER VI3 ;
  RECT 1915.340 6.340 1915.540 6.540 ;
  LAYER VI3 ;
  RECT 1915.340 5.940 1915.540 6.140 ;
  LAYER VI3 ;
  RECT 1914.940 6.340 1915.140 6.540 ;
  LAYER VI3 ;
  RECT 1914.940 5.940 1915.140 6.140 ;
  LAYER VI3 ;
  RECT 1914.540 6.340 1914.740 6.540 ;
  LAYER VI3 ;
  RECT 1914.540 5.940 1914.740 6.140 ;
  LAYER VI3 ;
  RECT 1914.140 6.340 1914.340 6.540 ;
  LAYER VI3 ;
  RECT 1914.140 5.940 1914.340 6.140 ;
  LAYER VI3 ;
  RECT 1913.740 6.340 1913.940 6.540 ;
  LAYER VI3 ;
  RECT 1913.740 5.940 1913.940 6.140 ;
  LAYER VI3 ;
  RECT 1913.340 6.340 1913.540 6.540 ;
  LAYER VI3 ;
  RECT 1913.340 5.940 1913.540 6.140 ;
  LAYER VI3 ;
  RECT 1912.940 6.340 1913.140 6.540 ;
  LAYER VI3 ;
  RECT 1912.940 5.940 1913.140 6.140 ;
  LAYER VI3 ;
  RECT 1912.540 6.340 1912.740 6.540 ;
  LAYER VI3 ;
  RECT 1912.540 5.940 1912.740 6.140 ;
  LAYER VI3 ;
  RECT 1912.140 6.340 1912.340 6.540 ;
  LAYER VI3 ;
  RECT 1912.140 5.940 1912.340 6.140 ;
  LAYER VI3 ;
  RECT 1911.740 6.340 1911.940 6.540 ;
  LAYER VI3 ;
  RECT 1911.740 5.940 1911.940 6.140 ;
  LAYER VI3 ;
  RECT 1911.340 6.340 1911.540 6.540 ;
  LAYER VI3 ;
  RECT 1911.340 5.940 1911.540 6.140 ;
  LAYER VI3 ;
  RECT 1910.940 6.340 1911.140 6.540 ;
  LAYER VI3 ;
  RECT 1910.940 5.940 1911.140 6.140 ;
  LAYER VI3 ;
  RECT 1910.540 6.340 1910.740 6.540 ;
  LAYER VI3 ;
  RECT 1910.540 5.940 1910.740 6.140 ;
  LAYER VI3 ;
  RECT 1910.140 6.340 1910.340 6.540 ;
  LAYER VI3 ;
  RECT 1910.140 5.940 1910.340 6.140 ;
  LAYER VI3 ;
  RECT 1929.980 5.880 1937.980 6.740 ;
  LAYER VI3 ;
  RECT 1937.580 6.340 1937.780 6.540 ;
  LAYER VI3 ;
  RECT 1937.580 5.940 1937.780 6.140 ;
  LAYER VI3 ;
  RECT 1937.180 6.340 1937.380 6.540 ;
  LAYER VI3 ;
  RECT 1937.180 5.940 1937.380 6.140 ;
  LAYER VI3 ;
  RECT 1936.780 6.340 1936.980 6.540 ;
  LAYER VI3 ;
  RECT 1936.780 5.940 1936.980 6.140 ;
  LAYER VI3 ;
  RECT 1936.380 6.340 1936.580 6.540 ;
  LAYER VI3 ;
  RECT 1936.380 5.940 1936.580 6.140 ;
  LAYER VI3 ;
  RECT 1935.980 6.340 1936.180 6.540 ;
  LAYER VI3 ;
  RECT 1935.980 5.940 1936.180 6.140 ;
  LAYER VI3 ;
  RECT 1935.580 6.340 1935.780 6.540 ;
  LAYER VI3 ;
  RECT 1935.580 5.940 1935.780 6.140 ;
  LAYER VI3 ;
  RECT 1935.180 6.340 1935.380 6.540 ;
  LAYER VI3 ;
  RECT 1935.180 5.940 1935.380 6.140 ;
  LAYER VI3 ;
  RECT 1934.780 6.340 1934.980 6.540 ;
  LAYER VI3 ;
  RECT 1934.780 5.940 1934.980 6.140 ;
  LAYER VI3 ;
  RECT 1934.380 6.340 1934.580 6.540 ;
  LAYER VI3 ;
  RECT 1934.380 5.940 1934.580 6.140 ;
  LAYER VI3 ;
  RECT 1933.980 6.340 1934.180 6.540 ;
  LAYER VI3 ;
  RECT 1933.980 5.940 1934.180 6.140 ;
  LAYER VI3 ;
  RECT 1933.580 6.340 1933.780 6.540 ;
  LAYER VI3 ;
  RECT 1933.580 5.940 1933.780 6.140 ;
  LAYER VI3 ;
  RECT 1933.180 6.340 1933.380 6.540 ;
  LAYER VI3 ;
  RECT 1933.180 5.940 1933.380 6.140 ;
  LAYER VI3 ;
  RECT 1932.780 6.340 1932.980 6.540 ;
  LAYER VI3 ;
  RECT 1932.780 5.940 1932.980 6.140 ;
  LAYER VI3 ;
  RECT 1932.380 6.340 1932.580 6.540 ;
  LAYER VI3 ;
  RECT 1932.380 5.940 1932.580 6.140 ;
  LAYER VI3 ;
  RECT 1931.980 6.340 1932.180 6.540 ;
  LAYER VI3 ;
  RECT 1931.980 5.940 1932.180 6.140 ;
  LAYER VI3 ;
  RECT 1931.580 6.340 1931.780 6.540 ;
  LAYER VI3 ;
  RECT 1931.580 5.940 1931.780 6.140 ;
  LAYER VI3 ;
  RECT 1931.180 6.340 1931.380 6.540 ;
  LAYER VI3 ;
  RECT 1931.180 5.940 1931.380 6.140 ;
  LAYER VI3 ;
  RECT 1930.780 6.340 1930.980 6.540 ;
  LAYER VI3 ;
  RECT 1930.780 5.940 1930.980 6.140 ;
  LAYER VI3 ;
  RECT 1930.380 6.340 1930.580 6.540 ;
  LAYER VI3 ;
  RECT 1930.380 5.940 1930.580 6.140 ;
  LAYER VI3 ;
  RECT 1929.980 6.340 1930.180 6.540 ;
  LAYER VI3 ;
  RECT 1929.980 5.940 1930.180 6.140 ;
  LAYER VI3 ;
  RECT 1951.060 5.880 1959.060 6.740 ;
  LAYER VI3 ;
  RECT 1958.660 6.340 1958.860 6.540 ;
  LAYER VI3 ;
  RECT 1958.660 5.940 1958.860 6.140 ;
  LAYER VI3 ;
  RECT 1958.260 6.340 1958.460 6.540 ;
  LAYER VI3 ;
  RECT 1958.260 5.940 1958.460 6.140 ;
  LAYER VI3 ;
  RECT 1957.860 6.340 1958.060 6.540 ;
  LAYER VI3 ;
  RECT 1957.860 5.940 1958.060 6.140 ;
  LAYER VI3 ;
  RECT 1957.460 6.340 1957.660 6.540 ;
  LAYER VI3 ;
  RECT 1957.460 5.940 1957.660 6.140 ;
  LAYER VI3 ;
  RECT 1957.060 6.340 1957.260 6.540 ;
  LAYER VI3 ;
  RECT 1957.060 5.940 1957.260 6.140 ;
  LAYER VI3 ;
  RECT 1956.660 6.340 1956.860 6.540 ;
  LAYER VI3 ;
  RECT 1956.660 5.940 1956.860 6.140 ;
  LAYER VI3 ;
  RECT 1956.260 6.340 1956.460 6.540 ;
  LAYER VI3 ;
  RECT 1956.260 5.940 1956.460 6.140 ;
  LAYER VI3 ;
  RECT 1955.860 6.340 1956.060 6.540 ;
  LAYER VI3 ;
  RECT 1955.860 5.940 1956.060 6.140 ;
  LAYER VI3 ;
  RECT 1955.460 6.340 1955.660 6.540 ;
  LAYER VI3 ;
  RECT 1955.460 5.940 1955.660 6.140 ;
  LAYER VI3 ;
  RECT 1955.060 6.340 1955.260 6.540 ;
  LAYER VI3 ;
  RECT 1955.060 5.940 1955.260 6.140 ;
  LAYER VI3 ;
  RECT 1954.660 6.340 1954.860 6.540 ;
  LAYER VI3 ;
  RECT 1954.660 5.940 1954.860 6.140 ;
  LAYER VI3 ;
  RECT 1954.260 6.340 1954.460 6.540 ;
  LAYER VI3 ;
  RECT 1954.260 5.940 1954.460 6.140 ;
  LAYER VI3 ;
  RECT 1953.860 6.340 1954.060 6.540 ;
  LAYER VI3 ;
  RECT 1953.860 5.940 1954.060 6.140 ;
  LAYER VI3 ;
  RECT 1953.460 6.340 1953.660 6.540 ;
  LAYER VI3 ;
  RECT 1953.460 5.940 1953.660 6.140 ;
  LAYER VI3 ;
  RECT 1953.060 6.340 1953.260 6.540 ;
  LAYER VI3 ;
  RECT 1953.060 5.940 1953.260 6.140 ;
  LAYER VI3 ;
  RECT 1952.660 6.340 1952.860 6.540 ;
  LAYER VI3 ;
  RECT 1952.660 5.940 1952.860 6.140 ;
  LAYER VI3 ;
  RECT 1952.260 6.340 1952.460 6.540 ;
  LAYER VI3 ;
  RECT 1952.260 5.940 1952.460 6.140 ;
  LAYER VI3 ;
  RECT 1951.860 6.340 1952.060 6.540 ;
  LAYER VI3 ;
  RECT 1951.860 5.940 1952.060 6.140 ;
  LAYER VI3 ;
  RECT 1951.460 6.340 1951.660 6.540 ;
  LAYER VI3 ;
  RECT 1951.460 5.940 1951.660 6.140 ;
  LAYER VI3 ;
  RECT 1951.060 6.340 1951.260 6.540 ;
  LAYER VI3 ;
  RECT 1951.060 5.940 1951.260 6.140 ;
  LAYER VI3 ;
  RECT 1970.900 5.880 1978.900 6.740 ;
  LAYER VI3 ;
  RECT 1978.500 6.340 1978.700 6.540 ;
  LAYER VI3 ;
  RECT 1978.500 5.940 1978.700 6.140 ;
  LAYER VI3 ;
  RECT 1978.100 6.340 1978.300 6.540 ;
  LAYER VI3 ;
  RECT 1978.100 5.940 1978.300 6.140 ;
  LAYER VI3 ;
  RECT 1977.700 6.340 1977.900 6.540 ;
  LAYER VI3 ;
  RECT 1977.700 5.940 1977.900 6.140 ;
  LAYER VI3 ;
  RECT 1977.300 6.340 1977.500 6.540 ;
  LAYER VI3 ;
  RECT 1977.300 5.940 1977.500 6.140 ;
  LAYER VI3 ;
  RECT 1976.900 6.340 1977.100 6.540 ;
  LAYER VI3 ;
  RECT 1976.900 5.940 1977.100 6.140 ;
  LAYER VI3 ;
  RECT 1976.500 6.340 1976.700 6.540 ;
  LAYER VI3 ;
  RECT 1976.500 5.940 1976.700 6.140 ;
  LAYER VI3 ;
  RECT 1976.100 6.340 1976.300 6.540 ;
  LAYER VI3 ;
  RECT 1976.100 5.940 1976.300 6.140 ;
  LAYER VI3 ;
  RECT 1975.700 6.340 1975.900 6.540 ;
  LAYER VI3 ;
  RECT 1975.700 5.940 1975.900 6.140 ;
  LAYER VI3 ;
  RECT 1975.300 6.340 1975.500 6.540 ;
  LAYER VI3 ;
  RECT 1975.300 5.940 1975.500 6.140 ;
  LAYER VI3 ;
  RECT 1974.900 6.340 1975.100 6.540 ;
  LAYER VI3 ;
  RECT 1974.900 5.940 1975.100 6.140 ;
  LAYER VI3 ;
  RECT 1974.500 6.340 1974.700 6.540 ;
  LAYER VI3 ;
  RECT 1974.500 5.940 1974.700 6.140 ;
  LAYER VI3 ;
  RECT 1974.100 6.340 1974.300 6.540 ;
  LAYER VI3 ;
  RECT 1974.100 5.940 1974.300 6.140 ;
  LAYER VI3 ;
  RECT 1973.700 6.340 1973.900 6.540 ;
  LAYER VI3 ;
  RECT 1973.700 5.940 1973.900 6.140 ;
  LAYER VI3 ;
  RECT 1973.300 6.340 1973.500 6.540 ;
  LAYER VI3 ;
  RECT 1973.300 5.940 1973.500 6.140 ;
  LAYER VI3 ;
  RECT 1972.900 6.340 1973.100 6.540 ;
  LAYER VI3 ;
  RECT 1972.900 5.940 1973.100 6.140 ;
  LAYER VI3 ;
  RECT 1972.500 6.340 1972.700 6.540 ;
  LAYER VI3 ;
  RECT 1972.500 5.940 1972.700 6.140 ;
  LAYER VI3 ;
  RECT 1972.100 6.340 1972.300 6.540 ;
  LAYER VI3 ;
  RECT 1972.100 5.940 1972.300 6.140 ;
  LAYER VI3 ;
  RECT 1971.700 6.340 1971.900 6.540 ;
  LAYER VI3 ;
  RECT 1971.700 5.940 1971.900 6.140 ;
  LAYER VI3 ;
  RECT 1971.300 6.340 1971.500 6.540 ;
  LAYER VI3 ;
  RECT 1971.300 5.940 1971.500 6.140 ;
  LAYER VI3 ;
  RECT 1970.900 6.340 1971.100 6.540 ;
  LAYER VI3 ;
  RECT 1970.900 5.940 1971.100 6.140 ;
  LAYER VI3 ;
  RECT 1991.980 5.880 1999.980 6.740 ;
  LAYER VI3 ;
  RECT 1999.580 6.340 1999.780 6.540 ;
  LAYER VI3 ;
  RECT 1999.580 5.940 1999.780 6.140 ;
  LAYER VI3 ;
  RECT 1999.180 6.340 1999.380 6.540 ;
  LAYER VI3 ;
  RECT 1999.180 5.940 1999.380 6.140 ;
  LAYER VI3 ;
  RECT 1998.780 6.340 1998.980 6.540 ;
  LAYER VI3 ;
  RECT 1998.780 5.940 1998.980 6.140 ;
  LAYER VI3 ;
  RECT 1998.380 6.340 1998.580 6.540 ;
  LAYER VI3 ;
  RECT 1998.380 5.940 1998.580 6.140 ;
  LAYER VI3 ;
  RECT 1997.980 6.340 1998.180 6.540 ;
  LAYER VI3 ;
  RECT 1997.980 5.940 1998.180 6.140 ;
  LAYER VI3 ;
  RECT 1997.580 6.340 1997.780 6.540 ;
  LAYER VI3 ;
  RECT 1997.580 5.940 1997.780 6.140 ;
  LAYER VI3 ;
  RECT 1997.180 6.340 1997.380 6.540 ;
  LAYER VI3 ;
  RECT 1997.180 5.940 1997.380 6.140 ;
  LAYER VI3 ;
  RECT 1996.780 6.340 1996.980 6.540 ;
  LAYER VI3 ;
  RECT 1996.780 5.940 1996.980 6.140 ;
  LAYER VI3 ;
  RECT 1996.380 6.340 1996.580 6.540 ;
  LAYER VI3 ;
  RECT 1996.380 5.940 1996.580 6.140 ;
  LAYER VI3 ;
  RECT 1995.980 6.340 1996.180 6.540 ;
  LAYER VI3 ;
  RECT 1995.980 5.940 1996.180 6.140 ;
  LAYER VI3 ;
  RECT 1995.580 6.340 1995.780 6.540 ;
  LAYER VI3 ;
  RECT 1995.580 5.940 1995.780 6.140 ;
  LAYER VI3 ;
  RECT 1995.180 6.340 1995.380 6.540 ;
  LAYER VI3 ;
  RECT 1995.180 5.940 1995.380 6.140 ;
  LAYER VI3 ;
  RECT 1994.780 6.340 1994.980 6.540 ;
  LAYER VI3 ;
  RECT 1994.780 5.940 1994.980 6.140 ;
  LAYER VI3 ;
  RECT 1994.380 6.340 1994.580 6.540 ;
  LAYER VI3 ;
  RECT 1994.380 5.940 1994.580 6.140 ;
  LAYER VI3 ;
  RECT 1993.980 6.340 1994.180 6.540 ;
  LAYER VI3 ;
  RECT 1993.980 5.940 1994.180 6.140 ;
  LAYER VI3 ;
  RECT 1993.580 6.340 1993.780 6.540 ;
  LAYER VI3 ;
  RECT 1993.580 5.940 1993.780 6.140 ;
  LAYER VI3 ;
  RECT 1993.180 6.340 1993.380 6.540 ;
  LAYER VI3 ;
  RECT 1993.180 5.940 1993.380 6.140 ;
  LAYER VI3 ;
  RECT 1992.780 6.340 1992.980 6.540 ;
  LAYER VI3 ;
  RECT 1992.780 5.940 1992.980 6.140 ;
  LAYER VI3 ;
  RECT 1992.380 6.340 1992.580 6.540 ;
  LAYER VI3 ;
  RECT 1992.380 5.940 1992.580 6.140 ;
  LAYER VI3 ;
  RECT 1991.980 6.340 1992.180 6.540 ;
  LAYER VI3 ;
  RECT 1991.980 5.940 1992.180 6.140 ;
  LAYER VI3 ;
  RECT 2011.820 5.880 2019.820 6.740 ;
  LAYER VI3 ;
  RECT 2019.420 6.340 2019.620 6.540 ;
  LAYER VI3 ;
  RECT 2019.420 5.940 2019.620 6.140 ;
  LAYER VI3 ;
  RECT 2019.020 6.340 2019.220 6.540 ;
  LAYER VI3 ;
  RECT 2019.020 5.940 2019.220 6.140 ;
  LAYER VI3 ;
  RECT 2018.620 6.340 2018.820 6.540 ;
  LAYER VI3 ;
  RECT 2018.620 5.940 2018.820 6.140 ;
  LAYER VI3 ;
  RECT 2018.220 6.340 2018.420 6.540 ;
  LAYER VI3 ;
  RECT 2018.220 5.940 2018.420 6.140 ;
  LAYER VI3 ;
  RECT 2017.820 6.340 2018.020 6.540 ;
  LAYER VI3 ;
  RECT 2017.820 5.940 2018.020 6.140 ;
  LAYER VI3 ;
  RECT 2017.420 6.340 2017.620 6.540 ;
  LAYER VI3 ;
  RECT 2017.420 5.940 2017.620 6.140 ;
  LAYER VI3 ;
  RECT 2017.020 6.340 2017.220 6.540 ;
  LAYER VI3 ;
  RECT 2017.020 5.940 2017.220 6.140 ;
  LAYER VI3 ;
  RECT 2016.620 6.340 2016.820 6.540 ;
  LAYER VI3 ;
  RECT 2016.620 5.940 2016.820 6.140 ;
  LAYER VI3 ;
  RECT 2016.220 6.340 2016.420 6.540 ;
  LAYER VI3 ;
  RECT 2016.220 5.940 2016.420 6.140 ;
  LAYER VI3 ;
  RECT 2015.820 6.340 2016.020 6.540 ;
  LAYER VI3 ;
  RECT 2015.820 5.940 2016.020 6.140 ;
  LAYER VI3 ;
  RECT 2015.420 6.340 2015.620 6.540 ;
  LAYER VI3 ;
  RECT 2015.420 5.940 2015.620 6.140 ;
  LAYER VI3 ;
  RECT 2015.020 6.340 2015.220 6.540 ;
  LAYER VI3 ;
  RECT 2015.020 5.940 2015.220 6.140 ;
  LAYER VI3 ;
  RECT 2014.620 6.340 2014.820 6.540 ;
  LAYER VI3 ;
  RECT 2014.620 5.940 2014.820 6.140 ;
  LAYER VI3 ;
  RECT 2014.220 6.340 2014.420 6.540 ;
  LAYER VI3 ;
  RECT 2014.220 5.940 2014.420 6.140 ;
  LAYER VI3 ;
  RECT 2013.820 6.340 2014.020 6.540 ;
  LAYER VI3 ;
  RECT 2013.820 5.940 2014.020 6.140 ;
  LAYER VI3 ;
  RECT 2013.420 6.340 2013.620 6.540 ;
  LAYER VI3 ;
  RECT 2013.420 5.940 2013.620 6.140 ;
  LAYER VI3 ;
  RECT 2013.020 6.340 2013.220 6.540 ;
  LAYER VI3 ;
  RECT 2013.020 5.940 2013.220 6.140 ;
  LAYER VI3 ;
  RECT 2012.620 6.340 2012.820 6.540 ;
  LAYER VI3 ;
  RECT 2012.620 5.940 2012.820 6.140 ;
  LAYER VI3 ;
  RECT 2012.220 6.340 2012.420 6.540 ;
  LAYER VI3 ;
  RECT 2012.220 5.940 2012.420 6.140 ;
  LAYER VI3 ;
  RECT 2011.820 6.340 2012.020 6.540 ;
  LAYER VI3 ;
  RECT 2011.820 5.940 2012.020 6.140 ;
  LAYER VI3 ;
  RECT 2032.900 5.880 2040.900 6.740 ;
  LAYER VI3 ;
  RECT 2040.500 6.340 2040.700 6.540 ;
  LAYER VI3 ;
  RECT 2040.500 5.940 2040.700 6.140 ;
  LAYER VI3 ;
  RECT 2040.100 6.340 2040.300 6.540 ;
  LAYER VI3 ;
  RECT 2040.100 5.940 2040.300 6.140 ;
  LAYER VI3 ;
  RECT 2039.700 6.340 2039.900 6.540 ;
  LAYER VI3 ;
  RECT 2039.700 5.940 2039.900 6.140 ;
  LAYER VI3 ;
  RECT 2039.300 6.340 2039.500 6.540 ;
  LAYER VI3 ;
  RECT 2039.300 5.940 2039.500 6.140 ;
  LAYER VI3 ;
  RECT 2038.900 6.340 2039.100 6.540 ;
  LAYER VI3 ;
  RECT 2038.900 5.940 2039.100 6.140 ;
  LAYER VI3 ;
  RECT 2038.500 6.340 2038.700 6.540 ;
  LAYER VI3 ;
  RECT 2038.500 5.940 2038.700 6.140 ;
  LAYER VI3 ;
  RECT 2038.100 6.340 2038.300 6.540 ;
  LAYER VI3 ;
  RECT 2038.100 5.940 2038.300 6.140 ;
  LAYER VI3 ;
  RECT 2037.700 6.340 2037.900 6.540 ;
  LAYER VI3 ;
  RECT 2037.700 5.940 2037.900 6.140 ;
  LAYER VI3 ;
  RECT 2037.300 6.340 2037.500 6.540 ;
  LAYER VI3 ;
  RECT 2037.300 5.940 2037.500 6.140 ;
  LAYER VI3 ;
  RECT 2036.900 6.340 2037.100 6.540 ;
  LAYER VI3 ;
  RECT 2036.900 5.940 2037.100 6.140 ;
  LAYER VI3 ;
  RECT 2036.500 6.340 2036.700 6.540 ;
  LAYER VI3 ;
  RECT 2036.500 5.940 2036.700 6.140 ;
  LAYER VI3 ;
  RECT 2036.100 6.340 2036.300 6.540 ;
  LAYER VI3 ;
  RECT 2036.100 5.940 2036.300 6.140 ;
  LAYER VI3 ;
  RECT 2035.700 6.340 2035.900 6.540 ;
  LAYER VI3 ;
  RECT 2035.700 5.940 2035.900 6.140 ;
  LAYER VI3 ;
  RECT 2035.300 6.340 2035.500 6.540 ;
  LAYER VI3 ;
  RECT 2035.300 5.940 2035.500 6.140 ;
  LAYER VI3 ;
  RECT 2034.900 6.340 2035.100 6.540 ;
  LAYER VI3 ;
  RECT 2034.900 5.940 2035.100 6.140 ;
  LAYER VI3 ;
  RECT 2034.500 6.340 2034.700 6.540 ;
  LAYER VI3 ;
  RECT 2034.500 5.940 2034.700 6.140 ;
  LAYER VI3 ;
  RECT 2034.100 6.340 2034.300 6.540 ;
  LAYER VI3 ;
  RECT 2034.100 5.940 2034.300 6.140 ;
  LAYER VI3 ;
  RECT 2033.700 6.340 2033.900 6.540 ;
  LAYER VI3 ;
  RECT 2033.700 5.940 2033.900 6.140 ;
  LAYER VI3 ;
  RECT 2033.300 6.340 2033.500 6.540 ;
  LAYER VI3 ;
  RECT 2033.300 5.940 2033.500 6.140 ;
  LAYER VI3 ;
  RECT 2032.900 6.340 2033.100 6.540 ;
  LAYER VI3 ;
  RECT 2032.900 5.940 2033.100 6.140 ;
  LAYER VI3 ;
  RECT 2052.740 5.880 2060.740 6.740 ;
  LAYER VI3 ;
  RECT 2060.340 6.340 2060.540 6.540 ;
  LAYER VI3 ;
  RECT 2060.340 5.940 2060.540 6.140 ;
  LAYER VI3 ;
  RECT 2059.940 6.340 2060.140 6.540 ;
  LAYER VI3 ;
  RECT 2059.940 5.940 2060.140 6.140 ;
  LAYER VI3 ;
  RECT 2059.540 6.340 2059.740 6.540 ;
  LAYER VI3 ;
  RECT 2059.540 5.940 2059.740 6.140 ;
  LAYER VI3 ;
  RECT 2059.140 6.340 2059.340 6.540 ;
  LAYER VI3 ;
  RECT 2059.140 5.940 2059.340 6.140 ;
  LAYER VI3 ;
  RECT 2058.740 6.340 2058.940 6.540 ;
  LAYER VI3 ;
  RECT 2058.740 5.940 2058.940 6.140 ;
  LAYER VI3 ;
  RECT 2058.340 6.340 2058.540 6.540 ;
  LAYER VI3 ;
  RECT 2058.340 5.940 2058.540 6.140 ;
  LAYER VI3 ;
  RECT 2057.940 6.340 2058.140 6.540 ;
  LAYER VI3 ;
  RECT 2057.940 5.940 2058.140 6.140 ;
  LAYER VI3 ;
  RECT 2057.540 6.340 2057.740 6.540 ;
  LAYER VI3 ;
  RECT 2057.540 5.940 2057.740 6.140 ;
  LAYER VI3 ;
  RECT 2057.140 6.340 2057.340 6.540 ;
  LAYER VI3 ;
  RECT 2057.140 5.940 2057.340 6.140 ;
  LAYER VI3 ;
  RECT 2056.740 6.340 2056.940 6.540 ;
  LAYER VI3 ;
  RECT 2056.740 5.940 2056.940 6.140 ;
  LAYER VI3 ;
  RECT 2056.340 6.340 2056.540 6.540 ;
  LAYER VI3 ;
  RECT 2056.340 5.940 2056.540 6.140 ;
  LAYER VI3 ;
  RECT 2055.940 6.340 2056.140 6.540 ;
  LAYER VI3 ;
  RECT 2055.940 5.940 2056.140 6.140 ;
  LAYER VI3 ;
  RECT 2055.540 6.340 2055.740 6.540 ;
  LAYER VI3 ;
  RECT 2055.540 5.940 2055.740 6.140 ;
  LAYER VI3 ;
  RECT 2055.140 6.340 2055.340 6.540 ;
  LAYER VI3 ;
  RECT 2055.140 5.940 2055.340 6.140 ;
  LAYER VI3 ;
  RECT 2054.740 6.340 2054.940 6.540 ;
  LAYER VI3 ;
  RECT 2054.740 5.940 2054.940 6.140 ;
  LAYER VI3 ;
  RECT 2054.340 6.340 2054.540 6.540 ;
  LAYER VI3 ;
  RECT 2054.340 5.940 2054.540 6.140 ;
  LAYER VI3 ;
  RECT 2053.940 6.340 2054.140 6.540 ;
  LAYER VI3 ;
  RECT 2053.940 5.940 2054.140 6.140 ;
  LAYER VI3 ;
  RECT 2053.540 6.340 2053.740 6.540 ;
  LAYER VI3 ;
  RECT 2053.540 5.940 2053.740 6.140 ;
  LAYER VI3 ;
  RECT 2053.140 6.340 2053.340 6.540 ;
  LAYER VI3 ;
  RECT 2053.140 5.940 2053.340 6.140 ;
  LAYER VI3 ;
  RECT 2052.740 6.340 2052.940 6.540 ;
  LAYER VI3 ;
  RECT 2052.740 5.940 2052.940 6.140 ;
  LAYER VI3 ;
  RECT 2073.820 5.880 2081.820 6.740 ;
  LAYER VI3 ;
  RECT 2081.420 6.340 2081.620 6.540 ;
  LAYER VI3 ;
  RECT 2081.420 5.940 2081.620 6.140 ;
  LAYER VI3 ;
  RECT 2081.020 6.340 2081.220 6.540 ;
  LAYER VI3 ;
  RECT 2081.020 5.940 2081.220 6.140 ;
  LAYER VI3 ;
  RECT 2080.620 6.340 2080.820 6.540 ;
  LAYER VI3 ;
  RECT 2080.620 5.940 2080.820 6.140 ;
  LAYER VI3 ;
  RECT 2080.220 6.340 2080.420 6.540 ;
  LAYER VI3 ;
  RECT 2080.220 5.940 2080.420 6.140 ;
  LAYER VI3 ;
  RECT 2079.820 6.340 2080.020 6.540 ;
  LAYER VI3 ;
  RECT 2079.820 5.940 2080.020 6.140 ;
  LAYER VI3 ;
  RECT 2079.420 6.340 2079.620 6.540 ;
  LAYER VI3 ;
  RECT 2079.420 5.940 2079.620 6.140 ;
  LAYER VI3 ;
  RECT 2079.020 6.340 2079.220 6.540 ;
  LAYER VI3 ;
  RECT 2079.020 5.940 2079.220 6.140 ;
  LAYER VI3 ;
  RECT 2078.620 6.340 2078.820 6.540 ;
  LAYER VI3 ;
  RECT 2078.620 5.940 2078.820 6.140 ;
  LAYER VI3 ;
  RECT 2078.220 6.340 2078.420 6.540 ;
  LAYER VI3 ;
  RECT 2078.220 5.940 2078.420 6.140 ;
  LAYER VI3 ;
  RECT 2077.820 6.340 2078.020 6.540 ;
  LAYER VI3 ;
  RECT 2077.820 5.940 2078.020 6.140 ;
  LAYER VI3 ;
  RECT 2077.420 6.340 2077.620 6.540 ;
  LAYER VI3 ;
  RECT 2077.420 5.940 2077.620 6.140 ;
  LAYER VI3 ;
  RECT 2077.020 6.340 2077.220 6.540 ;
  LAYER VI3 ;
  RECT 2077.020 5.940 2077.220 6.140 ;
  LAYER VI3 ;
  RECT 2076.620 6.340 2076.820 6.540 ;
  LAYER VI3 ;
  RECT 2076.620 5.940 2076.820 6.140 ;
  LAYER VI3 ;
  RECT 2076.220 6.340 2076.420 6.540 ;
  LAYER VI3 ;
  RECT 2076.220 5.940 2076.420 6.140 ;
  LAYER VI3 ;
  RECT 2075.820 6.340 2076.020 6.540 ;
  LAYER VI3 ;
  RECT 2075.820 5.940 2076.020 6.140 ;
  LAYER VI3 ;
  RECT 2075.420 6.340 2075.620 6.540 ;
  LAYER VI3 ;
  RECT 2075.420 5.940 2075.620 6.140 ;
  LAYER VI3 ;
  RECT 2075.020 6.340 2075.220 6.540 ;
  LAYER VI3 ;
  RECT 2075.020 5.940 2075.220 6.140 ;
  LAYER VI3 ;
  RECT 2074.620 6.340 2074.820 6.540 ;
  LAYER VI3 ;
  RECT 2074.620 5.940 2074.820 6.140 ;
  LAYER VI3 ;
  RECT 2074.220 6.340 2074.420 6.540 ;
  LAYER VI3 ;
  RECT 2074.220 5.940 2074.420 6.140 ;
  LAYER VI3 ;
  RECT 2073.820 6.340 2074.020 6.540 ;
  LAYER VI3 ;
  RECT 2073.820 5.940 2074.020 6.140 ;
  LAYER VI3 ;
  RECT 2093.660 5.880 2101.660 6.740 ;
  LAYER VI3 ;
  RECT 2101.260 6.340 2101.460 6.540 ;
  LAYER VI3 ;
  RECT 2101.260 5.940 2101.460 6.140 ;
  LAYER VI3 ;
  RECT 2100.860 6.340 2101.060 6.540 ;
  LAYER VI3 ;
  RECT 2100.860 5.940 2101.060 6.140 ;
  LAYER VI3 ;
  RECT 2100.460 6.340 2100.660 6.540 ;
  LAYER VI3 ;
  RECT 2100.460 5.940 2100.660 6.140 ;
  LAYER VI3 ;
  RECT 2100.060 6.340 2100.260 6.540 ;
  LAYER VI3 ;
  RECT 2100.060 5.940 2100.260 6.140 ;
  LAYER VI3 ;
  RECT 2099.660 6.340 2099.860 6.540 ;
  LAYER VI3 ;
  RECT 2099.660 5.940 2099.860 6.140 ;
  LAYER VI3 ;
  RECT 2099.260 6.340 2099.460 6.540 ;
  LAYER VI3 ;
  RECT 2099.260 5.940 2099.460 6.140 ;
  LAYER VI3 ;
  RECT 2098.860 6.340 2099.060 6.540 ;
  LAYER VI3 ;
  RECT 2098.860 5.940 2099.060 6.140 ;
  LAYER VI3 ;
  RECT 2098.460 6.340 2098.660 6.540 ;
  LAYER VI3 ;
  RECT 2098.460 5.940 2098.660 6.140 ;
  LAYER VI3 ;
  RECT 2098.060 6.340 2098.260 6.540 ;
  LAYER VI3 ;
  RECT 2098.060 5.940 2098.260 6.140 ;
  LAYER VI3 ;
  RECT 2097.660 6.340 2097.860 6.540 ;
  LAYER VI3 ;
  RECT 2097.660 5.940 2097.860 6.140 ;
  LAYER VI3 ;
  RECT 2097.260 6.340 2097.460 6.540 ;
  LAYER VI3 ;
  RECT 2097.260 5.940 2097.460 6.140 ;
  LAYER VI3 ;
  RECT 2096.860 6.340 2097.060 6.540 ;
  LAYER VI3 ;
  RECT 2096.860 5.940 2097.060 6.140 ;
  LAYER VI3 ;
  RECT 2096.460 6.340 2096.660 6.540 ;
  LAYER VI3 ;
  RECT 2096.460 5.940 2096.660 6.140 ;
  LAYER VI3 ;
  RECT 2096.060 6.340 2096.260 6.540 ;
  LAYER VI3 ;
  RECT 2096.060 5.940 2096.260 6.140 ;
  LAYER VI3 ;
  RECT 2095.660 6.340 2095.860 6.540 ;
  LAYER VI3 ;
  RECT 2095.660 5.940 2095.860 6.140 ;
  LAYER VI3 ;
  RECT 2095.260 6.340 2095.460 6.540 ;
  LAYER VI3 ;
  RECT 2095.260 5.940 2095.460 6.140 ;
  LAYER VI3 ;
  RECT 2094.860 6.340 2095.060 6.540 ;
  LAYER VI3 ;
  RECT 2094.860 5.940 2095.060 6.140 ;
  LAYER VI3 ;
  RECT 2094.460 6.340 2094.660 6.540 ;
  LAYER VI3 ;
  RECT 2094.460 5.940 2094.660 6.140 ;
  LAYER VI3 ;
  RECT 2094.060 6.340 2094.260 6.540 ;
  LAYER VI3 ;
  RECT 2094.060 5.940 2094.260 6.140 ;
  LAYER VI3 ;
  RECT 2093.660 6.340 2093.860 6.540 ;
  LAYER VI3 ;
  RECT 2093.660 5.940 2093.860 6.140 ;
  LAYER VI3 ;
  RECT 2114.740 5.880 2122.740 6.740 ;
  LAYER VI3 ;
  RECT 2122.340 6.340 2122.540 6.540 ;
  LAYER VI3 ;
  RECT 2122.340 5.940 2122.540 6.140 ;
  LAYER VI3 ;
  RECT 2121.940 6.340 2122.140 6.540 ;
  LAYER VI3 ;
  RECT 2121.940 5.940 2122.140 6.140 ;
  LAYER VI3 ;
  RECT 2121.540 6.340 2121.740 6.540 ;
  LAYER VI3 ;
  RECT 2121.540 5.940 2121.740 6.140 ;
  LAYER VI3 ;
  RECT 2121.140 6.340 2121.340 6.540 ;
  LAYER VI3 ;
  RECT 2121.140 5.940 2121.340 6.140 ;
  LAYER VI3 ;
  RECT 2120.740 6.340 2120.940 6.540 ;
  LAYER VI3 ;
  RECT 2120.740 5.940 2120.940 6.140 ;
  LAYER VI3 ;
  RECT 2120.340 6.340 2120.540 6.540 ;
  LAYER VI3 ;
  RECT 2120.340 5.940 2120.540 6.140 ;
  LAYER VI3 ;
  RECT 2119.940 6.340 2120.140 6.540 ;
  LAYER VI3 ;
  RECT 2119.940 5.940 2120.140 6.140 ;
  LAYER VI3 ;
  RECT 2119.540 6.340 2119.740 6.540 ;
  LAYER VI3 ;
  RECT 2119.540 5.940 2119.740 6.140 ;
  LAYER VI3 ;
  RECT 2119.140 6.340 2119.340 6.540 ;
  LAYER VI3 ;
  RECT 2119.140 5.940 2119.340 6.140 ;
  LAYER VI3 ;
  RECT 2118.740 6.340 2118.940 6.540 ;
  LAYER VI3 ;
  RECT 2118.740 5.940 2118.940 6.140 ;
  LAYER VI3 ;
  RECT 2118.340 6.340 2118.540 6.540 ;
  LAYER VI3 ;
  RECT 2118.340 5.940 2118.540 6.140 ;
  LAYER VI3 ;
  RECT 2117.940 6.340 2118.140 6.540 ;
  LAYER VI3 ;
  RECT 2117.940 5.940 2118.140 6.140 ;
  LAYER VI3 ;
  RECT 2117.540 6.340 2117.740 6.540 ;
  LAYER VI3 ;
  RECT 2117.540 5.940 2117.740 6.140 ;
  LAYER VI3 ;
  RECT 2117.140 6.340 2117.340 6.540 ;
  LAYER VI3 ;
  RECT 2117.140 5.940 2117.340 6.140 ;
  LAYER VI3 ;
  RECT 2116.740 6.340 2116.940 6.540 ;
  LAYER VI3 ;
  RECT 2116.740 5.940 2116.940 6.140 ;
  LAYER VI3 ;
  RECT 2116.340 6.340 2116.540 6.540 ;
  LAYER VI3 ;
  RECT 2116.340 5.940 2116.540 6.140 ;
  LAYER VI3 ;
  RECT 2115.940 6.340 2116.140 6.540 ;
  LAYER VI3 ;
  RECT 2115.940 5.940 2116.140 6.140 ;
  LAYER VI3 ;
  RECT 2115.540 6.340 2115.740 6.540 ;
  LAYER VI3 ;
  RECT 2115.540 5.940 2115.740 6.140 ;
  LAYER VI3 ;
  RECT 2115.140 6.340 2115.340 6.540 ;
  LAYER VI3 ;
  RECT 2115.140 5.940 2115.340 6.140 ;
  LAYER VI3 ;
  RECT 2114.740 6.340 2114.940 6.540 ;
  LAYER VI3 ;
  RECT 2114.740 5.940 2114.940 6.140 ;
  LAYER VI3 ;
  RECT 2134.580 5.880 2142.580 6.740 ;
  LAYER VI3 ;
  RECT 2142.180 6.340 2142.380 6.540 ;
  LAYER VI3 ;
  RECT 2142.180 5.940 2142.380 6.140 ;
  LAYER VI3 ;
  RECT 2141.780 6.340 2141.980 6.540 ;
  LAYER VI3 ;
  RECT 2141.780 5.940 2141.980 6.140 ;
  LAYER VI3 ;
  RECT 2141.380 6.340 2141.580 6.540 ;
  LAYER VI3 ;
  RECT 2141.380 5.940 2141.580 6.140 ;
  LAYER VI3 ;
  RECT 2140.980 6.340 2141.180 6.540 ;
  LAYER VI3 ;
  RECT 2140.980 5.940 2141.180 6.140 ;
  LAYER VI3 ;
  RECT 2140.580 6.340 2140.780 6.540 ;
  LAYER VI3 ;
  RECT 2140.580 5.940 2140.780 6.140 ;
  LAYER VI3 ;
  RECT 2140.180 6.340 2140.380 6.540 ;
  LAYER VI3 ;
  RECT 2140.180 5.940 2140.380 6.140 ;
  LAYER VI3 ;
  RECT 2139.780 6.340 2139.980 6.540 ;
  LAYER VI3 ;
  RECT 2139.780 5.940 2139.980 6.140 ;
  LAYER VI3 ;
  RECT 2139.380 6.340 2139.580 6.540 ;
  LAYER VI3 ;
  RECT 2139.380 5.940 2139.580 6.140 ;
  LAYER VI3 ;
  RECT 2138.980 6.340 2139.180 6.540 ;
  LAYER VI3 ;
  RECT 2138.980 5.940 2139.180 6.140 ;
  LAYER VI3 ;
  RECT 2138.580 6.340 2138.780 6.540 ;
  LAYER VI3 ;
  RECT 2138.580 5.940 2138.780 6.140 ;
  LAYER VI3 ;
  RECT 2138.180 6.340 2138.380 6.540 ;
  LAYER VI3 ;
  RECT 2138.180 5.940 2138.380 6.140 ;
  LAYER VI3 ;
  RECT 2137.780 6.340 2137.980 6.540 ;
  LAYER VI3 ;
  RECT 2137.780 5.940 2137.980 6.140 ;
  LAYER VI3 ;
  RECT 2137.380 6.340 2137.580 6.540 ;
  LAYER VI3 ;
  RECT 2137.380 5.940 2137.580 6.140 ;
  LAYER VI3 ;
  RECT 2136.980 6.340 2137.180 6.540 ;
  LAYER VI3 ;
  RECT 2136.980 5.940 2137.180 6.140 ;
  LAYER VI3 ;
  RECT 2136.580 6.340 2136.780 6.540 ;
  LAYER VI3 ;
  RECT 2136.580 5.940 2136.780 6.140 ;
  LAYER VI3 ;
  RECT 2136.180 6.340 2136.380 6.540 ;
  LAYER VI3 ;
  RECT 2136.180 5.940 2136.380 6.140 ;
  LAYER VI3 ;
  RECT 2135.780 6.340 2135.980 6.540 ;
  LAYER VI3 ;
  RECT 2135.780 5.940 2135.980 6.140 ;
  LAYER VI3 ;
  RECT 2135.380 6.340 2135.580 6.540 ;
  LAYER VI3 ;
  RECT 2135.380 5.940 2135.580 6.140 ;
  LAYER VI3 ;
  RECT 2134.980 6.340 2135.180 6.540 ;
  LAYER VI3 ;
  RECT 2134.980 5.940 2135.180 6.140 ;
  LAYER VI3 ;
  RECT 2134.580 6.340 2134.780 6.540 ;
  LAYER VI3 ;
  RECT 2134.580 5.940 2134.780 6.140 ;
  LAYER VI3 ;
  RECT 2155.660 5.880 2163.660 6.740 ;
  LAYER VI3 ;
  RECT 2163.260 6.340 2163.460 6.540 ;
  LAYER VI3 ;
  RECT 2163.260 5.940 2163.460 6.140 ;
  LAYER VI3 ;
  RECT 2162.860 6.340 2163.060 6.540 ;
  LAYER VI3 ;
  RECT 2162.860 5.940 2163.060 6.140 ;
  LAYER VI3 ;
  RECT 2162.460 6.340 2162.660 6.540 ;
  LAYER VI3 ;
  RECT 2162.460 5.940 2162.660 6.140 ;
  LAYER VI3 ;
  RECT 2162.060 6.340 2162.260 6.540 ;
  LAYER VI3 ;
  RECT 2162.060 5.940 2162.260 6.140 ;
  LAYER VI3 ;
  RECT 2161.660 6.340 2161.860 6.540 ;
  LAYER VI3 ;
  RECT 2161.660 5.940 2161.860 6.140 ;
  LAYER VI3 ;
  RECT 2161.260 6.340 2161.460 6.540 ;
  LAYER VI3 ;
  RECT 2161.260 5.940 2161.460 6.140 ;
  LAYER VI3 ;
  RECT 2160.860 6.340 2161.060 6.540 ;
  LAYER VI3 ;
  RECT 2160.860 5.940 2161.060 6.140 ;
  LAYER VI3 ;
  RECT 2160.460 6.340 2160.660 6.540 ;
  LAYER VI3 ;
  RECT 2160.460 5.940 2160.660 6.140 ;
  LAYER VI3 ;
  RECT 2160.060 6.340 2160.260 6.540 ;
  LAYER VI3 ;
  RECT 2160.060 5.940 2160.260 6.140 ;
  LAYER VI3 ;
  RECT 2159.660 6.340 2159.860 6.540 ;
  LAYER VI3 ;
  RECT 2159.660 5.940 2159.860 6.140 ;
  LAYER VI3 ;
  RECT 2159.260 6.340 2159.460 6.540 ;
  LAYER VI3 ;
  RECT 2159.260 5.940 2159.460 6.140 ;
  LAYER VI3 ;
  RECT 2158.860 6.340 2159.060 6.540 ;
  LAYER VI3 ;
  RECT 2158.860 5.940 2159.060 6.140 ;
  LAYER VI3 ;
  RECT 2158.460 6.340 2158.660 6.540 ;
  LAYER VI3 ;
  RECT 2158.460 5.940 2158.660 6.140 ;
  LAYER VI3 ;
  RECT 2158.060 6.340 2158.260 6.540 ;
  LAYER VI3 ;
  RECT 2158.060 5.940 2158.260 6.140 ;
  LAYER VI3 ;
  RECT 2157.660 6.340 2157.860 6.540 ;
  LAYER VI3 ;
  RECT 2157.660 5.940 2157.860 6.140 ;
  LAYER VI3 ;
  RECT 2157.260 6.340 2157.460 6.540 ;
  LAYER VI3 ;
  RECT 2157.260 5.940 2157.460 6.140 ;
  LAYER VI3 ;
  RECT 2156.860 6.340 2157.060 6.540 ;
  LAYER VI3 ;
  RECT 2156.860 5.940 2157.060 6.140 ;
  LAYER VI3 ;
  RECT 2156.460 6.340 2156.660 6.540 ;
  LAYER VI3 ;
  RECT 2156.460 5.940 2156.660 6.140 ;
  LAYER VI3 ;
  RECT 2156.060 6.340 2156.260 6.540 ;
  LAYER VI3 ;
  RECT 2156.060 5.940 2156.260 6.140 ;
  LAYER VI3 ;
  RECT 2155.660 6.340 2155.860 6.540 ;
  LAYER VI3 ;
  RECT 2155.660 5.940 2155.860 6.140 ;
  LAYER VI3 ;
  RECT 2175.500 5.880 2183.500 6.740 ;
  LAYER VI3 ;
  RECT 2183.100 6.340 2183.300 6.540 ;
  LAYER VI3 ;
  RECT 2183.100 5.940 2183.300 6.140 ;
  LAYER VI3 ;
  RECT 2182.700 6.340 2182.900 6.540 ;
  LAYER VI3 ;
  RECT 2182.700 5.940 2182.900 6.140 ;
  LAYER VI3 ;
  RECT 2182.300 6.340 2182.500 6.540 ;
  LAYER VI3 ;
  RECT 2182.300 5.940 2182.500 6.140 ;
  LAYER VI3 ;
  RECT 2181.900 6.340 2182.100 6.540 ;
  LAYER VI3 ;
  RECT 2181.900 5.940 2182.100 6.140 ;
  LAYER VI3 ;
  RECT 2181.500 6.340 2181.700 6.540 ;
  LAYER VI3 ;
  RECT 2181.500 5.940 2181.700 6.140 ;
  LAYER VI3 ;
  RECT 2181.100 6.340 2181.300 6.540 ;
  LAYER VI3 ;
  RECT 2181.100 5.940 2181.300 6.140 ;
  LAYER VI3 ;
  RECT 2180.700 6.340 2180.900 6.540 ;
  LAYER VI3 ;
  RECT 2180.700 5.940 2180.900 6.140 ;
  LAYER VI3 ;
  RECT 2180.300 6.340 2180.500 6.540 ;
  LAYER VI3 ;
  RECT 2180.300 5.940 2180.500 6.140 ;
  LAYER VI3 ;
  RECT 2179.900 6.340 2180.100 6.540 ;
  LAYER VI3 ;
  RECT 2179.900 5.940 2180.100 6.140 ;
  LAYER VI3 ;
  RECT 2179.500 6.340 2179.700 6.540 ;
  LAYER VI3 ;
  RECT 2179.500 5.940 2179.700 6.140 ;
  LAYER VI3 ;
  RECT 2179.100 6.340 2179.300 6.540 ;
  LAYER VI3 ;
  RECT 2179.100 5.940 2179.300 6.140 ;
  LAYER VI3 ;
  RECT 2178.700 6.340 2178.900 6.540 ;
  LAYER VI3 ;
  RECT 2178.700 5.940 2178.900 6.140 ;
  LAYER VI3 ;
  RECT 2178.300 6.340 2178.500 6.540 ;
  LAYER VI3 ;
  RECT 2178.300 5.940 2178.500 6.140 ;
  LAYER VI3 ;
  RECT 2177.900 6.340 2178.100 6.540 ;
  LAYER VI3 ;
  RECT 2177.900 5.940 2178.100 6.140 ;
  LAYER VI3 ;
  RECT 2177.500 6.340 2177.700 6.540 ;
  LAYER VI3 ;
  RECT 2177.500 5.940 2177.700 6.140 ;
  LAYER VI3 ;
  RECT 2177.100 6.340 2177.300 6.540 ;
  LAYER VI3 ;
  RECT 2177.100 5.940 2177.300 6.140 ;
  LAYER VI3 ;
  RECT 2176.700 6.340 2176.900 6.540 ;
  LAYER VI3 ;
  RECT 2176.700 5.940 2176.900 6.140 ;
  LAYER VI3 ;
  RECT 2176.300 6.340 2176.500 6.540 ;
  LAYER VI3 ;
  RECT 2176.300 5.940 2176.500 6.140 ;
  LAYER VI3 ;
  RECT 2175.900 6.340 2176.100 6.540 ;
  LAYER VI3 ;
  RECT 2175.900 5.940 2176.100 6.140 ;
  LAYER VI3 ;
  RECT 2175.500 6.340 2175.700 6.540 ;
  LAYER VI3 ;
  RECT 2175.500 5.940 2175.700 6.140 ;
  LAYER VI3 ;
  RECT 2196.580 5.880 2204.580 6.740 ;
  LAYER VI3 ;
  RECT 2204.180 6.340 2204.380 6.540 ;
  LAYER VI3 ;
  RECT 2204.180 5.940 2204.380 6.140 ;
  LAYER VI3 ;
  RECT 2203.780 6.340 2203.980 6.540 ;
  LAYER VI3 ;
  RECT 2203.780 5.940 2203.980 6.140 ;
  LAYER VI3 ;
  RECT 2203.380 6.340 2203.580 6.540 ;
  LAYER VI3 ;
  RECT 2203.380 5.940 2203.580 6.140 ;
  LAYER VI3 ;
  RECT 2202.980 6.340 2203.180 6.540 ;
  LAYER VI3 ;
  RECT 2202.980 5.940 2203.180 6.140 ;
  LAYER VI3 ;
  RECT 2202.580 6.340 2202.780 6.540 ;
  LAYER VI3 ;
  RECT 2202.580 5.940 2202.780 6.140 ;
  LAYER VI3 ;
  RECT 2202.180 6.340 2202.380 6.540 ;
  LAYER VI3 ;
  RECT 2202.180 5.940 2202.380 6.140 ;
  LAYER VI3 ;
  RECT 2201.780 6.340 2201.980 6.540 ;
  LAYER VI3 ;
  RECT 2201.780 5.940 2201.980 6.140 ;
  LAYER VI3 ;
  RECT 2201.380 6.340 2201.580 6.540 ;
  LAYER VI3 ;
  RECT 2201.380 5.940 2201.580 6.140 ;
  LAYER VI3 ;
  RECT 2200.980 6.340 2201.180 6.540 ;
  LAYER VI3 ;
  RECT 2200.980 5.940 2201.180 6.140 ;
  LAYER VI3 ;
  RECT 2200.580 6.340 2200.780 6.540 ;
  LAYER VI3 ;
  RECT 2200.580 5.940 2200.780 6.140 ;
  LAYER VI3 ;
  RECT 2200.180 6.340 2200.380 6.540 ;
  LAYER VI3 ;
  RECT 2200.180 5.940 2200.380 6.140 ;
  LAYER VI3 ;
  RECT 2199.780 6.340 2199.980 6.540 ;
  LAYER VI3 ;
  RECT 2199.780 5.940 2199.980 6.140 ;
  LAYER VI3 ;
  RECT 2199.380 6.340 2199.580 6.540 ;
  LAYER VI3 ;
  RECT 2199.380 5.940 2199.580 6.140 ;
  LAYER VI3 ;
  RECT 2198.980 6.340 2199.180 6.540 ;
  LAYER VI3 ;
  RECT 2198.980 5.940 2199.180 6.140 ;
  LAYER VI3 ;
  RECT 2198.580 6.340 2198.780 6.540 ;
  LAYER VI3 ;
  RECT 2198.580 5.940 2198.780 6.140 ;
  LAYER VI3 ;
  RECT 2198.180 6.340 2198.380 6.540 ;
  LAYER VI3 ;
  RECT 2198.180 5.940 2198.380 6.140 ;
  LAYER VI3 ;
  RECT 2197.780 6.340 2197.980 6.540 ;
  LAYER VI3 ;
  RECT 2197.780 5.940 2197.980 6.140 ;
  LAYER VI3 ;
  RECT 2197.380 6.340 2197.580 6.540 ;
  LAYER VI3 ;
  RECT 2197.380 5.940 2197.580 6.140 ;
  LAYER VI3 ;
  RECT 2196.980 6.340 2197.180 6.540 ;
  LAYER VI3 ;
  RECT 2196.980 5.940 2197.180 6.140 ;
  LAYER VI3 ;
  RECT 2196.580 6.340 2196.780 6.540 ;
  LAYER VI3 ;
  RECT 2196.580 5.940 2196.780 6.140 ;
  LAYER VI3 ;
  RECT 2216.420 5.880 2224.420 6.740 ;
  LAYER VI3 ;
  RECT 2224.020 6.340 2224.220 6.540 ;
  LAYER VI3 ;
  RECT 2224.020 5.940 2224.220 6.140 ;
  LAYER VI3 ;
  RECT 2223.620 6.340 2223.820 6.540 ;
  LAYER VI3 ;
  RECT 2223.620 5.940 2223.820 6.140 ;
  LAYER VI3 ;
  RECT 2223.220 6.340 2223.420 6.540 ;
  LAYER VI3 ;
  RECT 2223.220 5.940 2223.420 6.140 ;
  LAYER VI3 ;
  RECT 2222.820 6.340 2223.020 6.540 ;
  LAYER VI3 ;
  RECT 2222.820 5.940 2223.020 6.140 ;
  LAYER VI3 ;
  RECT 2222.420 6.340 2222.620 6.540 ;
  LAYER VI3 ;
  RECT 2222.420 5.940 2222.620 6.140 ;
  LAYER VI3 ;
  RECT 2222.020 6.340 2222.220 6.540 ;
  LAYER VI3 ;
  RECT 2222.020 5.940 2222.220 6.140 ;
  LAYER VI3 ;
  RECT 2221.620 6.340 2221.820 6.540 ;
  LAYER VI3 ;
  RECT 2221.620 5.940 2221.820 6.140 ;
  LAYER VI3 ;
  RECT 2221.220 6.340 2221.420 6.540 ;
  LAYER VI3 ;
  RECT 2221.220 5.940 2221.420 6.140 ;
  LAYER VI3 ;
  RECT 2220.820 6.340 2221.020 6.540 ;
  LAYER VI3 ;
  RECT 2220.820 5.940 2221.020 6.140 ;
  LAYER VI3 ;
  RECT 2220.420 6.340 2220.620 6.540 ;
  LAYER VI3 ;
  RECT 2220.420 5.940 2220.620 6.140 ;
  LAYER VI3 ;
  RECT 2220.020 6.340 2220.220 6.540 ;
  LAYER VI3 ;
  RECT 2220.020 5.940 2220.220 6.140 ;
  LAYER VI3 ;
  RECT 2219.620 6.340 2219.820 6.540 ;
  LAYER VI3 ;
  RECT 2219.620 5.940 2219.820 6.140 ;
  LAYER VI3 ;
  RECT 2219.220 6.340 2219.420 6.540 ;
  LAYER VI3 ;
  RECT 2219.220 5.940 2219.420 6.140 ;
  LAYER VI3 ;
  RECT 2218.820 6.340 2219.020 6.540 ;
  LAYER VI3 ;
  RECT 2218.820 5.940 2219.020 6.140 ;
  LAYER VI3 ;
  RECT 2218.420 6.340 2218.620 6.540 ;
  LAYER VI3 ;
  RECT 2218.420 5.940 2218.620 6.140 ;
  LAYER VI3 ;
  RECT 2218.020 6.340 2218.220 6.540 ;
  LAYER VI3 ;
  RECT 2218.020 5.940 2218.220 6.140 ;
  LAYER VI3 ;
  RECT 2217.620 6.340 2217.820 6.540 ;
  LAYER VI3 ;
  RECT 2217.620 5.940 2217.820 6.140 ;
  LAYER VI3 ;
  RECT 2217.220 6.340 2217.420 6.540 ;
  LAYER VI3 ;
  RECT 2217.220 5.940 2217.420 6.140 ;
  LAYER VI3 ;
  RECT 2216.820 6.340 2217.020 6.540 ;
  LAYER VI3 ;
  RECT 2216.820 5.940 2217.020 6.140 ;
  LAYER VI3 ;
  RECT 2216.420 6.340 2216.620 6.540 ;
  LAYER VI3 ;
  RECT 2216.420 5.940 2216.620 6.140 ;
  LAYER VI3 ;
  RECT 2237.500 5.880 2245.500 6.740 ;
  LAYER VI3 ;
  RECT 2245.100 6.340 2245.300 6.540 ;
  LAYER VI3 ;
  RECT 2245.100 5.940 2245.300 6.140 ;
  LAYER VI3 ;
  RECT 2244.700 6.340 2244.900 6.540 ;
  LAYER VI3 ;
  RECT 2244.700 5.940 2244.900 6.140 ;
  LAYER VI3 ;
  RECT 2244.300 6.340 2244.500 6.540 ;
  LAYER VI3 ;
  RECT 2244.300 5.940 2244.500 6.140 ;
  LAYER VI3 ;
  RECT 2243.900 6.340 2244.100 6.540 ;
  LAYER VI3 ;
  RECT 2243.900 5.940 2244.100 6.140 ;
  LAYER VI3 ;
  RECT 2243.500 6.340 2243.700 6.540 ;
  LAYER VI3 ;
  RECT 2243.500 5.940 2243.700 6.140 ;
  LAYER VI3 ;
  RECT 2243.100 6.340 2243.300 6.540 ;
  LAYER VI3 ;
  RECT 2243.100 5.940 2243.300 6.140 ;
  LAYER VI3 ;
  RECT 2242.700 6.340 2242.900 6.540 ;
  LAYER VI3 ;
  RECT 2242.700 5.940 2242.900 6.140 ;
  LAYER VI3 ;
  RECT 2242.300 6.340 2242.500 6.540 ;
  LAYER VI3 ;
  RECT 2242.300 5.940 2242.500 6.140 ;
  LAYER VI3 ;
  RECT 2241.900 6.340 2242.100 6.540 ;
  LAYER VI3 ;
  RECT 2241.900 5.940 2242.100 6.140 ;
  LAYER VI3 ;
  RECT 2241.500 6.340 2241.700 6.540 ;
  LAYER VI3 ;
  RECT 2241.500 5.940 2241.700 6.140 ;
  LAYER VI3 ;
  RECT 2241.100 6.340 2241.300 6.540 ;
  LAYER VI3 ;
  RECT 2241.100 5.940 2241.300 6.140 ;
  LAYER VI3 ;
  RECT 2240.700 6.340 2240.900 6.540 ;
  LAYER VI3 ;
  RECT 2240.700 5.940 2240.900 6.140 ;
  LAYER VI3 ;
  RECT 2240.300 6.340 2240.500 6.540 ;
  LAYER VI3 ;
  RECT 2240.300 5.940 2240.500 6.140 ;
  LAYER VI3 ;
  RECT 2239.900 6.340 2240.100 6.540 ;
  LAYER VI3 ;
  RECT 2239.900 5.940 2240.100 6.140 ;
  LAYER VI3 ;
  RECT 2239.500 6.340 2239.700 6.540 ;
  LAYER VI3 ;
  RECT 2239.500 5.940 2239.700 6.140 ;
  LAYER VI3 ;
  RECT 2239.100 6.340 2239.300 6.540 ;
  LAYER VI3 ;
  RECT 2239.100 5.940 2239.300 6.140 ;
  LAYER VI3 ;
  RECT 2238.700 6.340 2238.900 6.540 ;
  LAYER VI3 ;
  RECT 2238.700 5.940 2238.900 6.140 ;
  LAYER VI3 ;
  RECT 2238.300 6.340 2238.500 6.540 ;
  LAYER VI3 ;
  RECT 2238.300 5.940 2238.500 6.140 ;
  LAYER VI3 ;
  RECT 2237.900 6.340 2238.100 6.540 ;
  LAYER VI3 ;
  RECT 2237.900 5.940 2238.100 6.140 ;
  LAYER VI3 ;
  RECT 2237.500 6.340 2237.700 6.540 ;
  LAYER VI3 ;
  RECT 2237.500 5.940 2237.700 6.140 ;
  LAYER VI3 ;
  RECT 2257.340 5.880 2265.340 6.740 ;
  LAYER VI3 ;
  RECT 2264.940 6.340 2265.140 6.540 ;
  LAYER VI3 ;
  RECT 2264.940 5.940 2265.140 6.140 ;
  LAYER VI3 ;
  RECT 2264.540 6.340 2264.740 6.540 ;
  LAYER VI3 ;
  RECT 2264.540 5.940 2264.740 6.140 ;
  LAYER VI3 ;
  RECT 2264.140 6.340 2264.340 6.540 ;
  LAYER VI3 ;
  RECT 2264.140 5.940 2264.340 6.140 ;
  LAYER VI3 ;
  RECT 2263.740 6.340 2263.940 6.540 ;
  LAYER VI3 ;
  RECT 2263.740 5.940 2263.940 6.140 ;
  LAYER VI3 ;
  RECT 2263.340 6.340 2263.540 6.540 ;
  LAYER VI3 ;
  RECT 2263.340 5.940 2263.540 6.140 ;
  LAYER VI3 ;
  RECT 2262.940 6.340 2263.140 6.540 ;
  LAYER VI3 ;
  RECT 2262.940 5.940 2263.140 6.140 ;
  LAYER VI3 ;
  RECT 2262.540 6.340 2262.740 6.540 ;
  LAYER VI3 ;
  RECT 2262.540 5.940 2262.740 6.140 ;
  LAYER VI3 ;
  RECT 2262.140 6.340 2262.340 6.540 ;
  LAYER VI3 ;
  RECT 2262.140 5.940 2262.340 6.140 ;
  LAYER VI3 ;
  RECT 2261.740 6.340 2261.940 6.540 ;
  LAYER VI3 ;
  RECT 2261.740 5.940 2261.940 6.140 ;
  LAYER VI3 ;
  RECT 2261.340 6.340 2261.540 6.540 ;
  LAYER VI3 ;
  RECT 2261.340 5.940 2261.540 6.140 ;
  LAYER VI3 ;
  RECT 2260.940 6.340 2261.140 6.540 ;
  LAYER VI3 ;
  RECT 2260.940 5.940 2261.140 6.140 ;
  LAYER VI3 ;
  RECT 2260.540 6.340 2260.740 6.540 ;
  LAYER VI3 ;
  RECT 2260.540 5.940 2260.740 6.140 ;
  LAYER VI3 ;
  RECT 2260.140 6.340 2260.340 6.540 ;
  LAYER VI3 ;
  RECT 2260.140 5.940 2260.340 6.140 ;
  LAYER VI3 ;
  RECT 2259.740 6.340 2259.940 6.540 ;
  LAYER VI3 ;
  RECT 2259.740 5.940 2259.940 6.140 ;
  LAYER VI3 ;
  RECT 2259.340 6.340 2259.540 6.540 ;
  LAYER VI3 ;
  RECT 2259.340 5.940 2259.540 6.140 ;
  LAYER VI3 ;
  RECT 2258.940 6.340 2259.140 6.540 ;
  LAYER VI3 ;
  RECT 2258.940 5.940 2259.140 6.140 ;
  LAYER VI3 ;
  RECT 2258.540 6.340 2258.740 6.540 ;
  LAYER VI3 ;
  RECT 2258.540 5.940 2258.740 6.140 ;
  LAYER VI3 ;
  RECT 2258.140 6.340 2258.340 6.540 ;
  LAYER VI3 ;
  RECT 2258.140 5.940 2258.340 6.140 ;
  LAYER VI3 ;
  RECT 2257.740 6.340 2257.940 6.540 ;
  LAYER VI3 ;
  RECT 2257.740 5.940 2257.940 6.140 ;
  LAYER VI3 ;
  RECT 2257.340 6.340 2257.540 6.540 ;
  LAYER VI3 ;
  RECT 2257.340 5.940 2257.540 6.140 ;
  LAYER VI3 ;
  RECT 2278.420 5.880 2286.420 6.740 ;
  LAYER VI3 ;
  RECT 2286.020 6.340 2286.220 6.540 ;
  LAYER VI3 ;
  RECT 2286.020 5.940 2286.220 6.140 ;
  LAYER VI3 ;
  RECT 2285.620 6.340 2285.820 6.540 ;
  LAYER VI3 ;
  RECT 2285.620 5.940 2285.820 6.140 ;
  LAYER VI3 ;
  RECT 2285.220 6.340 2285.420 6.540 ;
  LAYER VI3 ;
  RECT 2285.220 5.940 2285.420 6.140 ;
  LAYER VI3 ;
  RECT 2284.820 6.340 2285.020 6.540 ;
  LAYER VI3 ;
  RECT 2284.820 5.940 2285.020 6.140 ;
  LAYER VI3 ;
  RECT 2284.420 6.340 2284.620 6.540 ;
  LAYER VI3 ;
  RECT 2284.420 5.940 2284.620 6.140 ;
  LAYER VI3 ;
  RECT 2284.020 6.340 2284.220 6.540 ;
  LAYER VI3 ;
  RECT 2284.020 5.940 2284.220 6.140 ;
  LAYER VI3 ;
  RECT 2283.620 6.340 2283.820 6.540 ;
  LAYER VI3 ;
  RECT 2283.620 5.940 2283.820 6.140 ;
  LAYER VI3 ;
  RECT 2283.220 6.340 2283.420 6.540 ;
  LAYER VI3 ;
  RECT 2283.220 5.940 2283.420 6.140 ;
  LAYER VI3 ;
  RECT 2282.820 6.340 2283.020 6.540 ;
  LAYER VI3 ;
  RECT 2282.820 5.940 2283.020 6.140 ;
  LAYER VI3 ;
  RECT 2282.420 6.340 2282.620 6.540 ;
  LAYER VI3 ;
  RECT 2282.420 5.940 2282.620 6.140 ;
  LAYER VI3 ;
  RECT 2282.020 6.340 2282.220 6.540 ;
  LAYER VI3 ;
  RECT 2282.020 5.940 2282.220 6.140 ;
  LAYER VI3 ;
  RECT 2281.620 6.340 2281.820 6.540 ;
  LAYER VI3 ;
  RECT 2281.620 5.940 2281.820 6.140 ;
  LAYER VI3 ;
  RECT 2281.220 6.340 2281.420 6.540 ;
  LAYER VI3 ;
  RECT 2281.220 5.940 2281.420 6.140 ;
  LAYER VI3 ;
  RECT 2280.820 6.340 2281.020 6.540 ;
  LAYER VI3 ;
  RECT 2280.820 5.940 2281.020 6.140 ;
  LAYER VI3 ;
  RECT 2280.420 6.340 2280.620 6.540 ;
  LAYER VI3 ;
  RECT 2280.420 5.940 2280.620 6.140 ;
  LAYER VI3 ;
  RECT 2280.020 6.340 2280.220 6.540 ;
  LAYER VI3 ;
  RECT 2280.020 5.940 2280.220 6.140 ;
  LAYER VI3 ;
  RECT 2279.620 6.340 2279.820 6.540 ;
  LAYER VI3 ;
  RECT 2279.620 5.940 2279.820 6.140 ;
  LAYER VI3 ;
  RECT 2279.220 6.340 2279.420 6.540 ;
  LAYER VI3 ;
  RECT 2279.220 5.940 2279.420 6.140 ;
  LAYER VI3 ;
  RECT 2278.820 6.340 2279.020 6.540 ;
  LAYER VI3 ;
  RECT 2278.820 5.940 2279.020 6.140 ;
  LAYER VI3 ;
  RECT 2278.420 6.340 2278.620 6.540 ;
  LAYER VI3 ;
  RECT 2278.420 5.940 2278.620 6.140 ;
  LAYER VI3 ;
  RECT 2298.260 5.880 2306.260 6.740 ;
  LAYER VI3 ;
  RECT 2305.860 6.340 2306.060 6.540 ;
  LAYER VI3 ;
  RECT 2305.860 5.940 2306.060 6.140 ;
  LAYER VI3 ;
  RECT 2305.460 6.340 2305.660 6.540 ;
  LAYER VI3 ;
  RECT 2305.460 5.940 2305.660 6.140 ;
  LAYER VI3 ;
  RECT 2305.060 6.340 2305.260 6.540 ;
  LAYER VI3 ;
  RECT 2305.060 5.940 2305.260 6.140 ;
  LAYER VI3 ;
  RECT 2304.660 6.340 2304.860 6.540 ;
  LAYER VI3 ;
  RECT 2304.660 5.940 2304.860 6.140 ;
  LAYER VI3 ;
  RECT 2304.260 6.340 2304.460 6.540 ;
  LAYER VI3 ;
  RECT 2304.260 5.940 2304.460 6.140 ;
  LAYER VI3 ;
  RECT 2303.860 6.340 2304.060 6.540 ;
  LAYER VI3 ;
  RECT 2303.860 5.940 2304.060 6.140 ;
  LAYER VI3 ;
  RECT 2303.460 6.340 2303.660 6.540 ;
  LAYER VI3 ;
  RECT 2303.460 5.940 2303.660 6.140 ;
  LAYER VI3 ;
  RECT 2303.060 6.340 2303.260 6.540 ;
  LAYER VI3 ;
  RECT 2303.060 5.940 2303.260 6.140 ;
  LAYER VI3 ;
  RECT 2302.660 6.340 2302.860 6.540 ;
  LAYER VI3 ;
  RECT 2302.660 5.940 2302.860 6.140 ;
  LAYER VI3 ;
  RECT 2302.260 6.340 2302.460 6.540 ;
  LAYER VI3 ;
  RECT 2302.260 5.940 2302.460 6.140 ;
  LAYER VI3 ;
  RECT 2301.860 6.340 2302.060 6.540 ;
  LAYER VI3 ;
  RECT 2301.860 5.940 2302.060 6.140 ;
  LAYER VI3 ;
  RECT 2301.460 6.340 2301.660 6.540 ;
  LAYER VI3 ;
  RECT 2301.460 5.940 2301.660 6.140 ;
  LAYER VI3 ;
  RECT 2301.060 6.340 2301.260 6.540 ;
  LAYER VI3 ;
  RECT 2301.060 5.940 2301.260 6.140 ;
  LAYER VI3 ;
  RECT 2300.660 6.340 2300.860 6.540 ;
  LAYER VI3 ;
  RECT 2300.660 5.940 2300.860 6.140 ;
  LAYER VI3 ;
  RECT 2300.260 6.340 2300.460 6.540 ;
  LAYER VI3 ;
  RECT 2300.260 5.940 2300.460 6.140 ;
  LAYER VI3 ;
  RECT 2299.860 6.340 2300.060 6.540 ;
  LAYER VI3 ;
  RECT 2299.860 5.940 2300.060 6.140 ;
  LAYER VI3 ;
  RECT 2299.460 6.340 2299.660 6.540 ;
  LAYER VI3 ;
  RECT 2299.460 5.940 2299.660 6.140 ;
  LAYER VI3 ;
  RECT 2299.060 6.340 2299.260 6.540 ;
  LAYER VI3 ;
  RECT 2299.060 5.940 2299.260 6.140 ;
  LAYER VI3 ;
  RECT 2298.660 6.340 2298.860 6.540 ;
  LAYER VI3 ;
  RECT 2298.660 5.940 2298.860 6.140 ;
  LAYER VI3 ;
  RECT 2298.260 6.340 2298.460 6.540 ;
  LAYER VI3 ;
  RECT 2298.260 5.940 2298.460 6.140 ;
  LAYER VI3 ;
  RECT 2319.340 5.880 2327.340 6.740 ;
  LAYER VI3 ;
  RECT 2326.940 6.340 2327.140 6.540 ;
  LAYER VI3 ;
  RECT 2326.940 5.940 2327.140 6.140 ;
  LAYER VI3 ;
  RECT 2326.540 6.340 2326.740 6.540 ;
  LAYER VI3 ;
  RECT 2326.540 5.940 2326.740 6.140 ;
  LAYER VI3 ;
  RECT 2326.140 6.340 2326.340 6.540 ;
  LAYER VI3 ;
  RECT 2326.140 5.940 2326.340 6.140 ;
  LAYER VI3 ;
  RECT 2325.740 6.340 2325.940 6.540 ;
  LAYER VI3 ;
  RECT 2325.740 5.940 2325.940 6.140 ;
  LAYER VI3 ;
  RECT 2325.340 6.340 2325.540 6.540 ;
  LAYER VI3 ;
  RECT 2325.340 5.940 2325.540 6.140 ;
  LAYER VI3 ;
  RECT 2324.940 6.340 2325.140 6.540 ;
  LAYER VI3 ;
  RECT 2324.940 5.940 2325.140 6.140 ;
  LAYER VI3 ;
  RECT 2324.540 6.340 2324.740 6.540 ;
  LAYER VI3 ;
  RECT 2324.540 5.940 2324.740 6.140 ;
  LAYER VI3 ;
  RECT 2324.140 6.340 2324.340 6.540 ;
  LAYER VI3 ;
  RECT 2324.140 5.940 2324.340 6.140 ;
  LAYER VI3 ;
  RECT 2323.740 6.340 2323.940 6.540 ;
  LAYER VI3 ;
  RECT 2323.740 5.940 2323.940 6.140 ;
  LAYER VI3 ;
  RECT 2323.340 6.340 2323.540 6.540 ;
  LAYER VI3 ;
  RECT 2323.340 5.940 2323.540 6.140 ;
  LAYER VI3 ;
  RECT 2322.940 6.340 2323.140 6.540 ;
  LAYER VI3 ;
  RECT 2322.940 5.940 2323.140 6.140 ;
  LAYER VI3 ;
  RECT 2322.540 6.340 2322.740 6.540 ;
  LAYER VI3 ;
  RECT 2322.540 5.940 2322.740 6.140 ;
  LAYER VI3 ;
  RECT 2322.140 6.340 2322.340 6.540 ;
  LAYER VI3 ;
  RECT 2322.140 5.940 2322.340 6.140 ;
  LAYER VI3 ;
  RECT 2321.740 6.340 2321.940 6.540 ;
  LAYER VI3 ;
  RECT 2321.740 5.940 2321.940 6.140 ;
  LAYER VI3 ;
  RECT 2321.340 6.340 2321.540 6.540 ;
  LAYER VI3 ;
  RECT 2321.340 5.940 2321.540 6.140 ;
  LAYER VI3 ;
  RECT 2320.940 6.340 2321.140 6.540 ;
  LAYER VI3 ;
  RECT 2320.940 5.940 2321.140 6.140 ;
  LAYER VI3 ;
  RECT 2320.540 6.340 2320.740 6.540 ;
  LAYER VI3 ;
  RECT 2320.540 5.940 2320.740 6.140 ;
  LAYER VI3 ;
  RECT 2320.140 6.340 2320.340 6.540 ;
  LAYER VI3 ;
  RECT 2320.140 5.940 2320.340 6.140 ;
  LAYER VI3 ;
  RECT 2319.740 6.340 2319.940 6.540 ;
  LAYER VI3 ;
  RECT 2319.740 5.940 2319.940 6.140 ;
  LAYER VI3 ;
  RECT 2319.340 6.340 2319.540 6.540 ;
  LAYER VI3 ;
  RECT 2319.340 5.940 2319.540 6.140 ;
  LAYER VI3 ;
  RECT 2339.180 5.880 2347.180 6.740 ;
  LAYER VI3 ;
  RECT 2346.780 6.340 2346.980 6.540 ;
  LAYER VI3 ;
  RECT 2346.780 5.940 2346.980 6.140 ;
  LAYER VI3 ;
  RECT 2346.380 6.340 2346.580 6.540 ;
  LAYER VI3 ;
  RECT 2346.380 5.940 2346.580 6.140 ;
  LAYER VI3 ;
  RECT 2345.980 6.340 2346.180 6.540 ;
  LAYER VI3 ;
  RECT 2345.980 5.940 2346.180 6.140 ;
  LAYER VI3 ;
  RECT 2345.580 6.340 2345.780 6.540 ;
  LAYER VI3 ;
  RECT 2345.580 5.940 2345.780 6.140 ;
  LAYER VI3 ;
  RECT 2345.180 6.340 2345.380 6.540 ;
  LAYER VI3 ;
  RECT 2345.180 5.940 2345.380 6.140 ;
  LAYER VI3 ;
  RECT 2344.780 6.340 2344.980 6.540 ;
  LAYER VI3 ;
  RECT 2344.780 5.940 2344.980 6.140 ;
  LAYER VI3 ;
  RECT 2344.380 6.340 2344.580 6.540 ;
  LAYER VI3 ;
  RECT 2344.380 5.940 2344.580 6.140 ;
  LAYER VI3 ;
  RECT 2343.980 6.340 2344.180 6.540 ;
  LAYER VI3 ;
  RECT 2343.980 5.940 2344.180 6.140 ;
  LAYER VI3 ;
  RECT 2343.580 6.340 2343.780 6.540 ;
  LAYER VI3 ;
  RECT 2343.580 5.940 2343.780 6.140 ;
  LAYER VI3 ;
  RECT 2343.180 6.340 2343.380 6.540 ;
  LAYER VI3 ;
  RECT 2343.180 5.940 2343.380 6.140 ;
  LAYER VI3 ;
  RECT 2342.780 6.340 2342.980 6.540 ;
  LAYER VI3 ;
  RECT 2342.780 5.940 2342.980 6.140 ;
  LAYER VI3 ;
  RECT 2342.380 6.340 2342.580 6.540 ;
  LAYER VI3 ;
  RECT 2342.380 5.940 2342.580 6.140 ;
  LAYER VI3 ;
  RECT 2341.980 6.340 2342.180 6.540 ;
  LAYER VI3 ;
  RECT 2341.980 5.940 2342.180 6.140 ;
  LAYER VI3 ;
  RECT 2341.580 6.340 2341.780 6.540 ;
  LAYER VI3 ;
  RECT 2341.580 5.940 2341.780 6.140 ;
  LAYER VI3 ;
  RECT 2341.180 6.340 2341.380 6.540 ;
  LAYER VI3 ;
  RECT 2341.180 5.940 2341.380 6.140 ;
  LAYER VI3 ;
  RECT 2340.780 6.340 2340.980 6.540 ;
  LAYER VI3 ;
  RECT 2340.780 5.940 2340.980 6.140 ;
  LAYER VI3 ;
  RECT 2340.380 6.340 2340.580 6.540 ;
  LAYER VI3 ;
  RECT 2340.380 5.940 2340.580 6.140 ;
  LAYER VI3 ;
  RECT 2339.980 6.340 2340.180 6.540 ;
  LAYER VI3 ;
  RECT 2339.980 5.940 2340.180 6.140 ;
  LAYER VI3 ;
  RECT 2339.580 6.340 2339.780 6.540 ;
  LAYER VI3 ;
  RECT 2339.580 5.940 2339.780 6.140 ;
  LAYER VI3 ;
  RECT 2339.180 6.340 2339.380 6.540 ;
  LAYER VI3 ;
  RECT 2339.180 5.940 2339.380 6.140 ;
  LAYER VI3 ;
  RECT 2360.260 5.880 2368.260 6.740 ;
  LAYER VI3 ;
  RECT 2367.860 6.340 2368.060 6.540 ;
  LAYER VI3 ;
  RECT 2367.860 5.940 2368.060 6.140 ;
  LAYER VI3 ;
  RECT 2367.460 6.340 2367.660 6.540 ;
  LAYER VI3 ;
  RECT 2367.460 5.940 2367.660 6.140 ;
  LAYER VI3 ;
  RECT 2367.060 6.340 2367.260 6.540 ;
  LAYER VI3 ;
  RECT 2367.060 5.940 2367.260 6.140 ;
  LAYER VI3 ;
  RECT 2366.660 6.340 2366.860 6.540 ;
  LAYER VI3 ;
  RECT 2366.660 5.940 2366.860 6.140 ;
  LAYER VI3 ;
  RECT 2366.260 6.340 2366.460 6.540 ;
  LAYER VI3 ;
  RECT 2366.260 5.940 2366.460 6.140 ;
  LAYER VI3 ;
  RECT 2365.860 6.340 2366.060 6.540 ;
  LAYER VI3 ;
  RECT 2365.860 5.940 2366.060 6.140 ;
  LAYER VI3 ;
  RECT 2365.460 6.340 2365.660 6.540 ;
  LAYER VI3 ;
  RECT 2365.460 5.940 2365.660 6.140 ;
  LAYER VI3 ;
  RECT 2365.060 6.340 2365.260 6.540 ;
  LAYER VI3 ;
  RECT 2365.060 5.940 2365.260 6.140 ;
  LAYER VI3 ;
  RECT 2364.660 6.340 2364.860 6.540 ;
  LAYER VI3 ;
  RECT 2364.660 5.940 2364.860 6.140 ;
  LAYER VI3 ;
  RECT 2364.260 6.340 2364.460 6.540 ;
  LAYER VI3 ;
  RECT 2364.260 5.940 2364.460 6.140 ;
  LAYER VI3 ;
  RECT 2363.860 6.340 2364.060 6.540 ;
  LAYER VI3 ;
  RECT 2363.860 5.940 2364.060 6.140 ;
  LAYER VI3 ;
  RECT 2363.460 6.340 2363.660 6.540 ;
  LAYER VI3 ;
  RECT 2363.460 5.940 2363.660 6.140 ;
  LAYER VI3 ;
  RECT 2363.060 6.340 2363.260 6.540 ;
  LAYER VI3 ;
  RECT 2363.060 5.940 2363.260 6.140 ;
  LAYER VI3 ;
  RECT 2362.660 6.340 2362.860 6.540 ;
  LAYER VI3 ;
  RECT 2362.660 5.940 2362.860 6.140 ;
  LAYER VI3 ;
  RECT 2362.260 6.340 2362.460 6.540 ;
  LAYER VI3 ;
  RECT 2362.260 5.940 2362.460 6.140 ;
  LAYER VI3 ;
  RECT 2361.860 6.340 2362.060 6.540 ;
  LAYER VI3 ;
  RECT 2361.860 5.940 2362.060 6.140 ;
  LAYER VI3 ;
  RECT 2361.460 6.340 2361.660 6.540 ;
  LAYER VI3 ;
  RECT 2361.460 5.940 2361.660 6.140 ;
  LAYER VI3 ;
  RECT 2361.060 6.340 2361.260 6.540 ;
  LAYER VI3 ;
  RECT 2361.060 5.940 2361.260 6.140 ;
  LAYER VI3 ;
  RECT 2360.660 6.340 2360.860 6.540 ;
  LAYER VI3 ;
  RECT 2360.660 5.940 2360.860 6.140 ;
  LAYER VI3 ;
  RECT 2360.260 6.340 2360.460 6.540 ;
  LAYER VI3 ;
  RECT 2360.260 5.940 2360.460 6.140 ;
  LAYER VI3 ;
  RECT 2380.100 5.880 2388.100 6.740 ;
  LAYER VI3 ;
  RECT 2387.700 6.340 2387.900 6.540 ;
  LAYER VI3 ;
  RECT 2387.700 5.940 2387.900 6.140 ;
  LAYER VI3 ;
  RECT 2387.300 6.340 2387.500 6.540 ;
  LAYER VI3 ;
  RECT 2387.300 5.940 2387.500 6.140 ;
  LAYER VI3 ;
  RECT 2386.900 6.340 2387.100 6.540 ;
  LAYER VI3 ;
  RECT 2386.900 5.940 2387.100 6.140 ;
  LAYER VI3 ;
  RECT 2386.500 6.340 2386.700 6.540 ;
  LAYER VI3 ;
  RECT 2386.500 5.940 2386.700 6.140 ;
  LAYER VI3 ;
  RECT 2386.100 6.340 2386.300 6.540 ;
  LAYER VI3 ;
  RECT 2386.100 5.940 2386.300 6.140 ;
  LAYER VI3 ;
  RECT 2385.700 6.340 2385.900 6.540 ;
  LAYER VI3 ;
  RECT 2385.700 5.940 2385.900 6.140 ;
  LAYER VI3 ;
  RECT 2385.300 6.340 2385.500 6.540 ;
  LAYER VI3 ;
  RECT 2385.300 5.940 2385.500 6.140 ;
  LAYER VI3 ;
  RECT 2384.900 6.340 2385.100 6.540 ;
  LAYER VI3 ;
  RECT 2384.900 5.940 2385.100 6.140 ;
  LAYER VI3 ;
  RECT 2384.500 6.340 2384.700 6.540 ;
  LAYER VI3 ;
  RECT 2384.500 5.940 2384.700 6.140 ;
  LAYER VI3 ;
  RECT 2384.100 6.340 2384.300 6.540 ;
  LAYER VI3 ;
  RECT 2384.100 5.940 2384.300 6.140 ;
  LAYER VI3 ;
  RECT 2383.700 6.340 2383.900 6.540 ;
  LAYER VI3 ;
  RECT 2383.700 5.940 2383.900 6.140 ;
  LAYER VI3 ;
  RECT 2383.300 6.340 2383.500 6.540 ;
  LAYER VI3 ;
  RECT 2383.300 5.940 2383.500 6.140 ;
  LAYER VI3 ;
  RECT 2382.900 6.340 2383.100 6.540 ;
  LAYER VI3 ;
  RECT 2382.900 5.940 2383.100 6.140 ;
  LAYER VI3 ;
  RECT 2382.500 6.340 2382.700 6.540 ;
  LAYER VI3 ;
  RECT 2382.500 5.940 2382.700 6.140 ;
  LAYER VI3 ;
  RECT 2382.100 6.340 2382.300 6.540 ;
  LAYER VI3 ;
  RECT 2382.100 5.940 2382.300 6.140 ;
  LAYER VI3 ;
  RECT 2381.700 6.340 2381.900 6.540 ;
  LAYER VI3 ;
  RECT 2381.700 5.940 2381.900 6.140 ;
  LAYER VI3 ;
  RECT 2381.300 6.340 2381.500 6.540 ;
  LAYER VI3 ;
  RECT 2381.300 5.940 2381.500 6.140 ;
  LAYER VI3 ;
  RECT 2380.900 6.340 2381.100 6.540 ;
  LAYER VI3 ;
  RECT 2380.900 5.940 2381.100 6.140 ;
  LAYER VI3 ;
  RECT 2380.500 6.340 2380.700 6.540 ;
  LAYER VI3 ;
  RECT 2380.500 5.940 2380.700 6.140 ;
  LAYER VI3 ;
  RECT 2380.100 6.340 2380.300 6.540 ;
  LAYER VI3 ;
  RECT 2380.100 5.940 2380.300 6.140 ;
  LAYER VI3 ;
  RECT 2401.180 5.880 2409.180 6.740 ;
  LAYER VI3 ;
  RECT 2408.780 6.340 2408.980 6.540 ;
  LAYER VI3 ;
  RECT 2408.780 5.940 2408.980 6.140 ;
  LAYER VI3 ;
  RECT 2408.380 6.340 2408.580 6.540 ;
  LAYER VI3 ;
  RECT 2408.380 5.940 2408.580 6.140 ;
  LAYER VI3 ;
  RECT 2407.980 6.340 2408.180 6.540 ;
  LAYER VI3 ;
  RECT 2407.980 5.940 2408.180 6.140 ;
  LAYER VI3 ;
  RECT 2407.580 6.340 2407.780 6.540 ;
  LAYER VI3 ;
  RECT 2407.580 5.940 2407.780 6.140 ;
  LAYER VI3 ;
  RECT 2407.180 6.340 2407.380 6.540 ;
  LAYER VI3 ;
  RECT 2407.180 5.940 2407.380 6.140 ;
  LAYER VI3 ;
  RECT 2406.780 6.340 2406.980 6.540 ;
  LAYER VI3 ;
  RECT 2406.780 5.940 2406.980 6.140 ;
  LAYER VI3 ;
  RECT 2406.380 6.340 2406.580 6.540 ;
  LAYER VI3 ;
  RECT 2406.380 5.940 2406.580 6.140 ;
  LAYER VI3 ;
  RECT 2405.980 6.340 2406.180 6.540 ;
  LAYER VI3 ;
  RECT 2405.980 5.940 2406.180 6.140 ;
  LAYER VI3 ;
  RECT 2405.580 6.340 2405.780 6.540 ;
  LAYER VI3 ;
  RECT 2405.580 5.940 2405.780 6.140 ;
  LAYER VI3 ;
  RECT 2405.180 6.340 2405.380 6.540 ;
  LAYER VI3 ;
  RECT 2405.180 5.940 2405.380 6.140 ;
  LAYER VI3 ;
  RECT 2404.780 6.340 2404.980 6.540 ;
  LAYER VI3 ;
  RECT 2404.780 5.940 2404.980 6.140 ;
  LAYER VI3 ;
  RECT 2404.380 6.340 2404.580 6.540 ;
  LAYER VI3 ;
  RECT 2404.380 5.940 2404.580 6.140 ;
  LAYER VI3 ;
  RECT 2403.980 6.340 2404.180 6.540 ;
  LAYER VI3 ;
  RECT 2403.980 5.940 2404.180 6.140 ;
  LAYER VI3 ;
  RECT 2403.580 6.340 2403.780 6.540 ;
  LAYER VI3 ;
  RECT 2403.580 5.940 2403.780 6.140 ;
  LAYER VI3 ;
  RECT 2403.180 6.340 2403.380 6.540 ;
  LAYER VI3 ;
  RECT 2403.180 5.940 2403.380 6.140 ;
  LAYER VI3 ;
  RECT 2402.780 6.340 2402.980 6.540 ;
  LAYER VI3 ;
  RECT 2402.780 5.940 2402.980 6.140 ;
  LAYER VI3 ;
  RECT 2402.380 6.340 2402.580 6.540 ;
  LAYER VI3 ;
  RECT 2402.380 5.940 2402.580 6.140 ;
  LAYER VI3 ;
  RECT 2401.980 6.340 2402.180 6.540 ;
  LAYER VI3 ;
  RECT 2401.980 5.940 2402.180 6.140 ;
  LAYER VI3 ;
  RECT 2401.580 6.340 2401.780 6.540 ;
  LAYER VI3 ;
  RECT 2401.580 5.940 2401.780 6.140 ;
  LAYER VI3 ;
  RECT 2401.180 6.340 2401.380 6.540 ;
  LAYER VI3 ;
  RECT 2401.180 5.940 2401.380 6.140 ;
  LAYER VI3 ;
  RECT 2421.020 5.880 2429.020 6.740 ;
  LAYER VI3 ;
  RECT 2428.620 6.340 2428.820 6.540 ;
  LAYER VI3 ;
  RECT 2428.620 5.940 2428.820 6.140 ;
  LAYER VI3 ;
  RECT 2428.220 6.340 2428.420 6.540 ;
  LAYER VI3 ;
  RECT 2428.220 5.940 2428.420 6.140 ;
  LAYER VI3 ;
  RECT 2427.820 6.340 2428.020 6.540 ;
  LAYER VI3 ;
  RECT 2427.820 5.940 2428.020 6.140 ;
  LAYER VI3 ;
  RECT 2427.420 6.340 2427.620 6.540 ;
  LAYER VI3 ;
  RECT 2427.420 5.940 2427.620 6.140 ;
  LAYER VI3 ;
  RECT 2427.020 6.340 2427.220 6.540 ;
  LAYER VI3 ;
  RECT 2427.020 5.940 2427.220 6.140 ;
  LAYER VI3 ;
  RECT 2426.620 6.340 2426.820 6.540 ;
  LAYER VI3 ;
  RECT 2426.620 5.940 2426.820 6.140 ;
  LAYER VI3 ;
  RECT 2426.220 6.340 2426.420 6.540 ;
  LAYER VI3 ;
  RECT 2426.220 5.940 2426.420 6.140 ;
  LAYER VI3 ;
  RECT 2425.820 6.340 2426.020 6.540 ;
  LAYER VI3 ;
  RECT 2425.820 5.940 2426.020 6.140 ;
  LAYER VI3 ;
  RECT 2425.420 6.340 2425.620 6.540 ;
  LAYER VI3 ;
  RECT 2425.420 5.940 2425.620 6.140 ;
  LAYER VI3 ;
  RECT 2425.020 6.340 2425.220 6.540 ;
  LAYER VI3 ;
  RECT 2425.020 5.940 2425.220 6.140 ;
  LAYER VI3 ;
  RECT 2424.620 6.340 2424.820 6.540 ;
  LAYER VI3 ;
  RECT 2424.620 5.940 2424.820 6.140 ;
  LAYER VI3 ;
  RECT 2424.220 6.340 2424.420 6.540 ;
  LAYER VI3 ;
  RECT 2424.220 5.940 2424.420 6.140 ;
  LAYER VI3 ;
  RECT 2423.820 6.340 2424.020 6.540 ;
  LAYER VI3 ;
  RECT 2423.820 5.940 2424.020 6.140 ;
  LAYER VI3 ;
  RECT 2423.420 6.340 2423.620 6.540 ;
  LAYER VI3 ;
  RECT 2423.420 5.940 2423.620 6.140 ;
  LAYER VI3 ;
  RECT 2423.020 6.340 2423.220 6.540 ;
  LAYER VI3 ;
  RECT 2423.020 5.940 2423.220 6.140 ;
  LAYER VI3 ;
  RECT 2422.620 6.340 2422.820 6.540 ;
  LAYER VI3 ;
  RECT 2422.620 5.940 2422.820 6.140 ;
  LAYER VI3 ;
  RECT 2422.220 6.340 2422.420 6.540 ;
  LAYER VI3 ;
  RECT 2422.220 5.940 2422.420 6.140 ;
  LAYER VI3 ;
  RECT 2421.820 6.340 2422.020 6.540 ;
  LAYER VI3 ;
  RECT 2421.820 5.940 2422.020 6.140 ;
  LAYER VI3 ;
  RECT 2421.420 6.340 2421.620 6.540 ;
  LAYER VI3 ;
  RECT 2421.420 5.940 2421.620 6.140 ;
  LAYER VI3 ;
  RECT 2421.020 6.340 2421.220 6.540 ;
  LAYER VI3 ;
  RECT 2421.020 5.940 2421.220 6.140 ;
  LAYER VI3 ;
  RECT 2442.100 5.880 2450.100 6.740 ;
  LAYER VI3 ;
  RECT 2449.700 6.340 2449.900 6.540 ;
  LAYER VI3 ;
  RECT 2449.700 5.940 2449.900 6.140 ;
  LAYER VI3 ;
  RECT 2449.300 6.340 2449.500 6.540 ;
  LAYER VI3 ;
  RECT 2449.300 5.940 2449.500 6.140 ;
  LAYER VI3 ;
  RECT 2448.900 6.340 2449.100 6.540 ;
  LAYER VI3 ;
  RECT 2448.900 5.940 2449.100 6.140 ;
  LAYER VI3 ;
  RECT 2448.500 6.340 2448.700 6.540 ;
  LAYER VI3 ;
  RECT 2448.500 5.940 2448.700 6.140 ;
  LAYER VI3 ;
  RECT 2448.100 6.340 2448.300 6.540 ;
  LAYER VI3 ;
  RECT 2448.100 5.940 2448.300 6.140 ;
  LAYER VI3 ;
  RECT 2447.700 6.340 2447.900 6.540 ;
  LAYER VI3 ;
  RECT 2447.700 5.940 2447.900 6.140 ;
  LAYER VI3 ;
  RECT 2447.300 6.340 2447.500 6.540 ;
  LAYER VI3 ;
  RECT 2447.300 5.940 2447.500 6.140 ;
  LAYER VI3 ;
  RECT 2446.900 6.340 2447.100 6.540 ;
  LAYER VI3 ;
  RECT 2446.900 5.940 2447.100 6.140 ;
  LAYER VI3 ;
  RECT 2446.500 6.340 2446.700 6.540 ;
  LAYER VI3 ;
  RECT 2446.500 5.940 2446.700 6.140 ;
  LAYER VI3 ;
  RECT 2446.100 6.340 2446.300 6.540 ;
  LAYER VI3 ;
  RECT 2446.100 5.940 2446.300 6.140 ;
  LAYER VI3 ;
  RECT 2445.700 6.340 2445.900 6.540 ;
  LAYER VI3 ;
  RECT 2445.700 5.940 2445.900 6.140 ;
  LAYER VI3 ;
  RECT 2445.300 6.340 2445.500 6.540 ;
  LAYER VI3 ;
  RECT 2445.300 5.940 2445.500 6.140 ;
  LAYER VI3 ;
  RECT 2444.900 6.340 2445.100 6.540 ;
  LAYER VI3 ;
  RECT 2444.900 5.940 2445.100 6.140 ;
  LAYER VI3 ;
  RECT 2444.500 6.340 2444.700 6.540 ;
  LAYER VI3 ;
  RECT 2444.500 5.940 2444.700 6.140 ;
  LAYER VI3 ;
  RECT 2444.100 6.340 2444.300 6.540 ;
  LAYER VI3 ;
  RECT 2444.100 5.940 2444.300 6.140 ;
  LAYER VI3 ;
  RECT 2443.700 6.340 2443.900 6.540 ;
  LAYER VI3 ;
  RECT 2443.700 5.940 2443.900 6.140 ;
  LAYER VI3 ;
  RECT 2443.300 6.340 2443.500 6.540 ;
  LAYER VI3 ;
  RECT 2443.300 5.940 2443.500 6.140 ;
  LAYER VI3 ;
  RECT 2442.900 6.340 2443.100 6.540 ;
  LAYER VI3 ;
  RECT 2442.900 5.940 2443.100 6.140 ;
  LAYER VI3 ;
  RECT 2442.500 6.340 2442.700 6.540 ;
  LAYER VI3 ;
  RECT 2442.500 5.940 2442.700 6.140 ;
  LAYER VI3 ;
  RECT 2442.100 6.340 2442.300 6.540 ;
  LAYER VI3 ;
  RECT 2442.100 5.940 2442.300 6.140 ;
  LAYER VI3 ;
  RECT 2461.940 5.880 2469.940 6.740 ;
  LAYER VI3 ;
  RECT 2469.540 6.340 2469.740 6.540 ;
  LAYER VI3 ;
  RECT 2469.540 5.940 2469.740 6.140 ;
  LAYER VI3 ;
  RECT 2469.140 6.340 2469.340 6.540 ;
  LAYER VI3 ;
  RECT 2469.140 5.940 2469.340 6.140 ;
  LAYER VI3 ;
  RECT 2468.740 6.340 2468.940 6.540 ;
  LAYER VI3 ;
  RECT 2468.740 5.940 2468.940 6.140 ;
  LAYER VI3 ;
  RECT 2468.340 6.340 2468.540 6.540 ;
  LAYER VI3 ;
  RECT 2468.340 5.940 2468.540 6.140 ;
  LAYER VI3 ;
  RECT 2467.940 6.340 2468.140 6.540 ;
  LAYER VI3 ;
  RECT 2467.940 5.940 2468.140 6.140 ;
  LAYER VI3 ;
  RECT 2467.540 6.340 2467.740 6.540 ;
  LAYER VI3 ;
  RECT 2467.540 5.940 2467.740 6.140 ;
  LAYER VI3 ;
  RECT 2467.140 6.340 2467.340 6.540 ;
  LAYER VI3 ;
  RECT 2467.140 5.940 2467.340 6.140 ;
  LAYER VI3 ;
  RECT 2466.740 6.340 2466.940 6.540 ;
  LAYER VI3 ;
  RECT 2466.740 5.940 2466.940 6.140 ;
  LAYER VI3 ;
  RECT 2466.340 6.340 2466.540 6.540 ;
  LAYER VI3 ;
  RECT 2466.340 5.940 2466.540 6.140 ;
  LAYER VI3 ;
  RECT 2465.940 6.340 2466.140 6.540 ;
  LAYER VI3 ;
  RECT 2465.940 5.940 2466.140 6.140 ;
  LAYER VI3 ;
  RECT 2465.540 6.340 2465.740 6.540 ;
  LAYER VI3 ;
  RECT 2465.540 5.940 2465.740 6.140 ;
  LAYER VI3 ;
  RECT 2465.140 6.340 2465.340 6.540 ;
  LAYER VI3 ;
  RECT 2465.140 5.940 2465.340 6.140 ;
  LAYER VI3 ;
  RECT 2464.740 6.340 2464.940 6.540 ;
  LAYER VI3 ;
  RECT 2464.740 5.940 2464.940 6.140 ;
  LAYER VI3 ;
  RECT 2464.340 6.340 2464.540 6.540 ;
  LAYER VI3 ;
  RECT 2464.340 5.940 2464.540 6.140 ;
  LAYER VI3 ;
  RECT 2463.940 6.340 2464.140 6.540 ;
  LAYER VI3 ;
  RECT 2463.940 5.940 2464.140 6.140 ;
  LAYER VI3 ;
  RECT 2463.540 6.340 2463.740 6.540 ;
  LAYER VI3 ;
  RECT 2463.540 5.940 2463.740 6.140 ;
  LAYER VI3 ;
  RECT 2463.140 6.340 2463.340 6.540 ;
  LAYER VI3 ;
  RECT 2463.140 5.940 2463.340 6.140 ;
  LAYER VI3 ;
  RECT 2462.740 6.340 2462.940 6.540 ;
  LAYER VI3 ;
  RECT 2462.740 5.940 2462.940 6.140 ;
  LAYER VI3 ;
  RECT 2462.340 6.340 2462.540 6.540 ;
  LAYER VI3 ;
  RECT 2462.340 5.940 2462.540 6.140 ;
  LAYER VI3 ;
  RECT 2461.940 6.340 2462.140 6.540 ;
  LAYER VI3 ;
  RECT 2461.940 5.940 2462.140 6.140 ;
  LAYER VI3 ;
  RECT 2483.020 5.880 2491.020 6.740 ;
  LAYER VI3 ;
  RECT 2490.620 6.340 2490.820 6.540 ;
  LAYER VI3 ;
  RECT 2490.620 5.940 2490.820 6.140 ;
  LAYER VI3 ;
  RECT 2490.220 6.340 2490.420 6.540 ;
  LAYER VI3 ;
  RECT 2490.220 5.940 2490.420 6.140 ;
  LAYER VI3 ;
  RECT 2489.820 6.340 2490.020 6.540 ;
  LAYER VI3 ;
  RECT 2489.820 5.940 2490.020 6.140 ;
  LAYER VI3 ;
  RECT 2489.420 6.340 2489.620 6.540 ;
  LAYER VI3 ;
  RECT 2489.420 5.940 2489.620 6.140 ;
  LAYER VI3 ;
  RECT 2489.020 6.340 2489.220 6.540 ;
  LAYER VI3 ;
  RECT 2489.020 5.940 2489.220 6.140 ;
  LAYER VI3 ;
  RECT 2488.620 6.340 2488.820 6.540 ;
  LAYER VI3 ;
  RECT 2488.620 5.940 2488.820 6.140 ;
  LAYER VI3 ;
  RECT 2488.220 6.340 2488.420 6.540 ;
  LAYER VI3 ;
  RECT 2488.220 5.940 2488.420 6.140 ;
  LAYER VI3 ;
  RECT 2487.820 6.340 2488.020 6.540 ;
  LAYER VI3 ;
  RECT 2487.820 5.940 2488.020 6.140 ;
  LAYER VI3 ;
  RECT 2487.420 6.340 2487.620 6.540 ;
  LAYER VI3 ;
  RECT 2487.420 5.940 2487.620 6.140 ;
  LAYER VI3 ;
  RECT 2487.020 6.340 2487.220 6.540 ;
  LAYER VI3 ;
  RECT 2487.020 5.940 2487.220 6.140 ;
  LAYER VI3 ;
  RECT 2486.620 6.340 2486.820 6.540 ;
  LAYER VI3 ;
  RECT 2486.620 5.940 2486.820 6.140 ;
  LAYER VI3 ;
  RECT 2486.220 6.340 2486.420 6.540 ;
  LAYER VI3 ;
  RECT 2486.220 5.940 2486.420 6.140 ;
  LAYER VI3 ;
  RECT 2485.820 6.340 2486.020 6.540 ;
  LAYER VI3 ;
  RECT 2485.820 5.940 2486.020 6.140 ;
  LAYER VI3 ;
  RECT 2485.420 6.340 2485.620 6.540 ;
  LAYER VI3 ;
  RECT 2485.420 5.940 2485.620 6.140 ;
  LAYER VI3 ;
  RECT 2485.020 6.340 2485.220 6.540 ;
  LAYER VI3 ;
  RECT 2485.020 5.940 2485.220 6.140 ;
  LAYER VI3 ;
  RECT 2484.620 6.340 2484.820 6.540 ;
  LAYER VI3 ;
  RECT 2484.620 5.940 2484.820 6.140 ;
  LAYER VI3 ;
  RECT 2484.220 6.340 2484.420 6.540 ;
  LAYER VI3 ;
  RECT 2484.220 5.940 2484.420 6.140 ;
  LAYER VI3 ;
  RECT 2483.820 6.340 2484.020 6.540 ;
  LAYER VI3 ;
  RECT 2483.820 5.940 2484.020 6.140 ;
  LAYER VI3 ;
  RECT 2483.420 6.340 2483.620 6.540 ;
  LAYER VI3 ;
  RECT 2483.420 5.940 2483.620 6.140 ;
  LAYER VI3 ;
  RECT 2483.020 6.340 2483.220 6.540 ;
  LAYER VI3 ;
  RECT 2483.020 5.940 2483.220 6.140 ;
  LAYER VI3 ;
  RECT 2502.860 5.880 2510.860 6.740 ;
  LAYER VI3 ;
  RECT 2510.460 6.340 2510.660 6.540 ;
  LAYER VI3 ;
  RECT 2510.460 5.940 2510.660 6.140 ;
  LAYER VI3 ;
  RECT 2510.060 6.340 2510.260 6.540 ;
  LAYER VI3 ;
  RECT 2510.060 5.940 2510.260 6.140 ;
  LAYER VI3 ;
  RECT 2509.660 6.340 2509.860 6.540 ;
  LAYER VI3 ;
  RECT 2509.660 5.940 2509.860 6.140 ;
  LAYER VI3 ;
  RECT 2509.260 6.340 2509.460 6.540 ;
  LAYER VI3 ;
  RECT 2509.260 5.940 2509.460 6.140 ;
  LAYER VI3 ;
  RECT 2508.860 6.340 2509.060 6.540 ;
  LAYER VI3 ;
  RECT 2508.860 5.940 2509.060 6.140 ;
  LAYER VI3 ;
  RECT 2508.460 6.340 2508.660 6.540 ;
  LAYER VI3 ;
  RECT 2508.460 5.940 2508.660 6.140 ;
  LAYER VI3 ;
  RECT 2508.060 6.340 2508.260 6.540 ;
  LAYER VI3 ;
  RECT 2508.060 5.940 2508.260 6.140 ;
  LAYER VI3 ;
  RECT 2507.660 6.340 2507.860 6.540 ;
  LAYER VI3 ;
  RECT 2507.660 5.940 2507.860 6.140 ;
  LAYER VI3 ;
  RECT 2507.260 6.340 2507.460 6.540 ;
  LAYER VI3 ;
  RECT 2507.260 5.940 2507.460 6.140 ;
  LAYER VI3 ;
  RECT 2506.860 6.340 2507.060 6.540 ;
  LAYER VI3 ;
  RECT 2506.860 5.940 2507.060 6.140 ;
  LAYER VI3 ;
  RECT 2506.460 6.340 2506.660 6.540 ;
  LAYER VI3 ;
  RECT 2506.460 5.940 2506.660 6.140 ;
  LAYER VI3 ;
  RECT 2506.060 6.340 2506.260 6.540 ;
  LAYER VI3 ;
  RECT 2506.060 5.940 2506.260 6.140 ;
  LAYER VI3 ;
  RECT 2505.660 6.340 2505.860 6.540 ;
  LAYER VI3 ;
  RECT 2505.660 5.940 2505.860 6.140 ;
  LAYER VI3 ;
  RECT 2505.260 6.340 2505.460 6.540 ;
  LAYER VI3 ;
  RECT 2505.260 5.940 2505.460 6.140 ;
  LAYER VI3 ;
  RECT 2504.860 6.340 2505.060 6.540 ;
  LAYER VI3 ;
  RECT 2504.860 5.940 2505.060 6.140 ;
  LAYER VI3 ;
  RECT 2504.460 6.340 2504.660 6.540 ;
  LAYER VI3 ;
  RECT 2504.460 5.940 2504.660 6.140 ;
  LAYER VI3 ;
  RECT 2504.060 6.340 2504.260 6.540 ;
  LAYER VI3 ;
  RECT 2504.060 5.940 2504.260 6.140 ;
  LAYER VI3 ;
  RECT 2503.660 6.340 2503.860 6.540 ;
  LAYER VI3 ;
  RECT 2503.660 5.940 2503.860 6.140 ;
  LAYER VI3 ;
  RECT 2503.260 6.340 2503.460 6.540 ;
  LAYER VI3 ;
  RECT 2503.260 5.940 2503.460 6.140 ;
  LAYER VI3 ;
  RECT 2502.860 6.340 2503.060 6.540 ;
  LAYER VI3 ;
  RECT 2502.860 5.940 2503.060 6.140 ;
  LAYER VI3 ;
  RECT 2523.940 5.880 2531.940 6.740 ;
  LAYER VI3 ;
  RECT 2531.540 6.340 2531.740 6.540 ;
  LAYER VI3 ;
  RECT 2531.540 5.940 2531.740 6.140 ;
  LAYER VI3 ;
  RECT 2531.140 6.340 2531.340 6.540 ;
  LAYER VI3 ;
  RECT 2531.140 5.940 2531.340 6.140 ;
  LAYER VI3 ;
  RECT 2530.740 6.340 2530.940 6.540 ;
  LAYER VI3 ;
  RECT 2530.740 5.940 2530.940 6.140 ;
  LAYER VI3 ;
  RECT 2530.340 6.340 2530.540 6.540 ;
  LAYER VI3 ;
  RECT 2530.340 5.940 2530.540 6.140 ;
  LAYER VI3 ;
  RECT 2529.940 6.340 2530.140 6.540 ;
  LAYER VI3 ;
  RECT 2529.940 5.940 2530.140 6.140 ;
  LAYER VI3 ;
  RECT 2529.540 6.340 2529.740 6.540 ;
  LAYER VI3 ;
  RECT 2529.540 5.940 2529.740 6.140 ;
  LAYER VI3 ;
  RECT 2529.140 6.340 2529.340 6.540 ;
  LAYER VI3 ;
  RECT 2529.140 5.940 2529.340 6.140 ;
  LAYER VI3 ;
  RECT 2528.740 6.340 2528.940 6.540 ;
  LAYER VI3 ;
  RECT 2528.740 5.940 2528.940 6.140 ;
  LAYER VI3 ;
  RECT 2528.340 6.340 2528.540 6.540 ;
  LAYER VI3 ;
  RECT 2528.340 5.940 2528.540 6.140 ;
  LAYER VI3 ;
  RECT 2527.940 6.340 2528.140 6.540 ;
  LAYER VI3 ;
  RECT 2527.940 5.940 2528.140 6.140 ;
  LAYER VI3 ;
  RECT 2527.540 6.340 2527.740 6.540 ;
  LAYER VI3 ;
  RECT 2527.540 5.940 2527.740 6.140 ;
  LAYER VI3 ;
  RECT 2527.140 6.340 2527.340 6.540 ;
  LAYER VI3 ;
  RECT 2527.140 5.940 2527.340 6.140 ;
  LAYER VI3 ;
  RECT 2526.740 6.340 2526.940 6.540 ;
  LAYER VI3 ;
  RECT 2526.740 5.940 2526.940 6.140 ;
  LAYER VI3 ;
  RECT 2526.340 6.340 2526.540 6.540 ;
  LAYER VI3 ;
  RECT 2526.340 5.940 2526.540 6.140 ;
  LAYER VI3 ;
  RECT 2525.940 6.340 2526.140 6.540 ;
  LAYER VI3 ;
  RECT 2525.940 5.940 2526.140 6.140 ;
  LAYER VI3 ;
  RECT 2525.540 6.340 2525.740 6.540 ;
  LAYER VI3 ;
  RECT 2525.540 5.940 2525.740 6.140 ;
  LAYER VI3 ;
  RECT 2525.140 6.340 2525.340 6.540 ;
  LAYER VI3 ;
  RECT 2525.140 5.940 2525.340 6.140 ;
  LAYER VI3 ;
  RECT 2524.740 6.340 2524.940 6.540 ;
  LAYER VI3 ;
  RECT 2524.740 5.940 2524.940 6.140 ;
  LAYER VI3 ;
  RECT 2524.340 6.340 2524.540 6.540 ;
  LAYER VI3 ;
  RECT 2524.340 5.940 2524.540 6.140 ;
  LAYER VI3 ;
  RECT 2523.940 6.340 2524.140 6.540 ;
  LAYER VI3 ;
  RECT 2523.940 5.940 2524.140 6.140 ;
  LAYER VI3 ;
  RECT 2543.780 5.880 2551.780 6.740 ;
  LAYER VI3 ;
  RECT 2551.380 6.340 2551.580 6.540 ;
  LAYER VI3 ;
  RECT 2551.380 5.940 2551.580 6.140 ;
  LAYER VI3 ;
  RECT 2550.980 6.340 2551.180 6.540 ;
  LAYER VI3 ;
  RECT 2550.980 5.940 2551.180 6.140 ;
  LAYER VI3 ;
  RECT 2550.580 6.340 2550.780 6.540 ;
  LAYER VI3 ;
  RECT 2550.580 5.940 2550.780 6.140 ;
  LAYER VI3 ;
  RECT 2550.180 6.340 2550.380 6.540 ;
  LAYER VI3 ;
  RECT 2550.180 5.940 2550.380 6.140 ;
  LAYER VI3 ;
  RECT 2549.780 6.340 2549.980 6.540 ;
  LAYER VI3 ;
  RECT 2549.780 5.940 2549.980 6.140 ;
  LAYER VI3 ;
  RECT 2549.380 6.340 2549.580 6.540 ;
  LAYER VI3 ;
  RECT 2549.380 5.940 2549.580 6.140 ;
  LAYER VI3 ;
  RECT 2548.980 6.340 2549.180 6.540 ;
  LAYER VI3 ;
  RECT 2548.980 5.940 2549.180 6.140 ;
  LAYER VI3 ;
  RECT 2548.580 6.340 2548.780 6.540 ;
  LAYER VI3 ;
  RECT 2548.580 5.940 2548.780 6.140 ;
  LAYER VI3 ;
  RECT 2548.180 6.340 2548.380 6.540 ;
  LAYER VI3 ;
  RECT 2548.180 5.940 2548.380 6.140 ;
  LAYER VI3 ;
  RECT 2547.780 6.340 2547.980 6.540 ;
  LAYER VI3 ;
  RECT 2547.780 5.940 2547.980 6.140 ;
  LAYER VI3 ;
  RECT 2547.380 6.340 2547.580 6.540 ;
  LAYER VI3 ;
  RECT 2547.380 5.940 2547.580 6.140 ;
  LAYER VI3 ;
  RECT 2546.980 6.340 2547.180 6.540 ;
  LAYER VI3 ;
  RECT 2546.980 5.940 2547.180 6.140 ;
  LAYER VI3 ;
  RECT 2546.580 6.340 2546.780 6.540 ;
  LAYER VI3 ;
  RECT 2546.580 5.940 2546.780 6.140 ;
  LAYER VI3 ;
  RECT 2546.180 6.340 2546.380 6.540 ;
  LAYER VI3 ;
  RECT 2546.180 5.940 2546.380 6.140 ;
  LAYER VI3 ;
  RECT 2545.780 6.340 2545.980 6.540 ;
  LAYER VI3 ;
  RECT 2545.780 5.940 2545.980 6.140 ;
  LAYER VI3 ;
  RECT 2545.380 6.340 2545.580 6.540 ;
  LAYER VI3 ;
  RECT 2545.380 5.940 2545.580 6.140 ;
  LAYER VI3 ;
  RECT 2544.980 6.340 2545.180 6.540 ;
  LAYER VI3 ;
  RECT 2544.980 5.940 2545.180 6.140 ;
  LAYER VI3 ;
  RECT 2544.580 6.340 2544.780 6.540 ;
  LAYER VI3 ;
  RECT 2544.580 5.940 2544.780 6.140 ;
  LAYER VI3 ;
  RECT 2544.180 6.340 2544.380 6.540 ;
  LAYER VI3 ;
  RECT 2544.180 5.940 2544.380 6.140 ;
  LAYER VI3 ;
  RECT 2543.780 6.340 2543.980 6.540 ;
  LAYER VI3 ;
  RECT 2543.780 5.940 2543.980 6.140 ;
  LAYER VI3 ;
  RECT 2564.860 5.880 2572.860 6.740 ;
  LAYER VI3 ;
  RECT 2572.460 6.340 2572.660 6.540 ;
  LAYER VI3 ;
  RECT 2572.460 5.940 2572.660 6.140 ;
  LAYER VI3 ;
  RECT 2572.060 6.340 2572.260 6.540 ;
  LAYER VI3 ;
  RECT 2572.060 5.940 2572.260 6.140 ;
  LAYER VI3 ;
  RECT 2571.660 6.340 2571.860 6.540 ;
  LAYER VI3 ;
  RECT 2571.660 5.940 2571.860 6.140 ;
  LAYER VI3 ;
  RECT 2571.260 6.340 2571.460 6.540 ;
  LAYER VI3 ;
  RECT 2571.260 5.940 2571.460 6.140 ;
  LAYER VI3 ;
  RECT 2570.860 6.340 2571.060 6.540 ;
  LAYER VI3 ;
  RECT 2570.860 5.940 2571.060 6.140 ;
  LAYER VI3 ;
  RECT 2570.460 6.340 2570.660 6.540 ;
  LAYER VI3 ;
  RECT 2570.460 5.940 2570.660 6.140 ;
  LAYER VI3 ;
  RECT 2570.060 6.340 2570.260 6.540 ;
  LAYER VI3 ;
  RECT 2570.060 5.940 2570.260 6.140 ;
  LAYER VI3 ;
  RECT 2569.660 6.340 2569.860 6.540 ;
  LAYER VI3 ;
  RECT 2569.660 5.940 2569.860 6.140 ;
  LAYER VI3 ;
  RECT 2569.260 6.340 2569.460 6.540 ;
  LAYER VI3 ;
  RECT 2569.260 5.940 2569.460 6.140 ;
  LAYER VI3 ;
  RECT 2568.860 6.340 2569.060 6.540 ;
  LAYER VI3 ;
  RECT 2568.860 5.940 2569.060 6.140 ;
  LAYER VI3 ;
  RECT 2568.460 6.340 2568.660 6.540 ;
  LAYER VI3 ;
  RECT 2568.460 5.940 2568.660 6.140 ;
  LAYER VI3 ;
  RECT 2568.060 6.340 2568.260 6.540 ;
  LAYER VI3 ;
  RECT 2568.060 5.940 2568.260 6.140 ;
  LAYER VI3 ;
  RECT 2567.660 6.340 2567.860 6.540 ;
  LAYER VI3 ;
  RECT 2567.660 5.940 2567.860 6.140 ;
  LAYER VI3 ;
  RECT 2567.260 6.340 2567.460 6.540 ;
  LAYER VI3 ;
  RECT 2567.260 5.940 2567.460 6.140 ;
  LAYER VI3 ;
  RECT 2566.860 6.340 2567.060 6.540 ;
  LAYER VI3 ;
  RECT 2566.860 5.940 2567.060 6.140 ;
  LAYER VI3 ;
  RECT 2566.460 6.340 2566.660 6.540 ;
  LAYER VI3 ;
  RECT 2566.460 5.940 2566.660 6.140 ;
  LAYER VI3 ;
  RECT 2566.060 6.340 2566.260 6.540 ;
  LAYER VI3 ;
  RECT 2566.060 5.940 2566.260 6.140 ;
  LAYER VI3 ;
  RECT 2565.660 6.340 2565.860 6.540 ;
  LAYER VI3 ;
  RECT 2565.660 5.940 2565.860 6.140 ;
  LAYER VI3 ;
  RECT 2565.260 6.340 2565.460 6.540 ;
  LAYER VI3 ;
  RECT 2565.260 5.940 2565.460 6.140 ;
  LAYER VI3 ;
  RECT 2564.860 6.340 2565.060 6.540 ;
  LAYER VI3 ;
  RECT 2564.860 5.940 2565.060 6.140 ;
  LAYER VI3 ;
  RECT 2584.700 5.880 2592.700 6.740 ;
  LAYER VI3 ;
  RECT 2592.300 6.340 2592.500 6.540 ;
  LAYER VI3 ;
  RECT 2592.300 5.940 2592.500 6.140 ;
  LAYER VI3 ;
  RECT 2591.900 6.340 2592.100 6.540 ;
  LAYER VI3 ;
  RECT 2591.900 5.940 2592.100 6.140 ;
  LAYER VI3 ;
  RECT 2591.500 6.340 2591.700 6.540 ;
  LAYER VI3 ;
  RECT 2591.500 5.940 2591.700 6.140 ;
  LAYER VI3 ;
  RECT 2591.100 6.340 2591.300 6.540 ;
  LAYER VI3 ;
  RECT 2591.100 5.940 2591.300 6.140 ;
  LAYER VI3 ;
  RECT 2590.700 6.340 2590.900 6.540 ;
  LAYER VI3 ;
  RECT 2590.700 5.940 2590.900 6.140 ;
  LAYER VI3 ;
  RECT 2590.300 6.340 2590.500 6.540 ;
  LAYER VI3 ;
  RECT 2590.300 5.940 2590.500 6.140 ;
  LAYER VI3 ;
  RECT 2589.900 6.340 2590.100 6.540 ;
  LAYER VI3 ;
  RECT 2589.900 5.940 2590.100 6.140 ;
  LAYER VI3 ;
  RECT 2589.500 6.340 2589.700 6.540 ;
  LAYER VI3 ;
  RECT 2589.500 5.940 2589.700 6.140 ;
  LAYER VI3 ;
  RECT 2589.100 6.340 2589.300 6.540 ;
  LAYER VI3 ;
  RECT 2589.100 5.940 2589.300 6.140 ;
  LAYER VI3 ;
  RECT 2588.700 6.340 2588.900 6.540 ;
  LAYER VI3 ;
  RECT 2588.700 5.940 2588.900 6.140 ;
  LAYER VI3 ;
  RECT 2588.300 6.340 2588.500 6.540 ;
  LAYER VI3 ;
  RECT 2588.300 5.940 2588.500 6.140 ;
  LAYER VI3 ;
  RECT 2587.900 6.340 2588.100 6.540 ;
  LAYER VI3 ;
  RECT 2587.900 5.940 2588.100 6.140 ;
  LAYER VI3 ;
  RECT 2587.500 6.340 2587.700 6.540 ;
  LAYER VI3 ;
  RECT 2587.500 5.940 2587.700 6.140 ;
  LAYER VI3 ;
  RECT 2587.100 6.340 2587.300 6.540 ;
  LAYER VI3 ;
  RECT 2587.100 5.940 2587.300 6.140 ;
  LAYER VI3 ;
  RECT 2586.700 6.340 2586.900 6.540 ;
  LAYER VI3 ;
  RECT 2586.700 5.940 2586.900 6.140 ;
  LAYER VI3 ;
  RECT 2586.300 6.340 2586.500 6.540 ;
  LAYER VI3 ;
  RECT 2586.300 5.940 2586.500 6.140 ;
  LAYER VI3 ;
  RECT 2585.900 6.340 2586.100 6.540 ;
  LAYER VI3 ;
  RECT 2585.900 5.940 2586.100 6.140 ;
  LAYER VI3 ;
  RECT 2585.500 6.340 2585.700 6.540 ;
  LAYER VI3 ;
  RECT 2585.500 5.940 2585.700 6.140 ;
  LAYER VI3 ;
  RECT 2585.100 6.340 2585.300 6.540 ;
  LAYER VI3 ;
  RECT 2585.100 5.940 2585.300 6.140 ;
  LAYER VI3 ;
  RECT 2584.700 6.340 2584.900 6.540 ;
  LAYER VI3 ;
  RECT 2584.700 5.940 2584.900 6.140 ;
  LAYER VI3 ;
  RECT 2605.780 5.880 2613.780 6.740 ;
  LAYER VI3 ;
  RECT 2613.380 6.340 2613.580 6.540 ;
  LAYER VI3 ;
  RECT 2613.380 5.940 2613.580 6.140 ;
  LAYER VI3 ;
  RECT 2612.980 6.340 2613.180 6.540 ;
  LAYER VI3 ;
  RECT 2612.980 5.940 2613.180 6.140 ;
  LAYER VI3 ;
  RECT 2612.580 6.340 2612.780 6.540 ;
  LAYER VI3 ;
  RECT 2612.580 5.940 2612.780 6.140 ;
  LAYER VI3 ;
  RECT 2612.180 6.340 2612.380 6.540 ;
  LAYER VI3 ;
  RECT 2612.180 5.940 2612.380 6.140 ;
  LAYER VI3 ;
  RECT 2611.780 6.340 2611.980 6.540 ;
  LAYER VI3 ;
  RECT 2611.780 5.940 2611.980 6.140 ;
  LAYER VI3 ;
  RECT 2611.380 6.340 2611.580 6.540 ;
  LAYER VI3 ;
  RECT 2611.380 5.940 2611.580 6.140 ;
  LAYER VI3 ;
  RECT 2610.980 6.340 2611.180 6.540 ;
  LAYER VI3 ;
  RECT 2610.980 5.940 2611.180 6.140 ;
  LAYER VI3 ;
  RECT 2610.580 6.340 2610.780 6.540 ;
  LAYER VI3 ;
  RECT 2610.580 5.940 2610.780 6.140 ;
  LAYER VI3 ;
  RECT 2610.180 6.340 2610.380 6.540 ;
  LAYER VI3 ;
  RECT 2610.180 5.940 2610.380 6.140 ;
  LAYER VI3 ;
  RECT 2609.780 6.340 2609.980 6.540 ;
  LAYER VI3 ;
  RECT 2609.780 5.940 2609.980 6.140 ;
  LAYER VI3 ;
  RECT 2609.380 6.340 2609.580 6.540 ;
  LAYER VI3 ;
  RECT 2609.380 5.940 2609.580 6.140 ;
  LAYER VI3 ;
  RECT 2608.980 6.340 2609.180 6.540 ;
  LAYER VI3 ;
  RECT 2608.980 5.940 2609.180 6.140 ;
  LAYER VI3 ;
  RECT 2608.580 6.340 2608.780 6.540 ;
  LAYER VI3 ;
  RECT 2608.580 5.940 2608.780 6.140 ;
  LAYER VI3 ;
  RECT 2608.180 6.340 2608.380 6.540 ;
  LAYER VI3 ;
  RECT 2608.180 5.940 2608.380 6.140 ;
  LAYER VI3 ;
  RECT 2607.780 6.340 2607.980 6.540 ;
  LAYER VI3 ;
  RECT 2607.780 5.940 2607.980 6.140 ;
  LAYER VI3 ;
  RECT 2607.380 6.340 2607.580 6.540 ;
  LAYER VI3 ;
  RECT 2607.380 5.940 2607.580 6.140 ;
  LAYER VI3 ;
  RECT 2606.980 6.340 2607.180 6.540 ;
  LAYER VI3 ;
  RECT 2606.980 5.940 2607.180 6.140 ;
  LAYER VI3 ;
  RECT 2606.580 6.340 2606.780 6.540 ;
  LAYER VI3 ;
  RECT 2606.580 5.940 2606.780 6.140 ;
  LAYER VI3 ;
  RECT 2606.180 6.340 2606.380 6.540 ;
  LAYER VI3 ;
  RECT 2606.180 5.940 2606.380 6.140 ;
  LAYER VI3 ;
  RECT 2605.780 6.340 2605.980 6.540 ;
  LAYER VI3 ;
  RECT 2605.780 5.940 2605.980 6.140 ;
  LAYER VI3 ;
  RECT 2625.620 5.880 2633.620 6.740 ;
  LAYER VI3 ;
  RECT 2633.220 6.340 2633.420 6.540 ;
  LAYER VI3 ;
  RECT 2633.220 5.940 2633.420 6.140 ;
  LAYER VI3 ;
  RECT 2632.820 6.340 2633.020 6.540 ;
  LAYER VI3 ;
  RECT 2632.820 5.940 2633.020 6.140 ;
  LAYER VI3 ;
  RECT 2632.420 6.340 2632.620 6.540 ;
  LAYER VI3 ;
  RECT 2632.420 5.940 2632.620 6.140 ;
  LAYER VI3 ;
  RECT 2632.020 6.340 2632.220 6.540 ;
  LAYER VI3 ;
  RECT 2632.020 5.940 2632.220 6.140 ;
  LAYER VI3 ;
  RECT 2631.620 6.340 2631.820 6.540 ;
  LAYER VI3 ;
  RECT 2631.620 5.940 2631.820 6.140 ;
  LAYER VI3 ;
  RECT 2631.220 6.340 2631.420 6.540 ;
  LAYER VI3 ;
  RECT 2631.220 5.940 2631.420 6.140 ;
  LAYER VI3 ;
  RECT 2630.820 6.340 2631.020 6.540 ;
  LAYER VI3 ;
  RECT 2630.820 5.940 2631.020 6.140 ;
  LAYER VI3 ;
  RECT 2630.420 6.340 2630.620 6.540 ;
  LAYER VI3 ;
  RECT 2630.420 5.940 2630.620 6.140 ;
  LAYER VI3 ;
  RECT 2630.020 6.340 2630.220 6.540 ;
  LAYER VI3 ;
  RECT 2630.020 5.940 2630.220 6.140 ;
  LAYER VI3 ;
  RECT 2629.620 6.340 2629.820 6.540 ;
  LAYER VI3 ;
  RECT 2629.620 5.940 2629.820 6.140 ;
  LAYER VI3 ;
  RECT 2629.220 6.340 2629.420 6.540 ;
  LAYER VI3 ;
  RECT 2629.220 5.940 2629.420 6.140 ;
  LAYER VI3 ;
  RECT 2628.820 6.340 2629.020 6.540 ;
  LAYER VI3 ;
  RECT 2628.820 5.940 2629.020 6.140 ;
  LAYER VI3 ;
  RECT 2628.420 6.340 2628.620 6.540 ;
  LAYER VI3 ;
  RECT 2628.420 5.940 2628.620 6.140 ;
  LAYER VI3 ;
  RECT 2628.020 6.340 2628.220 6.540 ;
  LAYER VI3 ;
  RECT 2628.020 5.940 2628.220 6.140 ;
  LAYER VI3 ;
  RECT 2627.620 6.340 2627.820 6.540 ;
  LAYER VI3 ;
  RECT 2627.620 5.940 2627.820 6.140 ;
  LAYER VI3 ;
  RECT 2627.220 6.340 2627.420 6.540 ;
  LAYER VI3 ;
  RECT 2627.220 5.940 2627.420 6.140 ;
  LAYER VI3 ;
  RECT 2626.820 6.340 2627.020 6.540 ;
  LAYER VI3 ;
  RECT 2626.820 5.940 2627.020 6.140 ;
  LAYER VI3 ;
  RECT 2626.420 6.340 2626.620 6.540 ;
  LAYER VI3 ;
  RECT 2626.420 5.940 2626.620 6.140 ;
  LAYER VI3 ;
  RECT 2626.020 6.340 2626.220 6.540 ;
  LAYER VI3 ;
  RECT 2626.020 5.940 2626.220 6.140 ;
  LAYER VI3 ;
  RECT 2625.620 6.340 2625.820 6.540 ;
  LAYER VI3 ;
  RECT 2625.620 5.940 2625.820 6.140 ;
  LAYER VI3 ;
  RECT 2646.700 5.880 2654.700 6.740 ;
  LAYER VI3 ;
  RECT 2654.300 6.340 2654.500 6.540 ;
  LAYER VI3 ;
  RECT 2654.300 5.940 2654.500 6.140 ;
  LAYER VI3 ;
  RECT 2653.900 6.340 2654.100 6.540 ;
  LAYER VI3 ;
  RECT 2653.900 5.940 2654.100 6.140 ;
  LAYER VI3 ;
  RECT 2653.500 6.340 2653.700 6.540 ;
  LAYER VI3 ;
  RECT 2653.500 5.940 2653.700 6.140 ;
  LAYER VI3 ;
  RECT 2653.100 6.340 2653.300 6.540 ;
  LAYER VI3 ;
  RECT 2653.100 5.940 2653.300 6.140 ;
  LAYER VI3 ;
  RECT 2652.700 6.340 2652.900 6.540 ;
  LAYER VI3 ;
  RECT 2652.700 5.940 2652.900 6.140 ;
  LAYER VI3 ;
  RECT 2652.300 6.340 2652.500 6.540 ;
  LAYER VI3 ;
  RECT 2652.300 5.940 2652.500 6.140 ;
  LAYER VI3 ;
  RECT 2651.900 6.340 2652.100 6.540 ;
  LAYER VI3 ;
  RECT 2651.900 5.940 2652.100 6.140 ;
  LAYER VI3 ;
  RECT 2651.500 6.340 2651.700 6.540 ;
  LAYER VI3 ;
  RECT 2651.500 5.940 2651.700 6.140 ;
  LAYER VI3 ;
  RECT 2651.100 6.340 2651.300 6.540 ;
  LAYER VI3 ;
  RECT 2651.100 5.940 2651.300 6.140 ;
  LAYER VI3 ;
  RECT 2650.700 6.340 2650.900 6.540 ;
  LAYER VI3 ;
  RECT 2650.700 5.940 2650.900 6.140 ;
  LAYER VI3 ;
  RECT 2650.300 6.340 2650.500 6.540 ;
  LAYER VI3 ;
  RECT 2650.300 5.940 2650.500 6.140 ;
  LAYER VI3 ;
  RECT 2649.900 6.340 2650.100 6.540 ;
  LAYER VI3 ;
  RECT 2649.900 5.940 2650.100 6.140 ;
  LAYER VI3 ;
  RECT 2649.500 6.340 2649.700 6.540 ;
  LAYER VI3 ;
  RECT 2649.500 5.940 2649.700 6.140 ;
  LAYER VI3 ;
  RECT 2649.100 6.340 2649.300 6.540 ;
  LAYER VI3 ;
  RECT 2649.100 5.940 2649.300 6.140 ;
  LAYER VI3 ;
  RECT 2648.700 6.340 2648.900 6.540 ;
  LAYER VI3 ;
  RECT 2648.700 5.940 2648.900 6.140 ;
  LAYER VI3 ;
  RECT 2648.300 6.340 2648.500 6.540 ;
  LAYER VI3 ;
  RECT 2648.300 5.940 2648.500 6.140 ;
  LAYER VI3 ;
  RECT 2647.900 6.340 2648.100 6.540 ;
  LAYER VI3 ;
  RECT 2647.900 5.940 2648.100 6.140 ;
  LAYER VI3 ;
  RECT 2647.500 6.340 2647.700 6.540 ;
  LAYER VI3 ;
  RECT 2647.500 5.940 2647.700 6.140 ;
  LAYER VI3 ;
  RECT 2647.100 6.340 2647.300 6.540 ;
  LAYER VI3 ;
  RECT 2647.100 5.940 2647.300 6.140 ;
  LAYER VI3 ;
  RECT 2646.700 6.340 2646.900 6.540 ;
  LAYER VI3 ;
  RECT 2646.700 5.940 2646.900 6.140 ;
  LAYER VI3 ;
  RECT 2666.540 5.880 2674.540 6.740 ;
  LAYER VI3 ;
  RECT 2674.140 6.340 2674.340 6.540 ;
  LAYER VI3 ;
  RECT 2674.140 5.940 2674.340 6.140 ;
  LAYER VI3 ;
  RECT 2673.740 6.340 2673.940 6.540 ;
  LAYER VI3 ;
  RECT 2673.740 5.940 2673.940 6.140 ;
  LAYER VI3 ;
  RECT 2673.340 6.340 2673.540 6.540 ;
  LAYER VI3 ;
  RECT 2673.340 5.940 2673.540 6.140 ;
  LAYER VI3 ;
  RECT 2672.940 6.340 2673.140 6.540 ;
  LAYER VI3 ;
  RECT 2672.940 5.940 2673.140 6.140 ;
  LAYER VI3 ;
  RECT 2672.540 6.340 2672.740 6.540 ;
  LAYER VI3 ;
  RECT 2672.540 5.940 2672.740 6.140 ;
  LAYER VI3 ;
  RECT 2672.140 6.340 2672.340 6.540 ;
  LAYER VI3 ;
  RECT 2672.140 5.940 2672.340 6.140 ;
  LAYER VI3 ;
  RECT 2671.740 6.340 2671.940 6.540 ;
  LAYER VI3 ;
  RECT 2671.740 5.940 2671.940 6.140 ;
  LAYER VI3 ;
  RECT 2671.340 6.340 2671.540 6.540 ;
  LAYER VI3 ;
  RECT 2671.340 5.940 2671.540 6.140 ;
  LAYER VI3 ;
  RECT 2670.940 6.340 2671.140 6.540 ;
  LAYER VI3 ;
  RECT 2670.940 5.940 2671.140 6.140 ;
  LAYER VI3 ;
  RECT 2670.540 6.340 2670.740 6.540 ;
  LAYER VI3 ;
  RECT 2670.540 5.940 2670.740 6.140 ;
  LAYER VI3 ;
  RECT 2670.140 6.340 2670.340 6.540 ;
  LAYER VI3 ;
  RECT 2670.140 5.940 2670.340 6.140 ;
  LAYER VI3 ;
  RECT 2669.740 6.340 2669.940 6.540 ;
  LAYER VI3 ;
  RECT 2669.740 5.940 2669.940 6.140 ;
  LAYER VI3 ;
  RECT 2669.340 6.340 2669.540 6.540 ;
  LAYER VI3 ;
  RECT 2669.340 5.940 2669.540 6.140 ;
  LAYER VI3 ;
  RECT 2668.940 6.340 2669.140 6.540 ;
  LAYER VI3 ;
  RECT 2668.940 5.940 2669.140 6.140 ;
  LAYER VI3 ;
  RECT 2668.540 6.340 2668.740 6.540 ;
  LAYER VI3 ;
  RECT 2668.540 5.940 2668.740 6.140 ;
  LAYER VI3 ;
  RECT 2668.140 6.340 2668.340 6.540 ;
  LAYER VI3 ;
  RECT 2668.140 5.940 2668.340 6.140 ;
  LAYER VI3 ;
  RECT 2667.740 6.340 2667.940 6.540 ;
  LAYER VI3 ;
  RECT 2667.740 5.940 2667.940 6.140 ;
  LAYER VI3 ;
  RECT 2667.340 6.340 2667.540 6.540 ;
  LAYER VI3 ;
  RECT 2667.340 5.940 2667.540 6.140 ;
  LAYER VI3 ;
  RECT 2666.940 6.340 2667.140 6.540 ;
  LAYER VI3 ;
  RECT 2666.940 5.940 2667.140 6.140 ;
  LAYER VI3 ;
  RECT 2666.540 6.340 2666.740 6.540 ;
  LAYER VI3 ;
  RECT 2666.540 5.940 2666.740 6.140 ;
  LAYER VI3 ;
  RECT 1343.440 5.880 1346.890 6.740 ;
  LAYER VI3 ;
  RECT 1346.640 6.340 1346.840 6.540 ;
  LAYER VI3 ;
  RECT 1346.640 5.940 1346.840 6.140 ;
  LAYER VI3 ;
  RECT 1346.240 6.340 1346.440 6.540 ;
  LAYER VI3 ;
  RECT 1346.240 5.940 1346.440 6.140 ;
  LAYER VI3 ;
  RECT 1345.840 6.340 1346.040 6.540 ;
  LAYER VI3 ;
  RECT 1345.840 5.940 1346.040 6.140 ;
  LAYER VI3 ;
  RECT 1345.440 6.340 1345.640 6.540 ;
  LAYER VI3 ;
  RECT 1345.440 5.940 1345.640 6.140 ;
  LAYER VI3 ;
  RECT 1345.040 6.340 1345.240 6.540 ;
  LAYER VI3 ;
  RECT 1345.040 5.940 1345.240 6.140 ;
  LAYER VI3 ;
  RECT 1344.640 6.340 1344.840 6.540 ;
  LAYER VI3 ;
  RECT 1344.640 5.940 1344.840 6.140 ;
  LAYER VI3 ;
  RECT 1344.240 6.340 1344.440 6.540 ;
  LAYER VI3 ;
  RECT 1344.240 5.940 1344.440 6.140 ;
  LAYER VI3 ;
  RECT 1343.840 6.340 1344.040 6.540 ;
  LAYER VI3 ;
  RECT 1343.840 5.940 1344.040 6.140 ;
  LAYER VI3 ;
  RECT 1343.440 6.340 1343.640 6.540 ;
  LAYER VI3 ;
  RECT 1343.440 5.940 1343.640 6.140 ;
  LAYER VI3 ;
  RECT 1352.290 5.880 1358.210 6.740 ;
  LAYER VI3 ;
  RECT 1357.890 6.340 1358.090 6.540 ;
  LAYER VI3 ;
  RECT 1357.890 5.940 1358.090 6.140 ;
  LAYER VI3 ;
  RECT 1357.490 6.340 1357.690 6.540 ;
  LAYER VI3 ;
  RECT 1357.490 5.940 1357.690 6.140 ;
  LAYER VI3 ;
  RECT 1357.090 6.340 1357.290 6.540 ;
  LAYER VI3 ;
  RECT 1357.090 5.940 1357.290 6.140 ;
  LAYER VI3 ;
  RECT 1356.690 6.340 1356.890 6.540 ;
  LAYER VI3 ;
  RECT 1356.690 5.940 1356.890 6.140 ;
  LAYER VI3 ;
  RECT 1356.290 6.340 1356.490 6.540 ;
  LAYER VI3 ;
  RECT 1356.290 5.940 1356.490 6.140 ;
  LAYER VI3 ;
  RECT 1355.890 6.340 1356.090 6.540 ;
  LAYER VI3 ;
  RECT 1355.890 5.940 1356.090 6.140 ;
  LAYER VI3 ;
  RECT 1355.490 6.340 1355.690 6.540 ;
  LAYER VI3 ;
  RECT 1355.490 5.940 1355.690 6.140 ;
  LAYER VI3 ;
  RECT 1355.090 6.340 1355.290 6.540 ;
  LAYER VI3 ;
  RECT 1355.090 5.940 1355.290 6.140 ;
  LAYER VI3 ;
  RECT 1354.690 6.340 1354.890 6.540 ;
  LAYER VI3 ;
  RECT 1354.690 5.940 1354.890 6.140 ;
  LAYER VI3 ;
  RECT 1354.290 6.340 1354.490 6.540 ;
  LAYER VI3 ;
  RECT 1354.290 5.940 1354.490 6.140 ;
  LAYER VI3 ;
  RECT 1353.890 6.340 1354.090 6.540 ;
  LAYER VI3 ;
  RECT 1353.890 5.940 1354.090 6.140 ;
  LAYER VI3 ;
  RECT 1353.490 6.340 1353.690 6.540 ;
  LAYER VI3 ;
  RECT 1353.490 5.940 1353.690 6.140 ;
  LAYER VI3 ;
  RECT 1353.090 6.340 1353.290 6.540 ;
  LAYER VI3 ;
  RECT 1353.090 5.940 1353.290 6.140 ;
  LAYER VI3 ;
  RECT 1352.690 6.340 1352.890 6.540 ;
  LAYER VI3 ;
  RECT 1352.690 5.940 1352.890 6.140 ;
  LAYER VI3 ;
  RECT 1352.290 6.340 1352.490 6.540 ;
  LAYER VI3 ;
  RECT 1352.290 5.940 1352.490 6.140 ;
  LAYER VI3 ;
  RECT 1335.160 5.880 1336.920 6.740 ;
  LAYER VI3 ;
  RECT 1336.360 6.340 1336.560 6.540 ;
  LAYER VI3 ;
  RECT 1336.360 5.940 1336.560 6.140 ;
  LAYER VI3 ;
  RECT 1335.960 6.340 1336.160 6.540 ;
  LAYER VI3 ;
  RECT 1335.960 5.940 1336.160 6.140 ;
  LAYER VI3 ;
  RECT 1335.560 6.340 1335.760 6.540 ;
  LAYER VI3 ;
  RECT 1335.560 5.940 1335.760 6.140 ;
  LAYER VI3 ;
  RECT 1335.160 6.340 1335.360 6.540 ;
  LAYER VI3 ;
  RECT 1335.160 5.940 1335.360 6.140 ;
  LAYER VI3 ;
  RECT 1329.820 5.880 1331.580 6.740 ;
  LAYER VI3 ;
  RECT 1331.020 6.340 1331.220 6.540 ;
  LAYER VI3 ;
  RECT 1331.020 5.940 1331.220 6.140 ;
  LAYER VI3 ;
  RECT 1330.620 6.340 1330.820 6.540 ;
  LAYER VI3 ;
  RECT 1330.620 5.940 1330.820 6.140 ;
  LAYER VI3 ;
  RECT 1330.220 6.340 1330.420 6.540 ;
  LAYER VI3 ;
  RECT 1330.220 5.940 1330.420 6.140 ;
  LAYER VI3 ;
  RECT 1329.820 6.340 1330.020 6.540 ;
  LAYER VI3 ;
  RECT 1329.820 5.940 1330.020 6.140 ;
  LAYER VI3 ;
  RECT 1325.820 5.880 1327.580 6.740 ;
  LAYER VI3 ;
  RECT 1327.020 6.340 1327.220 6.540 ;
  LAYER VI3 ;
  RECT 1327.020 5.940 1327.220 6.140 ;
  LAYER VI3 ;
  RECT 1326.620 6.340 1326.820 6.540 ;
  LAYER VI3 ;
  RECT 1326.620 5.940 1326.820 6.140 ;
  LAYER VI3 ;
  RECT 1326.220 6.340 1326.420 6.540 ;
  LAYER VI3 ;
  RECT 1326.220 5.940 1326.420 6.140 ;
  LAYER VI3 ;
  RECT 1325.820 6.340 1326.020 6.540 ;
  LAYER VI3 ;
  RECT 1325.820 5.940 1326.020 6.140 ;
  LAYER VI3 ;
  RECT 1321.820 5.880 1323.580 6.740 ;
  LAYER VI3 ;
  RECT 1323.020 6.340 1323.220 6.540 ;
  LAYER VI3 ;
  RECT 1323.020 5.940 1323.220 6.140 ;
  LAYER VI3 ;
  RECT 1322.620 6.340 1322.820 6.540 ;
  LAYER VI3 ;
  RECT 1322.620 5.940 1322.820 6.140 ;
  LAYER VI3 ;
  RECT 1322.220 6.340 1322.420 6.540 ;
  LAYER VI3 ;
  RECT 1322.220 5.940 1322.420 6.140 ;
  LAYER VI3 ;
  RECT 1321.820 6.340 1322.020 6.540 ;
  LAYER VI3 ;
  RECT 1321.820 5.940 1322.020 6.140 ;
  LAYER VI3 ;
  RECT 1317.820 5.880 1319.580 6.740 ;
  LAYER VI3 ;
  RECT 1319.020 6.340 1319.220 6.540 ;
  LAYER VI3 ;
  RECT 1319.020 5.940 1319.220 6.140 ;
  LAYER VI3 ;
  RECT 1318.620 6.340 1318.820 6.540 ;
  LAYER VI3 ;
  RECT 1318.620 5.940 1318.820 6.140 ;
  LAYER VI3 ;
  RECT 1318.220 6.340 1318.420 6.540 ;
  LAYER VI3 ;
  RECT 1318.220 5.940 1318.420 6.140 ;
  LAYER VI3 ;
  RECT 1317.820 6.340 1318.020 6.540 ;
  LAYER VI3 ;
  RECT 1317.820 5.940 1318.020 6.140 ;
  LAYER VI3 ;
  RECT 4.280 57.100 5.140 61.420 ;
  LAYER VI3 ;
  RECT 4.740 61.100 4.940 61.300 ;
  LAYER VI3 ;
  RECT 4.740 60.700 4.940 60.900 ;
  LAYER VI3 ;
  RECT 4.740 60.300 4.940 60.500 ;
  LAYER VI3 ;
  RECT 4.740 59.900 4.940 60.100 ;
  LAYER VI3 ;
  RECT 4.740 59.500 4.940 59.700 ;
  LAYER VI3 ;
  RECT 4.740 59.100 4.940 59.300 ;
  LAYER VI3 ;
  RECT 4.740 58.700 4.940 58.900 ;
  LAYER VI3 ;
  RECT 4.740 58.300 4.940 58.500 ;
  LAYER VI3 ;
  RECT 4.740 57.900 4.940 58.100 ;
  LAYER VI3 ;
  RECT 4.740 57.500 4.940 57.700 ;
  LAYER VI3 ;
  RECT 4.740 57.100 4.940 57.300 ;
  LAYER VI3 ;
  RECT 4.340 61.100 4.540 61.300 ;
  LAYER VI3 ;
  RECT 4.340 60.700 4.540 60.900 ;
  LAYER VI3 ;
  RECT 4.340 60.300 4.540 60.500 ;
  LAYER VI3 ;
  RECT 4.340 59.900 4.540 60.100 ;
  LAYER VI3 ;
  RECT 4.340 59.500 4.540 59.700 ;
  LAYER VI3 ;
  RECT 4.340 59.100 4.540 59.300 ;
  LAYER VI3 ;
  RECT 4.340 58.700 4.540 58.900 ;
  LAYER VI3 ;
  RECT 4.340 58.300 4.540 58.500 ;
  LAYER VI3 ;
  RECT 4.340 57.900 4.540 58.100 ;
  LAYER VI3 ;
  RECT 4.340 57.500 4.540 57.700 ;
  LAYER VI3 ;
  RECT 4.340 57.100 4.540 57.300 ;
  LAYER VI2 ;
  RECT 4.280 57.100 5.140 61.420 ;
  LAYER VI2 ;
  RECT 4.740 61.100 4.940 61.300 ;
  LAYER VI2 ;
  RECT 4.740 60.700 4.940 60.900 ;
  LAYER VI2 ;
  RECT 4.740 60.300 4.940 60.500 ;
  LAYER VI2 ;
  RECT 4.740 59.900 4.940 60.100 ;
  LAYER VI2 ;
  RECT 4.740 59.500 4.940 59.700 ;
  LAYER VI2 ;
  RECT 4.740 59.100 4.940 59.300 ;
  LAYER VI2 ;
  RECT 4.740 58.700 4.940 58.900 ;
  LAYER VI2 ;
  RECT 4.740 58.300 4.940 58.500 ;
  LAYER VI2 ;
  RECT 4.740 57.900 4.940 58.100 ;
  LAYER VI2 ;
  RECT 4.740 57.500 4.940 57.700 ;
  LAYER VI2 ;
  RECT 4.740 57.100 4.940 57.300 ;
  LAYER VI2 ;
  RECT 4.340 61.100 4.540 61.300 ;
  LAYER VI2 ;
  RECT 4.340 60.700 4.540 60.900 ;
  LAYER VI2 ;
  RECT 4.340 60.300 4.540 60.500 ;
  LAYER VI2 ;
  RECT 4.340 59.900 4.540 60.100 ;
  LAYER VI2 ;
  RECT 4.340 59.500 4.540 59.700 ;
  LAYER VI2 ;
  RECT 4.340 59.100 4.540 59.300 ;
  LAYER VI2 ;
  RECT 4.340 58.700 4.540 58.900 ;
  LAYER VI2 ;
  RECT 4.340 58.300 4.540 58.500 ;
  LAYER VI2 ;
  RECT 4.340 57.900 4.540 58.100 ;
  LAYER VI2 ;
  RECT 4.340 57.500 4.540 57.700 ;
  LAYER VI2 ;
  RECT 4.340 57.100 4.540 57.300 ;
  LAYER VI3 ;
  RECT 4.280 45.560 5.140 46.160 ;
  LAYER VI3 ;
  RECT 4.680 45.620 4.880 45.820 ;
  LAYER VI3 ;
  RECT 4.280 45.620 4.480 45.820 ;
  LAYER VI2 ;
  RECT 4.280 45.560 5.140 46.160 ;
  LAYER VI2 ;
  RECT 4.680 45.620 4.880 45.820 ;
  LAYER VI2 ;
  RECT 4.280 45.620 4.480 45.820 ;
  LAYER VI3 ;
  RECT 4.280 39.480 5.140 40.080 ;
  LAYER VI3 ;
  RECT 4.680 39.540 4.880 39.740 ;
  LAYER VI3 ;
  RECT 4.280 39.540 4.480 39.740 ;
  LAYER VI2 ;
  RECT 4.280 39.480 5.140 40.080 ;
  LAYER VI2 ;
  RECT 4.680 39.540 4.880 39.740 ;
  LAYER VI2 ;
  RECT 4.280 39.540 4.480 39.740 ;
  LAYER VI3 ;
  RECT 4.280 36.320 5.140 37.320 ;
  LAYER VI3 ;
  RECT 4.740 36.720 4.940 36.920 ;
  LAYER VI3 ;
  RECT 4.740 36.320 4.940 36.520 ;
  LAYER VI3 ;
  RECT 4.340 36.720 4.540 36.920 ;
  LAYER VI3 ;
  RECT 4.340 36.320 4.540 36.520 ;
  LAYER VI2 ;
  RECT 4.280 36.320 5.140 37.320 ;
  LAYER VI2 ;
  RECT 4.740 36.720 4.940 36.920 ;
  LAYER VI2 ;
  RECT 4.740 36.320 4.940 36.520 ;
  LAYER VI2 ;
  RECT 4.340 36.720 4.540 36.920 ;
  LAYER VI2 ;
  RECT 4.340 36.320 4.540 36.520 ;
  LAYER VI3 ;
  RECT 4.280 24.170 5.140 25.170 ;
  LAYER VI3 ;
  RECT 4.740 24.570 4.940 24.770 ;
  LAYER VI3 ;
  RECT 4.740 24.170 4.940 24.370 ;
  LAYER VI3 ;
  RECT 4.340 24.570 4.540 24.770 ;
  LAYER VI3 ;
  RECT 4.340 24.170 4.540 24.370 ;
  LAYER VI2 ;
  RECT 4.280 24.170 5.140 25.170 ;
  LAYER VI2 ;
  RECT 4.740 24.570 4.940 24.770 ;
  LAYER VI2 ;
  RECT 4.740 24.170 4.940 24.370 ;
  LAYER VI2 ;
  RECT 4.340 24.570 4.540 24.770 ;
  LAYER VI2 ;
  RECT 4.340 24.170 4.540 24.370 ;
  LAYER VI3 ;
  RECT 4.280 21.230 5.140 22.070 ;
  LAYER VI3 ;
  RECT 4.680 21.690 4.880 21.890 ;
  LAYER VI3 ;
  RECT 4.680 21.290 4.880 21.490 ;
  LAYER VI3 ;
  RECT 4.280 21.690 4.480 21.890 ;
  LAYER VI3 ;
  RECT 4.280 21.290 4.480 21.490 ;
  LAYER VI2 ;
  RECT 4.280 21.230 5.140 22.070 ;
  LAYER VI2 ;
  RECT 4.680 21.690 4.880 21.890 ;
  LAYER VI2 ;
  RECT 4.680 21.290 4.880 21.490 ;
  LAYER VI2 ;
  RECT 4.280 21.690 4.480 21.890 ;
  LAYER VI2 ;
  RECT 4.280 21.290 4.480 21.490 ;
  LAYER VI3 ;
  RECT 4.280 18.730 5.140 19.730 ;
  LAYER VI3 ;
  RECT 4.740 19.130 4.940 19.330 ;
  LAYER VI3 ;
  RECT 4.740 18.730 4.940 18.930 ;
  LAYER VI3 ;
  RECT 4.340 19.130 4.540 19.330 ;
  LAYER VI3 ;
  RECT 4.340 18.730 4.540 18.930 ;
  LAYER VI2 ;
  RECT 4.280 18.730 5.140 19.730 ;
  LAYER VI2 ;
  RECT 4.740 19.130 4.940 19.330 ;
  LAYER VI2 ;
  RECT 4.740 18.730 4.940 18.930 ;
  LAYER VI2 ;
  RECT 4.340 19.130 4.540 19.330 ;
  LAYER VI2 ;
  RECT 4.340 18.730 4.540 18.930 ;
  LAYER VI3 ;
  RECT 4.280 14.200 5.140 15.200 ;
  LAYER VI3 ;
  RECT 4.740 14.600 4.940 14.800 ;
  LAYER VI3 ;
  RECT 4.740 14.200 4.940 14.400 ;
  LAYER VI3 ;
  RECT 4.340 14.600 4.540 14.800 ;
  LAYER VI3 ;
  RECT 4.340 14.200 4.540 14.400 ;
  LAYER VI2 ;
  RECT 4.280 14.200 5.140 15.200 ;
  LAYER VI2 ;
  RECT 4.740 14.600 4.940 14.800 ;
  LAYER VI2 ;
  RECT 4.740 14.200 4.940 14.400 ;
  LAYER VI2 ;
  RECT 4.340 14.600 4.540 14.800 ;
  LAYER VI2 ;
  RECT 4.340 14.200 4.540 14.400 ;
  LAYER VI3 ;
  RECT 4.280 9.570 5.140 11.170 ;
  LAYER VI3 ;
  RECT 4.740 10.770 4.940 10.970 ;
  LAYER VI3 ;
  RECT 4.740 10.370 4.940 10.570 ;
  LAYER VI3 ;
  RECT 4.740 9.970 4.940 10.170 ;
  LAYER VI3 ;
  RECT 4.740 9.570 4.940 9.770 ;
  LAYER VI3 ;
  RECT 4.340 10.770 4.540 10.970 ;
  LAYER VI3 ;
  RECT 4.340 10.370 4.540 10.570 ;
  LAYER VI3 ;
  RECT 4.340 9.970 4.540 10.170 ;
  LAYER VI3 ;
  RECT 4.340 9.570 4.540 9.770 ;
  LAYER VI2 ;
  RECT 4.280 9.570 5.140 11.170 ;
  LAYER VI2 ;
  RECT 4.740 10.770 4.940 10.970 ;
  LAYER VI2 ;
  RECT 4.740 10.370 4.940 10.570 ;
  LAYER VI2 ;
  RECT 4.740 9.970 4.940 10.170 ;
  LAYER VI2 ;
  RECT 4.740 9.570 4.940 9.770 ;
  LAYER VI2 ;
  RECT 4.340 10.770 4.540 10.970 ;
  LAYER VI2 ;
  RECT 4.340 10.370 4.540 10.570 ;
  LAYER VI2 ;
  RECT 4.340 9.970 4.540 10.170 ;
  LAYER VI2 ;
  RECT 4.340 9.570 4.540 9.770 ;
  LAYER VI3 ;
  RECT 5.420 5.880 6.560 6.740 ;
  LAYER VI3 ;
  RECT 6.220 6.340 6.420 6.540 ;
  LAYER VI3 ;
  RECT 6.220 5.940 6.420 6.140 ;
  LAYER VI3 ;
  RECT 5.820 6.340 6.020 6.540 ;
  LAYER VI3 ;
  RECT 5.820 5.940 6.020 6.140 ;
  LAYER VI3 ;
  RECT 5.420 6.340 5.620 6.540 ;
  LAYER VI3 ;
  RECT 5.420 5.940 5.620 6.140 ;
  LAYER VI3 ;
  RECT 8.360 5.880 16.360 6.740 ;
  LAYER VI3 ;
  RECT 15.960 6.340 16.160 6.540 ;
  LAYER VI3 ;
  RECT 15.960 5.940 16.160 6.140 ;
  LAYER VI3 ;
  RECT 15.560 6.340 15.760 6.540 ;
  LAYER VI3 ;
  RECT 15.560 5.940 15.760 6.140 ;
  LAYER VI3 ;
  RECT 15.160 6.340 15.360 6.540 ;
  LAYER VI3 ;
  RECT 15.160 5.940 15.360 6.140 ;
  LAYER VI3 ;
  RECT 14.760 6.340 14.960 6.540 ;
  LAYER VI3 ;
  RECT 14.760 5.940 14.960 6.140 ;
  LAYER VI3 ;
  RECT 14.360 6.340 14.560 6.540 ;
  LAYER VI3 ;
  RECT 14.360 5.940 14.560 6.140 ;
  LAYER VI3 ;
  RECT 13.960 6.340 14.160 6.540 ;
  LAYER VI3 ;
  RECT 13.960 5.940 14.160 6.140 ;
  LAYER VI3 ;
  RECT 13.560 6.340 13.760 6.540 ;
  LAYER VI3 ;
  RECT 13.560 5.940 13.760 6.140 ;
  LAYER VI3 ;
  RECT 13.160 6.340 13.360 6.540 ;
  LAYER VI3 ;
  RECT 13.160 5.940 13.360 6.140 ;
  LAYER VI3 ;
  RECT 12.760 6.340 12.960 6.540 ;
  LAYER VI3 ;
  RECT 12.760 5.940 12.960 6.140 ;
  LAYER VI3 ;
  RECT 12.360 6.340 12.560 6.540 ;
  LAYER VI3 ;
  RECT 12.360 5.940 12.560 6.140 ;
  LAYER VI3 ;
  RECT 11.960 6.340 12.160 6.540 ;
  LAYER VI3 ;
  RECT 11.960 5.940 12.160 6.140 ;
  LAYER VI3 ;
  RECT 11.560 6.340 11.760 6.540 ;
  LAYER VI3 ;
  RECT 11.560 5.940 11.760 6.140 ;
  LAYER VI3 ;
  RECT 11.160 6.340 11.360 6.540 ;
  LAYER VI3 ;
  RECT 11.160 5.940 11.360 6.140 ;
  LAYER VI3 ;
  RECT 10.760 6.340 10.960 6.540 ;
  LAYER VI3 ;
  RECT 10.760 5.940 10.960 6.140 ;
  LAYER VI3 ;
  RECT 10.360 6.340 10.560 6.540 ;
  LAYER VI3 ;
  RECT 10.360 5.940 10.560 6.140 ;
  LAYER VI3 ;
  RECT 9.960 6.340 10.160 6.540 ;
  LAYER VI3 ;
  RECT 9.960 5.940 10.160 6.140 ;
  LAYER VI3 ;
  RECT 9.560 6.340 9.760 6.540 ;
  LAYER VI3 ;
  RECT 9.560 5.940 9.760 6.140 ;
  LAYER VI3 ;
  RECT 9.160 6.340 9.360 6.540 ;
  LAYER VI3 ;
  RECT 9.160 5.940 9.360 6.140 ;
  LAYER VI3 ;
  RECT 8.760 6.340 8.960 6.540 ;
  LAYER VI3 ;
  RECT 8.760 5.940 8.960 6.140 ;
  LAYER VI3 ;
  RECT 8.360 6.340 8.560 6.540 ;
  LAYER VI3 ;
  RECT 8.360 5.940 8.560 6.140 ;
  LAYER VI3 ;
  RECT 28.200 5.880 36.200 6.740 ;
  LAYER VI3 ;
  RECT 35.800 6.340 36.000 6.540 ;
  LAYER VI3 ;
  RECT 35.800 5.940 36.000 6.140 ;
  LAYER VI3 ;
  RECT 35.400 6.340 35.600 6.540 ;
  LAYER VI3 ;
  RECT 35.400 5.940 35.600 6.140 ;
  LAYER VI3 ;
  RECT 35.000 6.340 35.200 6.540 ;
  LAYER VI3 ;
  RECT 35.000 5.940 35.200 6.140 ;
  LAYER VI3 ;
  RECT 34.600 6.340 34.800 6.540 ;
  LAYER VI3 ;
  RECT 34.600 5.940 34.800 6.140 ;
  LAYER VI3 ;
  RECT 34.200 6.340 34.400 6.540 ;
  LAYER VI3 ;
  RECT 34.200 5.940 34.400 6.140 ;
  LAYER VI3 ;
  RECT 33.800 6.340 34.000 6.540 ;
  LAYER VI3 ;
  RECT 33.800 5.940 34.000 6.140 ;
  LAYER VI3 ;
  RECT 33.400 6.340 33.600 6.540 ;
  LAYER VI3 ;
  RECT 33.400 5.940 33.600 6.140 ;
  LAYER VI3 ;
  RECT 33.000 6.340 33.200 6.540 ;
  LAYER VI3 ;
  RECT 33.000 5.940 33.200 6.140 ;
  LAYER VI3 ;
  RECT 32.600 6.340 32.800 6.540 ;
  LAYER VI3 ;
  RECT 32.600 5.940 32.800 6.140 ;
  LAYER VI3 ;
  RECT 32.200 6.340 32.400 6.540 ;
  LAYER VI3 ;
  RECT 32.200 5.940 32.400 6.140 ;
  LAYER VI3 ;
  RECT 31.800 6.340 32.000 6.540 ;
  LAYER VI3 ;
  RECT 31.800 5.940 32.000 6.140 ;
  LAYER VI3 ;
  RECT 31.400 6.340 31.600 6.540 ;
  LAYER VI3 ;
  RECT 31.400 5.940 31.600 6.140 ;
  LAYER VI3 ;
  RECT 31.000 6.340 31.200 6.540 ;
  LAYER VI3 ;
  RECT 31.000 5.940 31.200 6.140 ;
  LAYER VI3 ;
  RECT 30.600 6.340 30.800 6.540 ;
  LAYER VI3 ;
  RECT 30.600 5.940 30.800 6.140 ;
  LAYER VI3 ;
  RECT 30.200 6.340 30.400 6.540 ;
  LAYER VI3 ;
  RECT 30.200 5.940 30.400 6.140 ;
  LAYER VI3 ;
  RECT 29.800 6.340 30.000 6.540 ;
  LAYER VI3 ;
  RECT 29.800 5.940 30.000 6.140 ;
  LAYER VI3 ;
  RECT 29.400 6.340 29.600 6.540 ;
  LAYER VI3 ;
  RECT 29.400 5.940 29.600 6.140 ;
  LAYER VI3 ;
  RECT 29.000 6.340 29.200 6.540 ;
  LAYER VI3 ;
  RECT 29.000 5.940 29.200 6.140 ;
  LAYER VI3 ;
  RECT 28.600 6.340 28.800 6.540 ;
  LAYER VI3 ;
  RECT 28.600 5.940 28.800 6.140 ;
  LAYER VI3 ;
  RECT 28.200 6.340 28.400 6.540 ;
  LAYER VI3 ;
  RECT 28.200 5.940 28.400 6.140 ;
  LAYER VI3 ;
  RECT 49.280 5.880 57.280 6.740 ;
  LAYER VI3 ;
  RECT 56.880 6.340 57.080 6.540 ;
  LAYER VI3 ;
  RECT 56.880 5.940 57.080 6.140 ;
  LAYER VI3 ;
  RECT 56.480 6.340 56.680 6.540 ;
  LAYER VI3 ;
  RECT 56.480 5.940 56.680 6.140 ;
  LAYER VI3 ;
  RECT 56.080 6.340 56.280 6.540 ;
  LAYER VI3 ;
  RECT 56.080 5.940 56.280 6.140 ;
  LAYER VI3 ;
  RECT 55.680 6.340 55.880 6.540 ;
  LAYER VI3 ;
  RECT 55.680 5.940 55.880 6.140 ;
  LAYER VI3 ;
  RECT 55.280 6.340 55.480 6.540 ;
  LAYER VI3 ;
  RECT 55.280 5.940 55.480 6.140 ;
  LAYER VI3 ;
  RECT 54.880 6.340 55.080 6.540 ;
  LAYER VI3 ;
  RECT 54.880 5.940 55.080 6.140 ;
  LAYER VI3 ;
  RECT 54.480 6.340 54.680 6.540 ;
  LAYER VI3 ;
  RECT 54.480 5.940 54.680 6.140 ;
  LAYER VI3 ;
  RECT 54.080 6.340 54.280 6.540 ;
  LAYER VI3 ;
  RECT 54.080 5.940 54.280 6.140 ;
  LAYER VI3 ;
  RECT 53.680 6.340 53.880 6.540 ;
  LAYER VI3 ;
  RECT 53.680 5.940 53.880 6.140 ;
  LAYER VI3 ;
  RECT 53.280 6.340 53.480 6.540 ;
  LAYER VI3 ;
  RECT 53.280 5.940 53.480 6.140 ;
  LAYER VI3 ;
  RECT 52.880 6.340 53.080 6.540 ;
  LAYER VI3 ;
  RECT 52.880 5.940 53.080 6.140 ;
  LAYER VI3 ;
  RECT 52.480 6.340 52.680 6.540 ;
  LAYER VI3 ;
  RECT 52.480 5.940 52.680 6.140 ;
  LAYER VI3 ;
  RECT 52.080 6.340 52.280 6.540 ;
  LAYER VI3 ;
  RECT 52.080 5.940 52.280 6.140 ;
  LAYER VI3 ;
  RECT 51.680 6.340 51.880 6.540 ;
  LAYER VI3 ;
  RECT 51.680 5.940 51.880 6.140 ;
  LAYER VI3 ;
  RECT 51.280 6.340 51.480 6.540 ;
  LAYER VI3 ;
  RECT 51.280 5.940 51.480 6.140 ;
  LAYER VI3 ;
  RECT 50.880 6.340 51.080 6.540 ;
  LAYER VI3 ;
  RECT 50.880 5.940 51.080 6.140 ;
  LAYER VI3 ;
  RECT 50.480 6.340 50.680 6.540 ;
  LAYER VI3 ;
  RECT 50.480 5.940 50.680 6.140 ;
  LAYER VI3 ;
  RECT 50.080 6.340 50.280 6.540 ;
  LAYER VI3 ;
  RECT 50.080 5.940 50.280 6.140 ;
  LAYER VI3 ;
  RECT 49.680 6.340 49.880 6.540 ;
  LAYER VI3 ;
  RECT 49.680 5.940 49.880 6.140 ;
  LAYER VI3 ;
  RECT 49.280 6.340 49.480 6.540 ;
  LAYER VI3 ;
  RECT 49.280 5.940 49.480 6.140 ;
  LAYER VI3 ;
  RECT 69.120 5.880 77.120 6.740 ;
  LAYER VI3 ;
  RECT 76.720 6.340 76.920 6.540 ;
  LAYER VI3 ;
  RECT 76.720 5.940 76.920 6.140 ;
  LAYER VI3 ;
  RECT 76.320 6.340 76.520 6.540 ;
  LAYER VI3 ;
  RECT 76.320 5.940 76.520 6.140 ;
  LAYER VI3 ;
  RECT 75.920 6.340 76.120 6.540 ;
  LAYER VI3 ;
  RECT 75.920 5.940 76.120 6.140 ;
  LAYER VI3 ;
  RECT 75.520 6.340 75.720 6.540 ;
  LAYER VI3 ;
  RECT 75.520 5.940 75.720 6.140 ;
  LAYER VI3 ;
  RECT 75.120 6.340 75.320 6.540 ;
  LAYER VI3 ;
  RECT 75.120 5.940 75.320 6.140 ;
  LAYER VI3 ;
  RECT 74.720 6.340 74.920 6.540 ;
  LAYER VI3 ;
  RECT 74.720 5.940 74.920 6.140 ;
  LAYER VI3 ;
  RECT 74.320 6.340 74.520 6.540 ;
  LAYER VI3 ;
  RECT 74.320 5.940 74.520 6.140 ;
  LAYER VI3 ;
  RECT 73.920 6.340 74.120 6.540 ;
  LAYER VI3 ;
  RECT 73.920 5.940 74.120 6.140 ;
  LAYER VI3 ;
  RECT 73.520 6.340 73.720 6.540 ;
  LAYER VI3 ;
  RECT 73.520 5.940 73.720 6.140 ;
  LAYER VI3 ;
  RECT 73.120 6.340 73.320 6.540 ;
  LAYER VI3 ;
  RECT 73.120 5.940 73.320 6.140 ;
  LAYER VI3 ;
  RECT 72.720 6.340 72.920 6.540 ;
  LAYER VI3 ;
  RECT 72.720 5.940 72.920 6.140 ;
  LAYER VI3 ;
  RECT 72.320 6.340 72.520 6.540 ;
  LAYER VI3 ;
  RECT 72.320 5.940 72.520 6.140 ;
  LAYER VI3 ;
  RECT 71.920 6.340 72.120 6.540 ;
  LAYER VI3 ;
  RECT 71.920 5.940 72.120 6.140 ;
  LAYER VI3 ;
  RECT 71.520 6.340 71.720 6.540 ;
  LAYER VI3 ;
  RECT 71.520 5.940 71.720 6.140 ;
  LAYER VI3 ;
  RECT 71.120 6.340 71.320 6.540 ;
  LAYER VI3 ;
  RECT 71.120 5.940 71.320 6.140 ;
  LAYER VI3 ;
  RECT 70.720 6.340 70.920 6.540 ;
  LAYER VI3 ;
  RECT 70.720 5.940 70.920 6.140 ;
  LAYER VI3 ;
  RECT 70.320 6.340 70.520 6.540 ;
  LAYER VI3 ;
  RECT 70.320 5.940 70.520 6.140 ;
  LAYER VI3 ;
  RECT 69.920 6.340 70.120 6.540 ;
  LAYER VI3 ;
  RECT 69.920 5.940 70.120 6.140 ;
  LAYER VI3 ;
  RECT 69.520 6.340 69.720 6.540 ;
  LAYER VI3 ;
  RECT 69.520 5.940 69.720 6.140 ;
  LAYER VI3 ;
  RECT 69.120 6.340 69.320 6.540 ;
  LAYER VI3 ;
  RECT 69.120 5.940 69.320 6.140 ;
  LAYER VI3 ;
  RECT 90.200 5.880 98.200 6.740 ;
  LAYER VI3 ;
  RECT 97.800 6.340 98.000 6.540 ;
  LAYER VI3 ;
  RECT 97.800 5.940 98.000 6.140 ;
  LAYER VI3 ;
  RECT 97.400 6.340 97.600 6.540 ;
  LAYER VI3 ;
  RECT 97.400 5.940 97.600 6.140 ;
  LAYER VI3 ;
  RECT 97.000 6.340 97.200 6.540 ;
  LAYER VI3 ;
  RECT 97.000 5.940 97.200 6.140 ;
  LAYER VI3 ;
  RECT 96.600 6.340 96.800 6.540 ;
  LAYER VI3 ;
  RECT 96.600 5.940 96.800 6.140 ;
  LAYER VI3 ;
  RECT 96.200 6.340 96.400 6.540 ;
  LAYER VI3 ;
  RECT 96.200 5.940 96.400 6.140 ;
  LAYER VI3 ;
  RECT 95.800 6.340 96.000 6.540 ;
  LAYER VI3 ;
  RECT 95.800 5.940 96.000 6.140 ;
  LAYER VI3 ;
  RECT 95.400 6.340 95.600 6.540 ;
  LAYER VI3 ;
  RECT 95.400 5.940 95.600 6.140 ;
  LAYER VI3 ;
  RECT 95.000 6.340 95.200 6.540 ;
  LAYER VI3 ;
  RECT 95.000 5.940 95.200 6.140 ;
  LAYER VI3 ;
  RECT 94.600 6.340 94.800 6.540 ;
  LAYER VI3 ;
  RECT 94.600 5.940 94.800 6.140 ;
  LAYER VI3 ;
  RECT 94.200 6.340 94.400 6.540 ;
  LAYER VI3 ;
  RECT 94.200 5.940 94.400 6.140 ;
  LAYER VI3 ;
  RECT 93.800 6.340 94.000 6.540 ;
  LAYER VI3 ;
  RECT 93.800 5.940 94.000 6.140 ;
  LAYER VI3 ;
  RECT 93.400 6.340 93.600 6.540 ;
  LAYER VI3 ;
  RECT 93.400 5.940 93.600 6.140 ;
  LAYER VI3 ;
  RECT 93.000 6.340 93.200 6.540 ;
  LAYER VI3 ;
  RECT 93.000 5.940 93.200 6.140 ;
  LAYER VI3 ;
  RECT 92.600 6.340 92.800 6.540 ;
  LAYER VI3 ;
  RECT 92.600 5.940 92.800 6.140 ;
  LAYER VI3 ;
  RECT 92.200 6.340 92.400 6.540 ;
  LAYER VI3 ;
  RECT 92.200 5.940 92.400 6.140 ;
  LAYER VI3 ;
  RECT 91.800 6.340 92.000 6.540 ;
  LAYER VI3 ;
  RECT 91.800 5.940 92.000 6.140 ;
  LAYER VI3 ;
  RECT 91.400 6.340 91.600 6.540 ;
  LAYER VI3 ;
  RECT 91.400 5.940 91.600 6.140 ;
  LAYER VI3 ;
  RECT 91.000 6.340 91.200 6.540 ;
  LAYER VI3 ;
  RECT 91.000 5.940 91.200 6.140 ;
  LAYER VI3 ;
  RECT 90.600 6.340 90.800 6.540 ;
  LAYER VI3 ;
  RECT 90.600 5.940 90.800 6.140 ;
  LAYER VI3 ;
  RECT 90.200 6.340 90.400 6.540 ;
  LAYER VI3 ;
  RECT 90.200 5.940 90.400 6.140 ;
  LAYER VI3 ;
  RECT 110.040 5.880 118.040 6.740 ;
  LAYER VI3 ;
  RECT 117.640 6.340 117.840 6.540 ;
  LAYER VI3 ;
  RECT 117.640 5.940 117.840 6.140 ;
  LAYER VI3 ;
  RECT 117.240 6.340 117.440 6.540 ;
  LAYER VI3 ;
  RECT 117.240 5.940 117.440 6.140 ;
  LAYER VI3 ;
  RECT 116.840 6.340 117.040 6.540 ;
  LAYER VI3 ;
  RECT 116.840 5.940 117.040 6.140 ;
  LAYER VI3 ;
  RECT 116.440 6.340 116.640 6.540 ;
  LAYER VI3 ;
  RECT 116.440 5.940 116.640 6.140 ;
  LAYER VI3 ;
  RECT 116.040 6.340 116.240 6.540 ;
  LAYER VI3 ;
  RECT 116.040 5.940 116.240 6.140 ;
  LAYER VI3 ;
  RECT 115.640 6.340 115.840 6.540 ;
  LAYER VI3 ;
  RECT 115.640 5.940 115.840 6.140 ;
  LAYER VI3 ;
  RECT 115.240 6.340 115.440 6.540 ;
  LAYER VI3 ;
  RECT 115.240 5.940 115.440 6.140 ;
  LAYER VI3 ;
  RECT 114.840 6.340 115.040 6.540 ;
  LAYER VI3 ;
  RECT 114.840 5.940 115.040 6.140 ;
  LAYER VI3 ;
  RECT 114.440 6.340 114.640 6.540 ;
  LAYER VI3 ;
  RECT 114.440 5.940 114.640 6.140 ;
  LAYER VI3 ;
  RECT 114.040 6.340 114.240 6.540 ;
  LAYER VI3 ;
  RECT 114.040 5.940 114.240 6.140 ;
  LAYER VI3 ;
  RECT 113.640 6.340 113.840 6.540 ;
  LAYER VI3 ;
  RECT 113.640 5.940 113.840 6.140 ;
  LAYER VI3 ;
  RECT 113.240 6.340 113.440 6.540 ;
  LAYER VI3 ;
  RECT 113.240 5.940 113.440 6.140 ;
  LAYER VI3 ;
  RECT 112.840 6.340 113.040 6.540 ;
  LAYER VI3 ;
  RECT 112.840 5.940 113.040 6.140 ;
  LAYER VI3 ;
  RECT 112.440 6.340 112.640 6.540 ;
  LAYER VI3 ;
  RECT 112.440 5.940 112.640 6.140 ;
  LAYER VI3 ;
  RECT 112.040 6.340 112.240 6.540 ;
  LAYER VI3 ;
  RECT 112.040 5.940 112.240 6.140 ;
  LAYER VI3 ;
  RECT 111.640 6.340 111.840 6.540 ;
  LAYER VI3 ;
  RECT 111.640 5.940 111.840 6.140 ;
  LAYER VI3 ;
  RECT 111.240 6.340 111.440 6.540 ;
  LAYER VI3 ;
  RECT 111.240 5.940 111.440 6.140 ;
  LAYER VI3 ;
  RECT 110.840 6.340 111.040 6.540 ;
  LAYER VI3 ;
  RECT 110.840 5.940 111.040 6.140 ;
  LAYER VI3 ;
  RECT 110.440 6.340 110.640 6.540 ;
  LAYER VI3 ;
  RECT 110.440 5.940 110.640 6.140 ;
  LAYER VI3 ;
  RECT 110.040 6.340 110.240 6.540 ;
  LAYER VI3 ;
  RECT 110.040 5.940 110.240 6.140 ;
  LAYER VI3 ;
  RECT 131.120 5.880 139.120 6.740 ;
  LAYER VI3 ;
  RECT 138.720 6.340 138.920 6.540 ;
  LAYER VI3 ;
  RECT 138.720 5.940 138.920 6.140 ;
  LAYER VI3 ;
  RECT 138.320 6.340 138.520 6.540 ;
  LAYER VI3 ;
  RECT 138.320 5.940 138.520 6.140 ;
  LAYER VI3 ;
  RECT 137.920 6.340 138.120 6.540 ;
  LAYER VI3 ;
  RECT 137.920 5.940 138.120 6.140 ;
  LAYER VI3 ;
  RECT 137.520 6.340 137.720 6.540 ;
  LAYER VI3 ;
  RECT 137.520 5.940 137.720 6.140 ;
  LAYER VI3 ;
  RECT 137.120 6.340 137.320 6.540 ;
  LAYER VI3 ;
  RECT 137.120 5.940 137.320 6.140 ;
  LAYER VI3 ;
  RECT 136.720 6.340 136.920 6.540 ;
  LAYER VI3 ;
  RECT 136.720 5.940 136.920 6.140 ;
  LAYER VI3 ;
  RECT 136.320 6.340 136.520 6.540 ;
  LAYER VI3 ;
  RECT 136.320 5.940 136.520 6.140 ;
  LAYER VI3 ;
  RECT 135.920 6.340 136.120 6.540 ;
  LAYER VI3 ;
  RECT 135.920 5.940 136.120 6.140 ;
  LAYER VI3 ;
  RECT 135.520 6.340 135.720 6.540 ;
  LAYER VI3 ;
  RECT 135.520 5.940 135.720 6.140 ;
  LAYER VI3 ;
  RECT 135.120 6.340 135.320 6.540 ;
  LAYER VI3 ;
  RECT 135.120 5.940 135.320 6.140 ;
  LAYER VI3 ;
  RECT 134.720 6.340 134.920 6.540 ;
  LAYER VI3 ;
  RECT 134.720 5.940 134.920 6.140 ;
  LAYER VI3 ;
  RECT 134.320 6.340 134.520 6.540 ;
  LAYER VI3 ;
  RECT 134.320 5.940 134.520 6.140 ;
  LAYER VI3 ;
  RECT 133.920 6.340 134.120 6.540 ;
  LAYER VI3 ;
  RECT 133.920 5.940 134.120 6.140 ;
  LAYER VI3 ;
  RECT 133.520 6.340 133.720 6.540 ;
  LAYER VI3 ;
  RECT 133.520 5.940 133.720 6.140 ;
  LAYER VI3 ;
  RECT 133.120 6.340 133.320 6.540 ;
  LAYER VI3 ;
  RECT 133.120 5.940 133.320 6.140 ;
  LAYER VI3 ;
  RECT 132.720 6.340 132.920 6.540 ;
  LAYER VI3 ;
  RECT 132.720 5.940 132.920 6.140 ;
  LAYER VI3 ;
  RECT 132.320 6.340 132.520 6.540 ;
  LAYER VI3 ;
  RECT 132.320 5.940 132.520 6.140 ;
  LAYER VI3 ;
  RECT 131.920 6.340 132.120 6.540 ;
  LAYER VI3 ;
  RECT 131.920 5.940 132.120 6.140 ;
  LAYER VI3 ;
  RECT 131.520 6.340 131.720 6.540 ;
  LAYER VI3 ;
  RECT 131.520 5.940 131.720 6.140 ;
  LAYER VI3 ;
  RECT 131.120 6.340 131.320 6.540 ;
  LAYER VI3 ;
  RECT 131.120 5.940 131.320 6.140 ;
  LAYER VI3 ;
  RECT 150.960 5.880 158.960 6.740 ;
  LAYER VI3 ;
  RECT 158.560 6.340 158.760 6.540 ;
  LAYER VI3 ;
  RECT 158.560 5.940 158.760 6.140 ;
  LAYER VI3 ;
  RECT 158.160 6.340 158.360 6.540 ;
  LAYER VI3 ;
  RECT 158.160 5.940 158.360 6.140 ;
  LAYER VI3 ;
  RECT 157.760 6.340 157.960 6.540 ;
  LAYER VI3 ;
  RECT 157.760 5.940 157.960 6.140 ;
  LAYER VI3 ;
  RECT 157.360 6.340 157.560 6.540 ;
  LAYER VI3 ;
  RECT 157.360 5.940 157.560 6.140 ;
  LAYER VI3 ;
  RECT 156.960 6.340 157.160 6.540 ;
  LAYER VI3 ;
  RECT 156.960 5.940 157.160 6.140 ;
  LAYER VI3 ;
  RECT 156.560 6.340 156.760 6.540 ;
  LAYER VI3 ;
  RECT 156.560 5.940 156.760 6.140 ;
  LAYER VI3 ;
  RECT 156.160 6.340 156.360 6.540 ;
  LAYER VI3 ;
  RECT 156.160 5.940 156.360 6.140 ;
  LAYER VI3 ;
  RECT 155.760 6.340 155.960 6.540 ;
  LAYER VI3 ;
  RECT 155.760 5.940 155.960 6.140 ;
  LAYER VI3 ;
  RECT 155.360 6.340 155.560 6.540 ;
  LAYER VI3 ;
  RECT 155.360 5.940 155.560 6.140 ;
  LAYER VI3 ;
  RECT 154.960 6.340 155.160 6.540 ;
  LAYER VI3 ;
  RECT 154.960 5.940 155.160 6.140 ;
  LAYER VI3 ;
  RECT 154.560 6.340 154.760 6.540 ;
  LAYER VI3 ;
  RECT 154.560 5.940 154.760 6.140 ;
  LAYER VI3 ;
  RECT 154.160 6.340 154.360 6.540 ;
  LAYER VI3 ;
  RECT 154.160 5.940 154.360 6.140 ;
  LAYER VI3 ;
  RECT 153.760 6.340 153.960 6.540 ;
  LAYER VI3 ;
  RECT 153.760 5.940 153.960 6.140 ;
  LAYER VI3 ;
  RECT 153.360 6.340 153.560 6.540 ;
  LAYER VI3 ;
  RECT 153.360 5.940 153.560 6.140 ;
  LAYER VI3 ;
  RECT 152.960 6.340 153.160 6.540 ;
  LAYER VI3 ;
  RECT 152.960 5.940 153.160 6.140 ;
  LAYER VI3 ;
  RECT 152.560 6.340 152.760 6.540 ;
  LAYER VI3 ;
  RECT 152.560 5.940 152.760 6.140 ;
  LAYER VI3 ;
  RECT 152.160 6.340 152.360 6.540 ;
  LAYER VI3 ;
  RECT 152.160 5.940 152.360 6.140 ;
  LAYER VI3 ;
  RECT 151.760 6.340 151.960 6.540 ;
  LAYER VI3 ;
  RECT 151.760 5.940 151.960 6.140 ;
  LAYER VI3 ;
  RECT 151.360 6.340 151.560 6.540 ;
  LAYER VI3 ;
  RECT 151.360 5.940 151.560 6.140 ;
  LAYER VI3 ;
  RECT 150.960 6.340 151.160 6.540 ;
  LAYER VI3 ;
  RECT 150.960 5.940 151.160 6.140 ;
  LAYER VI3 ;
  RECT 172.040 5.880 180.040 6.740 ;
  LAYER VI3 ;
  RECT 179.640 6.340 179.840 6.540 ;
  LAYER VI3 ;
  RECT 179.640 5.940 179.840 6.140 ;
  LAYER VI3 ;
  RECT 179.240 6.340 179.440 6.540 ;
  LAYER VI3 ;
  RECT 179.240 5.940 179.440 6.140 ;
  LAYER VI3 ;
  RECT 178.840 6.340 179.040 6.540 ;
  LAYER VI3 ;
  RECT 178.840 5.940 179.040 6.140 ;
  LAYER VI3 ;
  RECT 178.440 6.340 178.640 6.540 ;
  LAYER VI3 ;
  RECT 178.440 5.940 178.640 6.140 ;
  LAYER VI3 ;
  RECT 178.040 6.340 178.240 6.540 ;
  LAYER VI3 ;
  RECT 178.040 5.940 178.240 6.140 ;
  LAYER VI3 ;
  RECT 177.640 6.340 177.840 6.540 ;
  LAYER VI3 ;
  RECT 177.640 5.940 177.840 6.140 ;
  LAYER VI3 ;
  RECT 177.240 6.340 177.440 6.540 ;
  LAYER VI3 ;
  RECT 177.240 5.940 177.440 6.140 ;
  LAYER VI3 ;
  RECT 176.840 6.340 177.040 6.540 ;
  LAYER VI3 ;
  RECT 176.840 5.940 177.040 6.140 ;
  LAYER VI3 ;
  RECT 176.440 6.340 176.640 6.540 ;
  LAYER VI3 ;
  RECT 176.440 5.940 176.640 6.140 ;
  LAYER VI3 ;
  RECT 176.040 6.340 176.240 6.540 ;
  LAYER VI3 ;
  RECT 176.040 5.940 176.240 6.140 ;
  LAYER VI3 ;
  RECT 175.640 6.340 175.840 6.540 ;
  LAYER VI3 ;
  RECT 175.640 5.940 175.840 6.140 ;
  LAYER VI3 ;
  RECT 175.240 6.340 175.440 6.540 ;
  LAYER VI3 ;
  RECT 175.240 5.940 175.440 6.140 ;
  LAYER VI3 ;
  RECT 174.840 6.340 175.040 6.540 ;
  LAYER VI3 ;
  RECT 174.840 5.940 175.040 6.140 ;
  LAYER VI3 ;
  RECT 174.440 6.340 174.640 6.540 ;
  LAYER VI3 ;
  RECT 174.440 5.940 174.640 6.140 ;
  LAYER VI3 ;
  RECT 174.040 6.340 174.240 6.540 ;
  LAYER VI3 ;
  RECT 174.040 5.940 174.240 6.140 ;
  LAYER VI3 ;
  RECT 173.640 6.340 173.840 6.540 ;
  LAYER VI3 ;
  RECT 173.640 5.940 173.840 6.140 ;
  LAYER VI3 ;
  RECT 173.240 6.340 173.440 6.540 ;
  LAYER VI3 ;
  RECT 173.240 5.940 173.440 6.140 ;
  LAYER VI3 ;
  RECT 172.840 6.340 173.040 6.540 ;
  LAYER VI3 ;
  RECT 172.840 5.940 173.040 6.140 ;
  LAYER VI3 ;
  RECT 172.440 6.340 172.640 6.540 ;
  LAYER VI3 ;
  RECT 172.440 5.940 172.640 6.140 ;
  LAYER VI3 ;
  RECT 172.040 6.340 172.240 6.540 ;
  LAYER VI3 ;
  RECT 172.040 5.940 172.240 6.140 ;
  LAYER VI3 ;
  RECT 191.880 5.880 199.880 6.740 ;
  LAYER VI3 ;
  RECT 199.480 6.340 199.680 6.540 ;
  LAYER VI3 ;
  RECT 199.480 5.940 199.680 6.140 ;
  LAYER VI3 ;
  RECT 199.080 6.340 199.280 6.540 ;
  LAYER VI3 ;
  RECT 199.080 5.940 199.280 6.140 ;
  LAYER VI3 ;
  RECT 198.680 6.340 198.880 6.540 ;
  LAYER VI3 ;
  RECT 198.680 5.940 198.880 6.140 ;
  LAYER VI3 ;
  RECT 198.280 6.340 198.480 6.540 ;
  LAYER VI3 ;
  RECT 198.280 5.940 198.480 6.140 ;
  LAYER VI3 ;
  RECT 197.880 6.340 198.080 6.540 ;
  LAYER VI3 ;
  RECT 197.880 5.940 198.080 6.140 ;
  LAYER VI3 ;
  RECT 197.480 6.340 197.680 6.540 ;
  LAYER VI3 ;
  RECT 197.480 5.940 197.680 6.140 ;
  LAYER VI3 ;
  RECT 197.080 6.340 197.280 6.540 ;
  LAYER VI3 ;
  RECT 197.080 5.940 197.280 6.140 ;
  LAYER VI3 ;
  RECT 196.680 6.340 196.880 6.540 ;
  LAYER VI3 ;
  RECT 196.680 5.940 196.880 6.140 ;
  LAYER VI3 ;
  RECT 196.280 6.340 196.480 6.540 ;
  LAYER VI3 ;
  RECT 196.280 5.940 196.480 6.140 ;
  LAYER VI3 ;
  RECT 195.880 6.340 196.080 6.540 ;
  LAYER VI3 ;
  RECT 195.880 5.940 196.080 6.140 ;
  LAYER VI3 ;
  RECT 195.480 6.340 195.680 6.540 ;
  LAYER VI3 ;
  RECT 195.480 5.940 195.680 6.140 ;
  LAYER VI3 ;
  RECT 195.080 6.340 195.280 6.540 ;
  LAYER VI3 ;
  RECT 195.080 5.940 195.280 6.140 ;
  LAYER VI3 ;
  RECT 194.680 6.340 194.880 6.540 ;
  LAYER VI3 ;
  RECT 194.680 5.940 194.880 6.140 ;
  LAYER VI3 ;
  RECT 194.280 6.340 194.480 6.540 ;
  LAYER VI3 ;
  RECT 194.280 5.940 194.480 6.140 ;
  LAYER VI3 ;
  RECT 193.880 6.340 194.080 6.540 ;
  LAYER VI3 ;
  RECT 193.880 5.940 194.080 6.140 ;
  LAYER VI3 ;
  RECT 193.480 6.340 193.680 6.540 ;
  LAYER VI3 ;
  RECT 193.480 5.940 193.680 6.140 ;
  LAYER VI3 ;
  RECT 193.080 6.340 193.280 6.540 ;
  LAYER VI3 ;
  RECT 193.080 5.940 193.280 6.140 ;
  LAYER VI3 ;
  RECT 192.680 6.340 192.880 6.540 ;
  LAYER VI3 ;
  RECT 192.680 5.940 192.880 6.140 ;
  LAYER VI3 ;
  RECT 192.280 6.340 192.480 6.540 ;
  LAYER VI3 ;
  RECT 192.280 5.940 192.480 6.140 ;
  LAYER VI3 ;
  RECT 191.880 6.340 192.080 6.540 ;
  LAYER VI3 ;
  RECT 191.880 5.940 192.080 6.140 ;
  LAYER VI3 ;
  RECT 212.960 5.880 220.960 6.740 ;
  LAYER VI3 ;
  RECT 220.560 6.340 220.760 6.540 ;
  LAYER VI3 ;
  RECT 220.560 5.940 220.760 6.140 ;
  LAYER VI3 ;
  RECT 220.160 6.340 220.360 6.540 ;
  LAYER VI3 ;
  RECT 220.160 5.940 220.360 6.140 ;
  LAYER VI3 ;
  RECT 219.760 6.340 219.960 6.540 ;
  LAYER VI3 ;
  RECT 219.760 5.940 219.960 6.140 ;
  LAYER VI3 ;
  RECT 219.360 6.340 219.560 6.540 ;
  LAYER VI3 ;
  RECT 219.360 5.940 219.560 6.140 ;
  LAYER VI3 ;
  RECT 218.960 6.340 219.160 6.540 ;
  LAYER VI3 ;
  RECT 218.960 5.940 219.160 6.140 ;
  LAYER VI3 ;
  RECT 218.560 6.340 218.760 6.540 ;
  LAYER VI3 ;
  RECT 218.560 5.940 218.760 6.140 ;
  LAYER VI3 ;
  RECT 218.160 6.340 218.360 6.540 ;
  LAYER VI3 ;
  RECT 218.160 5.940 218.360 6.140 ;
  LAYER VI3 ;
  RECT 217.760 6.340 217.960 6.540 ;
  LAYER VI3 ;
  RECT 217.760 5.940 217.960 6.140 ;
  LAYER VI3 ;
  RECT 217.360 6.340 217.560 6.540 ;
  LAYER VI3 ;
  RECT 217.360 5.940 217.560 6.140 ;
  LAYER VI3 ;
  RECT 216.960 6.340 217.160 6.540 ;
  LAYER VI3 ;
  RECT 216.960 5.940 217.160 6.140 ;
  LAYER VI3 ;
  RECT 216.560 6.340 216.760 6.540 ;
  LAYER VI3 ;
  RECT 216.560 5.940 216.760 6.140 ;
  LAYER VI3 ;
  RECT 216.160 6.340 216.360 6.540 ;
  LAYER VI3 ;
  RECT 216.160 5.940 216.360 6.140 ;
  LAYER VI3 ;
  RECT 215.760 6.340 215.960 6.540 ;
  LAYER VI3 ;
  RECT 215.760 5.940 215.960 6.140 ;
  LAYER VI3 ;
  RECT 215.360 6.340 215.560 6.540 ;
  LAYER VI3 ;
  RECT 215.360 5.940 215.560 6.140 ;
  LAYER VI3 ;
  RECT 214.960 6.340 215.160 6.540 ;
  LAYER VI3 ;
  RECT 214.960 5.940 215.160 6.140 ;
  LAYER VI3 ;
  RECT 214.560 6.340 214.760 6.540 ;
  LAYER VI3 ;
  RECT 214.560 5.940 214.760 6.140 ;
  LAYER VI3 ;
  RECT 214.160 6.340 214.360 6.540 ;
  LAYER VI3 ;
  RECT 214.160 5.940 214.360 6.140 ;
  LAYER VI3 ;
  RECT 213.760 6.340 213.960 6.540 ;
  LAYER VI3 ;
  RECT 213.760 5.940 213.960 6.140 ;
  LAYER VI3 ;
  RECT 213.360 6.340 213.560 6.540 ;
  LAYER VI3 ;
  RECT 213.360 5.940 213.560 6.140 ;
  LAYER VI3 ;
  RECT 212.960 6.340 213.160 6.540 ;
  LAYER VI3 ;
  RECT 212.960 5.940 213.160 6.140 ;
  LAYER VI3 ;
  RECT 232.800 5.880 240.800 6.740 ;
  LAYER VI3 ;
  RECT 240.400 6.340 240.600 6.540 ;
  LAYER VI3 ;
  RECT 240.400 5.940 240.600 6.140 ;
  LAYER VI3 ;
  RECT 240.000 6.340 240.200 6.540 ;
  LAYER VI3 ;
  RECT 240.000 5.940 240.200 6.140 ;
  LAYER VI3 ;
  RECT 239.600 6.340 239.800 6.540 ;
  LAYER VI3 ;
  RECT 239.600 5.940 239.800 6.140 ;
  LAYER VI3 ;
  RECT 239.200 6.340 239.400 6.540 ;
  LAYER VI3 ;
  RECT 239.200 5.940 239.400 6.140 ;
  LAYER VI3 ;
  RECT 238.800 6.340 239.000 6.540 ;
  LAYER VI3 ;
  RECT 238.800 5.940 239.000 6.140 ;
  LAYER VI3 ;
  RECT 238.400 6.340 238.600 6.540 ;
  LAYER VI3 ;
  RECT 238.400 5.940 238.600 6.140 ;
  LAYER VI3 ;
  RECT 238.000 6.340 238.200 6.540 ;
  LAYER VI3 ;
  RECT 238.000 5.940 238.200 6.140 ;
  LAYER VI3 ;
  RECT 237.600 6.340 237.800 6.540 ;
  LAYER VI3 ;
  RECT 237.600 5.940 237.800 6.140 ;
  LAYER VI3 ;
  RECT 237.200 6.340 237.400 6.540 ;
  LAYER VI3 ;
  RECT 237.200 5.940 237.400 6.140 ;
  LAYER VI3 ;
  RECT 236.800 6.340 237.000 6.540 ;
  LAYER VI3 ;
  RECT 236.800 5.940 237.000 6.140 ;
  LAYER VI3 ;
  RECT 236.400 6.340 236.600 6.540 ;
  LAYER VI3 ;
  RECT 236.400 5.940 236.600 6.140 ;
  LAYER VI3 ;
  RECT 236.000 6.340 236.200 6.540 ;
  LAYER VI3 ;
  RECT 236.000 5.940 236.200 6.140 ;
  LAYER VI3 ;
  RECT 235.600 6.340 235.800 6.540 ;
  LAYER VI3 ;
  RECT 235.600 5.940 235.800 6.140 ;
  LAYER VI3 ;
  RECT 235.200 6.340 235.400 6.540 ;
  LAYER VI3 ;
  RECT 235.200 5.940 235.400 6.140 ;
  LAYER VI3 ;
  RECT 234.800 6.340 235.000 6.540 ;
  LAYER VI3 ;
  RECT 234.800 5.940 235.000 6.140 ;
  LAYER VI3 ;
  RECT 234.400 6.340 234.600 6.540 ;
  LAYER VI3 ;
  RECT 234.400 5.940 234.600 6.140 ;
  LAYER VI3 ;
  RECT 234.000 6.340 234.200 6.540 ;
  LAYER VI3 ;
  RECT 234.000 5.940 234.200 6.140 ;
  LAYER VI3 ;
  RECT 233.600 6.340 233.800 6.540 ;
  LAYER VI3 ;
  RECT 233.600 5.940 233.800 6.140 ;
  LAYER VI3 ;
  RECT 233.200 6.340 233.400 6.540 ;
  LAYER VI3 ;
  RECT 233.200 5.940 233.400 6.140 ;
  LAYER VI3 ;
  RECT 232.800 6.340 233.000 6.540 ;
  LAYER VI3 ;
  RECT 232.800 5.940 233.000 6.140 ;
  LAYER VI3 ;
  RECT 253.880 5.880 261.880 6.740 ;
  LAYER VI3 ;
  RECT 261.480 6.340 261.680 6.540 ;
  LAYER VI3 ;
  RECT 261.480 5.940 261.680 6.140 ;
  LAYER VI3 ;
  RECT 261.080 6.340 261.280 6.540 ;
  LAYER VI3 ;
  RECT 261.080 5.940 261.280 6.140 ;
  LAYER VI3 ;
  RECT 260.680 6.340 260.880 6.540 ;
  LAYER VI3 ;
  RECT 260.680 5.940 260.880 6.140 ;
  LAYER VI3 ;
  RECT 260.280 6.340 260.480 6.540 ;
  LAYER VI3 ;
  RECT 260.280 5.940 260.480 6.140 ;
  LAYER VI3 ;
  RECT 259.880 6.340 260.080 6.540 ;
  LAYER VI3 ;
  RECT 259.880 5.940 260.080 6.140 ;
  LAYER VI3 ;
  RECT 259.480 6.340 259.680 6.540 ;
  LAYER VI3 ;
  RECT 259.480 5.940 259.680 6.140 ;
  LAYER VI3 ;
  RECT 259.080 6.340 259.280 6.540 ;
  LAYER VI3 ;
  RECT 259.080 5.940 259.280 6.140 ;
  LAYER VI3 ;
  RECT 258.680 6.340 258.880 6.540 ;
  LAYER VI3 ;
  RECT 258.680 5.940 258.880 6.140 ;
  LAYER VI3 ;
  RECT 258.280 6.340 258.480 6.540 ;
  LAYER VI3 ;
  RECT 258.280 5.940 258.480 6.140 ;
  LAYER VI3 ;
  RECT 257.880 6.340 258.080 6.540 ;
  LAYER VI3 ;
  RECT 257.880 5.940 258.080 6.140 ;
  LAYER VI3 ;
  RECT 257.480 6.340 257.680 6.540 ;
  LAYER VI3 ;
  RECT 257.480 5.940 257.680 6.140 ;
  LAYER VI3 ;
  RECT 257.080 6.340 257.280 6.540 ;
  LAYER VI3 ;
  RECT 257.080 5.940 257.280 6.140 ;
  LAYER VI3 ;
  RECT 256.680 6.340 256.880 6.540 ;
  LAYER VI3 ;
  RECT 256.680 5.940 256.880 6.140 ;
  LAYER VI3 ;
  RECT 256.280 6.340 256.480 6.540 ;
  LAYER VI3 ;
  RECT 256.280 5.940 256.480 6.140 ;
  LAYER VI3 ;
  RECT 255.880 6.340 256.080 6.540 ;
  LAYER VI3 ;
  RECT 255.880 5.940 256.080 6.140 ;
  LAYER VI3 ;
  RECT 255.480 6.340 255.680 6.540 ;
  LAYER VI3 ;
  RECT 255.480 5.940 255.680 6.140 ;
  LAYER VI3 ;
  RECT 255.080 6.340 255.280 6.540 ;
  LAYER VI3 ;
  RECT 255.080 5.940 255.280 6.140 ;
  LAYER VI3 ;
  RECT 254.680 6.340 254.880 6.540 ;
  LAYER VI3 ;
  RECT 254.680 5.940 254.880 6.140 ;
  LAYER VI3 ;
  RECT 254.280 6.340 254.480 6.540 ;
  LAYER VI3 ;
  RECT 254.280 5.940 254.480 6.140 ;
  LAYER VI3 ;
  RECT 253.880 6.340 254.080 6.540 ;
  LAYER VI3 ;
  RECT 253.880 5.940 254.080 6.140 ;
  LAYER VI3 ;
  RECT 273.720 5.880 281.720 6.740 ;
  LAYER VI3 ;
  RECT 281.320 6.340 281.520 6.540 ;
  LAYER VI3 ;
  RECT 281.320 5.940 281.520 6.140 ;
  LAYER VI3 ;
  RECT 280.920 6.340 281.120 6.540 ;
  LAYER VI3 ;
  RECT 280.920 5.940 281.120 6.140 ;
  LAYER VI3 ;
  RECT 280.520 6.340 280.720 6.540 ;
  LAYER VI3 ;
  RECT 280.520 5.940 280.720 6.140 ;
  LAYER VI3 ;
  RECT 280.120 6.340 280.320 6.540 ;
  LAYER VI3 ;
  RECT 280.120 5.940 280.320 6.140 ;
  LAYER VI3 ;
  RECT 279.720 6.340 279.920 6.540 ;
  LAYER VI3 ;
  RECT 279.720 5.940 279.920 6.140 ;
  LAYER VI3 ;
  RECT 279.320 6.340 279.520 6.540 ;
  LAYER VI3 ;
  RECT 279.320 5.940 279.520 6.140 ;
  LAYER VI3 ;
  RECT 278.920 6.340 279.120 6.540 ;
  LAYER VI3 ;
  RECT 278.920 5.940 279.120 6.140 ;
  LAYER VI3 ;
  RECT 278.520 6.340 278.720 6.540 ;
  LAYER VI3 ;
  RECT 278.520 5.940 278.720 6.140 ;
  LAYER VI3 ;
  RECT 278.120 6.340 278.320 6.540 ;
  LAYER VI3 ;
  RECT 278.120 5.940 278.320 6.140 ;
  LAYER VI3 ;
  RECT 277.720 6.340 277.920 6.540 ;
  LAYER VI3 ;
  RECT 277.720 5.940 277.920 6.140 ;
  LAYER VI3 ;
  RECT 277.320 6.340 277.520 6.540 ;
  LAYER VI3 ;
  RECT 277.320 5.940 277.520 6.140 ;
  LAYER VI3 ;
  RECT 276.920 6.340 277.120 6.540 ;
  LAYER VI3 ;
  RECT 276.920 5.940 277.120 6.140 ;
  LAYER VI3 ;
  RECT 276.520 6.340 276.720 6.540 ;
  LAYER VI3 ;
  RECT 276.520 5.940 276.720 6.140 ;
  LAYER VI3 ;
  RECT 276.120 6.340 276.320 6.540 ;
  LAYER VI3 ;
  RECT 276.120 5.940 276.320 6.140 ;
  LAYER VI3 ;
  RECT 275.720 6.340 275.920 6.540 ;
  LAYER VI3 ;
  RECT 275.720 5.940 275.920 6.140 ;
  LAYER VI3 ;
  RECT 275.320 6.340 275.520 6.540 ;
  LAYER VI3 ;
  RECT 275.320 5.940 275.520 6.140 ;
  LAYER VI3 ;
  RECT 274.920 6.340 275.120 6.540 ;
  LAYER VI3 ;
  RECT 274.920 5.940 275.120 6.140 ;
  LAYER VI3 ;
  RECT 274.520 6.340 274.720 6.540 ;
  LAYER VI3 ;
  RECT 274.520 5.940 274.720 6.140 ;
  LAYER VI3 ;
  RECT 274.120 6.340 274.320 6.540 ;
  LAYER VI3 ;
  RECT 274.120 5.940 274.320 6.140 ;
  LAYER VI3 ;
  RECT 273.720 6.340 273.920 6.540 ;
  LAYER VI3 ;
  RECT 273.720 5.940 273.920 6.140 ;
  LAYER VI3 ;
  RECT 294.800 5.880 302.800 6.740 ;
  LAYER VI3 ;
  RECT 302.400 6.340 302.600 6.540 ;
  LAYER VI3 ;
  RECT 302.400 5.940 302.600 6.140 ;
  LAYER VI3 ;
  RECT 302.000 6.340 302.200 6.540 ;
  LAYER VI3 ;
  RECT 302.000 5.940 302.200 6.140 ;
  LAYER VI3 ;
  RECT 301.600 6.340 301.800 6.540 ;
  LAYER VI3 ;
  RECT 301.600 5.940 301.800 6.140 ;
  LAYER VI3 ;
  RECT 301.200 6.340 301.400 6.540 ;
  LAYER VI3 ;
  RECT 301.200 5.940 301.400 6.140 ;
  LAYER VI3 ;
  RECT 300.800 6.340 301.000 6.540 ;
  LAYER VI3 ;
  RECT 300.800 5.940 301.000 6.140 ;
  LAYER VI3 ;
  RECT 300.400 6.340 300.600 6.540 ;
  LAYER VI3 ;
  RECT 300.400 5.940 300.600 6.140 ;
  LAYER VI3 ;
  RECT 300.000 6.340 300.200 6.540 ;
  LAYER VI3 ;
  RECT 300.000 5.940 300.200 6.140 ;
  LAYER VI3 ;
  RECT 299.600 6.340 299.800 6.540 ;
  LAYER VI3 ;
  RECT 299.600 5.940 299.800 6.140 ;
  LAYER VI3 ;
  RECT 299.200 6.340 299.400 6.540 ;
  LAYER VI3 ;
  RECT 299.200 5.940 299.400 6.140 ;
  LAYER VI3 ;
  RECT 298.800 6.340 299.000 6.540 ;
  LAYER VI3 ;
  RECT 298.800 5.940 299.000 6.140 ;
  LAYER VI3 ;
  RECT 298.400 6.340 298.600 6.540 ;
  LAYER VI3 ;
  RECT 298.400 5.940 298.600 6.140 ;
  LAYER VI3 ;
  RECT 298.000 6.340 298.200 6.540 ;
  LAYER VI3 ;
  RECT 298.000 5.940 298.200 6.140 ;
  LAYER VI3 ;
  RECT 297.600 6.340 297.800 6.540 ;
  LAYER VI3 ;
  RECT 297.600 5.940 297.800 6.140 ;
  LAYER VI3 ;
  RECT 297.200 6.340 297.400 6.540 ;
  LAYER VI3 ;
  RECT 297.200 5.940 297.400 6.140 ;
  LAYER VI3 ;
  RECT 296.800 6.340 297.000 6.540 ;
  LAYER VI3 ;
  RECT 296.800 5.940 297.000 6.140 ;
  LAYER VI3 ;
  RECT 296.400 6.340 296.600 6.540 ;
  LAYER VI3 ;
  RECT 296.400 5.940 296.600 6.140 ;
  LAYER VI3 ;
  RECT 296.000 6.340 296.200 6.540 ;
  LAYER VI3 ;
  RECT 296.000 5.940 296.200 6.140 ;
  LAYER VI3 ;
  RECT 295.600 6.340 295.800 6.540 ;
  LAYER VI3 ;
  RECT 295.600 5.940 295.800 6.140 ;
  LAYER VI3 ;
  RECT 295.200 6.340 295.400 6.540 ;
  LAYER VI3 ;
  RECT 295.200 5.940 295.400 6.140 ;
  LAYER VI3 ;
  RECT 294.800 6.340 295.000 6.540 ;
  LAYER VI3 ;
  RECT 294.800 5.940 295.000 6.140 ;
  LAYER VI3 ;
  RECT 314.640 5.880 322.640 6.740 ;
  LAYER VI3 ;
  RECT 322.240 6.340 322.440 6.540 ;
  LAYER VI3 ;
  RECT 322.240 5.940 322.440 6.140 ;
  LAYER VI3 ;
  RECT 321.840 6.340 322.040 6.540 ;
  LAYER VI3 ;
  RECT 321.840 5.940 322.040 6.140 ;
  LAYER VI3 ;
  RECT 321.440 6.340 321.640 6.540 ;
  LAYER VI3 ;
  RECT 321.440 5.940 321.640 6.140 ;
  LAYER VI3 ;
  RECT 321.040 6.340 321.240 6.540 ;
  LAYER VI3 ;
  RECT 321.040 5.940 321.240 6.140 ;
  LAYER VI3 ;
  RECT 320.640 6.340 320.840 6.540 ;
  LAYER VI3 ;
  RECT 320.640 5.940 320.840 6.140 ;
  LAYER VI3 ;
  RECT 320.240 6.340 320.440 6.540 ;
  LAYER VI3 ;
  RECT 320.240 5.940 320.440 6.140 ;
  LAYER VI3 ;
  RECT 319.840 6.340 320.040 6.540 ;
  LAYER VI3 ;
  RECT 319.840 5.940 320.040 6.140 ;
  LAYER VI3 ;
  RECT 319.440 6.340 319.640 6.540 ;
  LAYER VI3 ;
  RECT 319.440 5.940 319.640 6.140 ;
  LAYER VI3 ;
  RECT 319.040 6.340 319.240 6.540 ;
  LAYER VI3 ;
  RECT 319.040 5.940 319.240 6.140 ;
  LAYER VI3 ;
  RECT 318.640 6.340 318.840 6.540 ;
  LAYER VI3 ;
  RECT 318.640 5.940 318.840 6.140 ;
  LAYER VI3 ;
  RECT 318.240 6.340 318.440 6.540 ;
  LAYER VI3 ;
  RECT 318.240 5.940 318.440 6.140 ;
  LAYER VI3 ;
  RECT 317.840 6.340 318.040 6.540 ;
  LAYER VI3 ;
  RECT 317.840 5.940 318.040 6.140 ;
  LAYER VI3 ;
  RECT 317.440 6.340 317.640 6.540 ;
  LAYER VI3 ;
  RECT 317.440 5.940 317.640 6.140 ;
  LAYER VI3 ;
  RECT 317.040 6.340 317.240 6.540 ;
  LAYER VI3 ;
  RECT 317.040 5.940 317.240 6.140 ;
  LAYER VI3 ;
  RECT 316.640 6.340 316.840 6.540 ;
  LAYER VI3 ;
  RECT 316.640 5.940 316.840 6.140 ;
  LAYER VI3 ;
  RECT 316.240 6.340 316.440 6.540 ;
  LAYER VI3 ;
  RECT 316.240 5.940 316.440 6.140 ;
  LAYER VI3 ;
  RECT 315.840 6.340 316.040 6.540 ;
  LAYER VI3 ;
  RECT 315.840 5.940 316.040 6.140 ;
  LAYER VI3 ;
  RECT 315.440 6.340 315.640 6.540 ;
  LAYER VI3 ;
  RECT 315.440 5.940 315.640 6.140 ;
  LAYER VI3 ;
  RECT 315.040 6.340 315.240 6.540 ;
  LAYER VI3 ;
  RECT 315.040 5.940 315.240 6.140 ;
  LAYER VI3 ;
  RECT 314.640 6.340 314.840 6.540 ;
  LAYER VI3 ;
  RECT 314.640 5.940 314.840 6.140 ;
  LAYER VI3 ;
  RECT 335.720 5.880 343.720 6.740 ;
  LAYER VI3 ;
  RECT 343.320 6.340 343.520 6.540 ;
  LAYER VI3 ;
  RECT 343.320 5.940 343.520 6.140 ;
  LAYER VI3 ;
  RECT 342.920 6.340 343.120 6.540 ;
  LAYER VI3 ;
  RECT 342.920 5.940 343.120 6.140 ;
  LAYER VI3 ;
  RECT 342.520 6.340 342.720 6.540 ;
  LAYER VI3 ;
  RECT 342.520 5.940 342.720 6.140 ;
  LAYER VI3 ;
  RECT 342.120 6.340 342.320 6.540 ;
  LAYER VI3 ;
  RECT 342.120 5.940 342.320 6.140 ;
  LAYER VI3 ;
  RECT 341.720 6.340 341.920 6.540 ;
  LAYER VI3 ;
  RECT 341.720 5.940 341.920 6.140 ;
  LAYER VI3 ;
  RECT 341.320 6.340 341.520 6.540 ;
  LAYER VI3 ;
  RECT 341.320 5.940 341.520 6.140 ;
  LAYER VI3 ;
  RECT 340.920 6.340 341.120 6.540 ;
  LAYER VI3 ;
  RECT 340.920 5.940 341.120 6.140 ;
  LAYER VI3 ;
  RECT 340.520 6.340 340.720 6.540 ;
  LAYER VI3 ;
  RECT 340.520 5.940 340.720 6.140 ;
  LAYER VI3 ;
  RECT 340.120 6.340 340.320 6.540 ;
  LAYER VI3 ;
  RECT 340.120 5.940 340.320 6.140 ;
  LAYER VI3 ;
  RECT 339.720 6.340 339.920 6.540 ;
  LAYER VI3 ;
  RECT 339.720 5.940 339.920 6.140 ;
  LAYER VI3 ;
  RECT 339.320 6.340 339.520 6.540 ;
  LAYER VI3 ;
  RECT 339.320 5.940 339.520 6.140 ;
  LAYER VI3 ;
  RECT 338.920 6.340 339.120 6.540 ;
  LAYER VI3 ;
  RECT 338.920 5.940 339.120 6.140 ;
  LAYER VI3 ;
  RECT 338.520 6.340 338.720 6.540 ;
  LAYER VI3 ;
  RECT 338.520 5.940 338.720 6.140 ;
  LAYER VI3 ;
  RECT 338.120 6.340 338.320 6.540 ;
  LAYER VI3 ;
  RECT 338.120 5.940 338.320 6.140 ;
  LAYER VI3 ;
  RECT 337.720 6.340 337.920 6.540 ;
  LAYER VI3 ;
  RECT 337.720 5.940 337.920 6.140 ;
  LAYER VI3 ;
  RECT 337.320 6.340 337.520 6.540 ;
  LAYER VI3 ;
  RECT 337.320 5.940 337.520 6.140 ;
  LAYER VI3 ;
  RECT 336.920 6.340 337.120 6.540 ;
  LAYER VI3 ;
  RECT 336.920 5.940 337.120 6.140 ;
  LAYER VI3 ;
  RECT 336.520 6.340 336.720 6.540 ;
  LAYER VI3 ;
  RECT 336.520 5.940 336.720 6.140 ;
  LAYER VI3 ;
  RECT 336.120 6.340 336.320 6.540 ;
  LAYER VI3 ;
  RECT 336.120 5.940 336.320 6.140 ;
  LAYER VI3 ;
  RECT 335.720 6.340 335.920 6.540 ;
  LAYER VI3 ;
  RECT 335.720 5.940 335.920 6.140 ;
  LAYER VI3 ;
  RECT 355.560 5.880 363.560 6.740 ;
  LAYER VI3 ;
  RECT 363.160 6.340 363.360 6.540 ;
  LAYER VI3 ;
  RECT 363.160 5.940 363.360 6.140 ;
  LAYER VI3 ;
  RECT 362.760 6.340 362.960 6.540 ;
  LAYER VI3 ;
  RECT 362.760 5.940 362.960 6.140 ;
  LAYER VI3 ;
  RECT 362.360 6.340 362.560 6.540 ;
  LAYER VI3 ;
  RECT 362.360 5.940 362.560 6.140 ;
  LAYER VI3 ;
  RECT 361.960 6.340 362.160 6.540 ;
  LAYER VI3 ;
  RECT 361.960 5.940 362.160 6.140 ;
  LAYER VI3 ;
  RECT 361.560 6.340 361.760 6.540 ;
  LAYER VI3 ;
  RECT 361.560 5.940 361.760 6.140 ;
  LAYER VI3 ;
  RECT 361.160 6.340 361.360 6.540 ;
  LAYER VI3 ;
  RECT 361.160 5.940 361.360 6.140 ;
  LAYER VI3 ;
  RECT 360.760 6.340 360.960 6.540 ;
  LAYER VI3 ;
  RECT 360.760 5.940 360.960 6.140 ;
  LAYER VI3 ;
  RECT 360.360 6.340 360.560 6.540 ;
  LAYER VI3 ;
  RECT 360.360 5.940 360.560 6.140 ;
  LAYER VI3 ;
  RECT 359.960 6.340 360.160 6.540 ;
  LAYER VI3 ;
  RECT 359.960 5.940 360.160 6.140 ;
  LAYER VI3 ;
  RECT 359.560 6.340 359.760 6.540 ;
  LAYER VI3 ;
  RECT 359.560 5.940 359.760 6.140 ;
  LAYER VI3 ;
  RECT 359.160 6.340 359.360 6.540 ;
  LAYER VI3 ;
  RECT 359.160 5.940 359.360 6.140 ;
  LAYER VI3 ;
  RECT 358.760 6.340 358.960 6.540 ;
  LAYER VI3 ;
  RECT 358.760 5.940 358.960 6.140 ;
  LAYER VI3 ;
  RECT 358.360 6.340 358.560 6.540 ;
  LAYER VI3 ;
  RECT 358.360 5.940 358.560 6.140 ;
  LAYER VI3 ;
  RECT 357.960 6.340 358.160 6.540 ;
  LAYER VI3 ;
  RECT 357.960 5.940 358.160 6.140 ;
  LAYER VI3 ;
  RECT 357.560 6.340 357.760 6.540 ;
  LAYER VI3 ;
  RECT 357.560 5.940 357.760 6.140 ;
  LAYER VI3 ;
  RECT 357.160 6.340 357.360 6.540 ;
  LAYER VI3 ;
  RECT 357.160 5.940 357.360 6.140 ;
  LAYER VI3 ;
  RECT 356.760 6.340 356.960 6.540 ;
  LAYER VI3 ;
  RECT 356.760 5.940 356.960 6.140 ;
  LAYER VI3 ;
  RECT 356.360 6.340 356.560 6.540 ;
  LAYER VI3 ;
  RECT 356.360 5.940 356.560 6.140 ;
  LAYER VI3 ;
  RECT 355.960 6.340 356.160 6.540 ;
  LAYER VI3 ;
  RECT 355.960 5.940 356.160 6.140 ;
  LAYER VI3 ;
  RECT 355.560 6.340 355.760 6.540 ;
  LAYER VI3 ;
  RECT 355.560 5.940 355.760 6.140 ;
  LAYER VI3 ;
  RECT 376.640 5.880 384.640 6.740 ;
  LAYER VI3 ;
  RECT 384.240 6.340 384.440 6.540 ;
  LAYER VI3 ;
  RECT 384.240 5.940 384.440 6.140 ;
  LAYER VI3 ;
  RECT 383.840 6.340 384.040 6.540 ;
  LAYER VI3 ;
  RECT 383.840 5.940 384.040 6.140 ;
  LAYER VI3 ;
  RECT 383.440 6.340 383.640 6.540 ;
  LAYER VI3 ;
  RECT 383.440 5.940 383.640 6.140 ;
  LAYER VI3 ;
  RECT 383.040 6.340 383.240 6.540 ;
  LAYER VI3 ;
  RECT 383.040 5.940 383.240 6.140 ;
  LAYER VI3 ;
  RECT 382.640 6.340 382.840 6.540 ;
  LAYER VI3 ;
  RECT 382.640 5.940 382.840 6.140 ;
  LAYER VI3 ;
  RECT 382.240 6.340 382.440 6.540 ;
  LAYER VI3 ;
  RECT 382.240 5.940 382.440 6.140 ;
  LAYER VI3 ;
  RECT 381.840 6.340 382.040 6.540 ;
  LAYER VI3 ;
  RECT 381.840 5.940 382.040 6.140 ;
  LAYER VI3 ;
  RECT 381.440 6.340 381.640 6.540 ;
  LAYER VI3 ;
  RECT 381.440 5.940 381.640 6.140 ;
  LAYER VI3 ;
  RECT 381.040 6.340 381.240 6.540 ;
  LAYER VI3 ;
  RECT 381.040 5.940 381.240 6.140 ;
  LAYER VI3 ;
  RECT 380.640 6.340 380.840 6.540 ;
  LAYER VI3 ;
  RECT 380.640 5.940 380.840 6.140 ;
  LAYER VI3 ;
  RECT 380.240 6.340 380.440 6.540 ;
  LAYER VI3 ;
  RECT 380.240 5.940 380.440 6.140 ;
  LAYER VI3 ;
  RECT 379.840 6.340 380.040 6.540 ;
  LAYER VI3 ;
  RECT 379.840 5.940 380.040 6.140 ;
  LAYER VI3 ;
  RECT 379.440 6.340 379.640 6.540 ;
  LAYER VI3 ;
  RECT 379.440 5.940 379.640 6.140 ;
  LAYER VI3 ;
  RECT 379.040 6.340 379.240 6.540 ;
  LAYER VI3 ;
  RECT 379.040 5.940 379.240 6.140 ;
  LAYER VI3 ;
  RECT 378.640 6.340 378.840 6.540 ;
  LAYER VI3 ;
  RECT 378.640 5.940 378.840 6.140 ;
  LAYER VI3 ;
  RECT 378.240 6.340 378.440 6.540 ;
  LAYER VI3 ;
  RECT 378.240 5.940 378.440 6.140 ;
  LAYER VI3 ;
  RECT 377.840 6.340 378.040 6.540 ;
  LAYER VI3 ;
  RECT 377.840 5.940 378.040 6.140 ;
  LAYER VI3 ;
  RECT 377.440 6.340 377.640 6.540 ;
  LAYER VI3 ;
  RECT 377.440 5.940 377.640 6.140 ;
  LAYER VI3 ;
  RECT 377.040 6.340 377.240 6.540 ;
  LAYER VI3 ;
  RECT 377.040 5.940 377.240 6.140 ;
  LAYER VI3 ;
  RECT 376.640 6.340 376.840 6.540 ;
  LAYER VI3 ;
  RECT 376.640 5.940 376.840 6.140 ;
  LAYER VI3 ;
  RECT 396.480 5.880 404.480 6.740 ;
  LAYER VI3 ;
  RECT 404.080 6.340 404.280 6.540 ;
  LAYER VI3 ;
  RECT 404.080 5.940 404.280 6.140 ;
  LAYER VI3 ;
  RECT 403.680 6.340 403.880 6.540 ;
  LAYER VI3 ;
  RECT 403.680 5.940 403.880 6.140 ;
  LAYER VI3 ;
  RECT 403.280 6.340 403.480 6.540 ;
  LAYER VI3 ;
  RECT 403.280 5.940 403.480 6.140 ;
  LAYER VI3 ;
  RECT 402.880 6.340 403.080 6.540 ;
  LAYER VI3 ;
  RECT 402.880 5.940 403.080 6.140 ;
  LAYER VI3 ;
  RECT 402.480 6.340 402.680 6.540 ;
  LAYER VI3 ;
  RECT 402.480 5.940 402.680 6.140 ;
  LAYER VI3 ;
  RECT 402.080 6.340 402.280 6.540 ;
  LAYER VI3 ;
  RECT 402.080 5.940 402.280 6.140 ;
  LAYER VI3 ;
  RECT 401.680 6.340 401.880 6.540 ;
  LAYER VI3 ;
  RECT 401.680 5.940 401.880 6.140 ;
  LAYER VI3 ;
  RECT 401.280 6.340 401.480 6.540 ;
  LAYER VI3 ;
  RECT 401.280 5.940 401.480 6.140 ;
  LAYER VI3 ;
  RECT 400.880 6.340 401.080 6.540 ;
  LAYER VI3 ;
  RECT 400.880 5.940 401.080 6.140 ;
  LAYER VI3 ;
  RECT 400.480 6.340 400.680 6.540 ;
  LAYER VI3 ;
  RECT 400.480 5.940 400.680 6.140 ;
  LAYER VI3 ;
  RECT 400.080 6.340 400.280 6.540 ;
  LAYER VI3 ;
  RECT 400.080 5.940 400.280 6.140 ;
  LAYER VI3 ;
  RECT 399.680 6.340 399.880 6.540 ;
  LAYER VI3 ;
  RECT 399.680 5.940 399.880 6.140 ;
  LAYER VI3 ;
  RECT 399.280 6.340 399.480 6.540 ;
  LAYER VI3 ;
  RECT 399.280 5.940 399.480 6.140 ;
  LAYER VI3 ;
  RECT 398.880 6.340 399.080 6.540 ;
  LAYER VI3 ;
  RECT 398.880 5.940 399.080 6.140 ;
  LAYER VI3 ;
  RECT 398.480 6.340 398.680 6.540 ;
  LAYER VI3 ;
  RECT 398.480 5.940 398.680 6.140 ;
  LAYER VI3 ;
  RECT 398.080 6.340 398.280 6.540 ;
  LAYER VI3 ;
  RECT 398.080 5.940 398.280 6.140 ;
  LAYER VI3 ;
  RECT 397.680 6.340 397.880 6.540 ;
  LAYER VI3 ;
  RECT 397.680 5.940 397.880 6.140 ;
  LAYER VI3 ;
  RECT 397.280 6.340 397.480 6.540 ;
  LAYER VI3 ;
  RECT 397.280 5.940 397.480 6.140 ;
  LAYER VI3 ;
  RECT 396.880 6.340 397.080 6.540 ;
  LAYER VI3 ;
  RECT 396.880 5.940 397.080 6.140 ;
  LAYER VI3 ;
  RECT 396.480 6.340 396.680 6.540 ;
  LAYER VI3 ;
  RECT 396.480 5.940 396.680 6.140 ;
  LAYER VI3 ;
  RECT 417.560 5.880 425.560 6.740 ;
  LAYER VI3 ;
  RECT 425.160 6.340 425.360 6.540 ;
  LAYER VI3 ;
  RECT 425.160 5.940 425.360 6.140 ;
  LAYER VI3 ;
  RECT 424.760 6.340 424.960 6.540 ;
  LAYER VI3 ;
  RECT 424.760 5.940 424.960 6.140 ;
  LAYER VI3 ;
  RECT 424.360 6.340 424.560 6.540 ;
  LAYER VI3 ;
  RECT 424.360 5.940 424.560 6.140 ;
  LAYER VI3 ;
  RECT 423.960 6.340 424.160 6.540 ;
  LAYER VI3 ;
  RECT 423.960 5.940 424.160 6.140 ;
  LAYER VI3 ;
  RECT 423.560 6.340 423.760 6.540 ;
  LAYER VI3 ;
  RECT 423.560 5.940 423.760 6.140 ;
  LAYER VI3 ;
  RECT 423.160 6.340 423.360 6.540 ;
  LAYER VI3 ;
  RECT 423.160 5.940 423.360 6.140 ;
  LAYER VI3 ;
  RECT 422.760 6.340 422.960 6.540 ;
  LAYER VI3 ;
  RECT 422.760 5.940 422.960 6.140 ;
  LAYER VI3 ;
  RECT 422.360 6.340 422.560 6.540 ;
  LAYER VI3 ;
  RECT 422.360 5.940 422.560 6.140 ;
  LAYER VI3 ;
  RECT 421.960 6.340 422.160 6.540 ;
  LAYER VI3 ;
  RECT 421.960 5.940 422.160 6.140 ;
  LAYER VI3 ;
  RECT 421.560 6.340 421.760 6.540 ;
  LAYER VI3 ;
  RECT 421.560 5.940 421.760 6.140 ;
  LAYER VI3 ;
  RECT 421.160 6.340 421.360 6.540 ;
  LAYER VI3 ;
  RECT 421.160 5.940 421.360 6.140 ;
  LAYER VI3 ;
  RECT 420.760 6.340 420.960 6.540 ;
  LAYER VI3 ;
  RECT 420.760 5.940 420.960 6.140 ;
  LAYER VI3 ;
  RECT 420.360 6.340 420.560 6.540 ;
  LAYER VI3 ;
  RECT 420.360 5.940 420.560 6.140 ;
  LAYER VI3 ;
  RECT 419.960 6.340 420.160 6.540 ;
  LAYER VI3 ;
  RECT 419.960 5.940 420.160 6.140 ;
  LAYER VI3 ;
  RECT 419.560 6.340 419.760 6.540 ;
  LAYER VI3 ;
  RECT 419.560 5.940 419.760 6.140 ;
  LAYER VI3 ;
  RECT 419.160 6.340 419.360 6.540 ;
  LAYER VI3 ;
  RECT 419.160 5.940 419.360 6.140 ;
  LAYER VI3 ;
  RECT 418.760 6.340 418.960 6.540 ;
  LAYER VI3 ;
  RECT 418.760 5.940 418.960 6.140 ;
  LAYER VI3 ;
  RECT 418.360 6.340 418.560 6.540 ;
  LAYER VI3 ;
  RECT 418.360 5.940 418.560 6.140 ;
  LAYER VI3 ;
  RECT 417.960 6.340 418.160 6.540 ;
  LAYER VI3 ;
  RECT 417.960 5.940 418.160 6.140 ;
  LAYER VI3 ;
  RECT 417.560 6.340 417.760 6.540 ;
  LAYER VI3 ;
  RECT 417.560 5.940 417.760 6.140 ;
  LAYER VI3 ;
  RECT 437.400 5.880 445.400 6.740 ;
  LAYER VI3 ;
  RECT 445.000 6.340 445.200 6.540 ;
  LAYER VI3 ;
  RECT 445.000 5.940 445.200 6.140 ;
  LAYER VI3 ;
  RECT 444.600 6.340 444.800 6.540 ;
  LAYER VI3 ;
  RECT 444.600 5.940 444.800 6.140 ;
  LAYER VI3 ;
  RECT 444.200 6.340 444.400 6.540 ;
  LAYER VI3 ;
  RECT 444.200 5.940 444.400 6.140 ;
  LAYER VI3 ;
  RECT 443.800 6.340 444.000 6.540 ;
  LAYER VI3 ;
  RECT 443.800 5.940 444.000 6.140 ;
  LAYER VI3 ;
  RECT 443.400 6.340 443.600 6.540 ;
  LAYER VI3 ;
  RECT 443.400 5.940 443.600 6.140 ;
  LAYER VI3 ;
  RECT 443.000 6.340 443.200 6.540 ;
  LAYER VI3 ;
  RECT 443.000 5.940 443.200 6.140 ;
  LAYER VI3 ;
  RECT 442.600 6.340 442.800 6.540 ;
  LAYER VI3 ;
  RECT 442.600 5.940 442.800 6.140 ;
  LAYER VI3 ;
  RECT 442.200 6.340 442.400 6.540 ;
  LAYER VI3 ;
  RECT 442.200 5.940 442.400 6.140 ;
  LAYER VI3 ;
  RECT 441.800 6.340 442.000 6.540 ;
  LAYER VI3 ;
  RECT 441.800 5.940 442.000 6.140 ;
  LAYER VI3 ;
  RECT 441.400 6.340 441.600 6.540 ;
  LAYER VI3 ;
  RECT 441.400 5.940 441.600 6.140 ;
  LAYER VI3 ;
  RECT 441.000 6.340 441.200 6.540 ;
  LAYER VI3 ;
  RECT 441.000 5.940 441.200 6.140 ;
  LAYER VI3 ;
  RECT 440.600 6.340 440.800 6.540 ;
  LAYER VI3 ;
  RECT 440.600 5.940 440.800 6.140 ;
  LAYER VI3 ;
  RECT 440.200 6.340 440.400 6.540 ;
  LAYER VI3 ;
  RECT 440.200 5.940 440.400 6.140 ;
  LAYER VI3 ;
  RECT 439.800 6.340 440.000 6.540 ;
  LAYER VI3 ;
  RECT 439.800 5.940 440.000 6.140 ;
  LAYER VI3 ;
  RECT 439.400 6.340 439.600 6.540 ;
  LAYER VI3 ;
  RECT 439.400 5.940 439.600 6.140 ;
  LAYER VI3 ;
  RECT 439.000 6.340 439.200 6.540 ;
  LAYER VI3 ;
  RECT 439.000 5.940 439.200 6.140 ;
  LAYER VI3 ;
  RECT 438.600 6.340 438.800 6.540 ;
  LAYER VI3 ;
  RECT 438.600 5.940 438.800 6.140 ;
  LAYER VI3 ;
  RECT 438.200 6.340 438.400 6.540 ;
  LAYER VI3 ;
  RECT 438.200 5.940 438.400 6.140 ;
  LAYER VI3 ;
  RECT 437.800 6.340 438.000 6.540 ;
  LAYER VI3 ;
  RECT 437.800 5.940 438.000 6.140 ;
  LAYER VI3 ;
  RECT 437.400 6.340 437.600 6.540 ;
  LAYER VI3 ;
  RECT 437.400 5.940 437.600 6.140 ;
  LAYER VI3 ;
  RECT 458.480 5.880 466.480 6.740 ;
  LAYER VI3 ;
  RECT 466.080 6.340 466.280 6.540 ;
  LAYER VI3 ;
  RECT 466.080 5.940 466.280 6.140 ;
  LAYER VI3 ;
  RECT 465.680 6.340 465.880 6.540 ;
  LAYER VI3 ;
  RECT 465.680 5.940 465.880 6.140 ;
  LAYER VI3 ;
  RECT 465.280 6.340 465.480 6.540 ;
  LAYER VI3 ;
  RECT 465.280 5.940 465.480 6.140 ;
  LAYER VI3 ;
  RECT 464.880 6.340 465.080 6.540 ;
  LAYER VI3 ;
  RECT 464.880 5.940 465.080 6.140 ;
  LAYER VI3 ;
  RECT 464.480 6.340 464.680 6.540 ;
  LAYER VI3 ;
  RECT 464.480 5.940 464.680 6.140 ;
  LAYER VI3 ;
  RECT 464.080 6.340 464.280 6.540 ;
  LAYER VI3 ;
  RECT 464.080 5.940 464.280 6.140 ;
  LAYER VI3 ;
  RECT 463.680 6.340 463.880 6.540 ;
  LAYER VI3 ;
  RECT 463.680 5.940 463.880 6.140 ;
  LAYER VI3 ;
  RECT 463.280 6.340 463.480 6.540 ;
  LAYER VI3 ;
  RECT 463.280 5.940 463.480 6.140 ;
  LAYER VI3 ;
  RECT 462.880 6.340 463.080 6.540 ;
  LAYER VI3 ;
  RECT 462.880 5.940 463.080 6.140 ;
  LAYER VI3 ;
  RECT 462.480 6.340 462.680 6.540 ;
  LAYER VI3 ;
  RECT 462.480 5.940 462.680 6.140 ;
  LAYER VI3 ;
  RECT 462.080 6.340 462.280 6.540 ;
  LAYER VI3 ;
  RECT 462.080 5.940 462.280 6.140 ;
  LAYER VI3 ;
  RECT 461.680 6.340 461.880 6.540 ;
  LAYER VI3 ;
  RECT 461.680 5.940 461.880 6.140 ;
  LAYER VI3 ;
  RECT 461.280 6.340 461.480 6.540 ;
  LAYER VI3 ;
  RECT 461.280 5.940 461.480 6.140 ;
  LAYER VI3 ;
  RECT 460.880 6.340 461.080 6.540 ;
  LAYER VI3 ;
  RECT 460.880 5.940 461.080 6.140 ;
  LAYER VI3 ;
  RECT 460.480 6.340 460.680 6.540 ;
  LAYER VI3 ;
  RECT 460.480 5.940 460.680 6.140 ;
  LAYER VI3 ;
  RECT 460.080 6.340 460.280 6.540 ;
  LAYER VI3 ;
  RECT 460.080 5.940 460.280 6.140 ;
  LAYER VI3 ;
  RECT 459.680 6.340 459.880 6.540 ;
  LAYER VI3 ;
  RECT 459.680 5.940 459.880 6.140 ;
  LAYER VI3 ;
  RECT 459.280 6.340 459.480 6.540 ;
  LAYER VI3 ;
  RECT 459.280 5.940 459.480 6.140 ;
  LAYER VI3 ;
  RECT 458.880 6.340 459.080 6.540 ;
  LAYER VI3 ;
  RECT 458.880 5.940 459.080 6.140 ;
  LAYER VI3 ;
  RECT 458.480 6.340 458.680 6.540 ;
  LAYER VI3 ;
  RECT 458.480 5.940 458.680 6.140 ;
  LAYER VI3 ;
  RECT 478.320 5.880 486.320 6.740 ;
  LAYER VI3 ;
  RECT 485.920 6.340 486.120 6.540 ;
  LAYER VI3 ;
  RECT 485.920 5.940 486.120 6.140 ;
  LAYER VI3 ;
  RECT 485.520 6.340 485.720 6.540 ;
  LAYER VI3 ;
  RECT 485.520 5.940 485.720 6.140 ;
  LAYER VI3 ;
  RECT 485.120 6.340 485.320 6.540 ;
  LAYER VI3 ;
  RECT 485.120 5.940 485.320 6.140 ;
  LAYER VI3 ;
  RECT 484.720 6.340 484.920 6.540 ;
  LAYER VI3 ;
  RECT 484.720 5.940 484.920 6.140 ;
  LAYER VI3 ;
  RECT 484.320 6.340 484.520 6.540 ;
  LAYER VI3 ;
  RECT 484.320 5.940 484.520 6.140 ;
  LAYER VI3 ;
  RECT 483.920 6.340 484.120 6.540 ;
  LAYER VI3 ;
  RECT 483.920 5.940 484.120 6.140 ;
  LAYER VI3 ;
  RECT 483.520 6.340 483.720 6.540 ;
  LAYER VI3 ;
  RECT 483.520 5.940 483.720 6.140 ;
  LAYER VI3 ;
  RECT 483.120 6.340 483.320 6.540 ;
  LAYER VI3 ;
  RECT 483.120 5.940 483.320 6.140 ;
  LAYER VI3 ;
  RECT 482.720 6.340 482.920 6.540 ;
  LAYER VI3 ;
  RECT 482.720 5.940 482.920 6.140 ;
  LAYER VI3 ;
  RECT 482.320 6.340 482.520 6.540 ;
  LAYER VI3 ;
  RECT 482.320 5.940 482.520 6.140 ;
  LAYER VI3 ;
  RECT 481.920 6.340 482.120 6.540 ;
  LAYER VI3 ;
  RECT 481.920 5.940 482.120 6.140 ;
  LAYER VI3 ;
  RECT 481.520 6.340 481.720 6.540 ;
  LAYER VI3 ;
  RECT 481.520 5.940 481.720 6.140 ;
  LAYER VI3 ;
  RECT 481.120 6.340 481.320 6.540 ;
  LAYER VI3 ;
  RECT 481.120 5.940 481.320 6.140 ;
  LAYER VI3 ;
  RECT 480.720 6.340 480.920 6.540 ;
  LAYER VI3 ;
  RECT 480.720 5.940 480.920 6.140 ;
  LAYER VI3 ;
  RECT 480.320 6.340 480.520 6.540 ;
  LAYER VI3 ;
  RECT 480.320 5.940 480.520 6.140 ;
  LAYER VI3 ;
  RECT 479.920 6.340 480.120 6.540 ;
  LAYER VI3 ;
  RECT 479.920 5.940 480.120 6.140 ;
  LAYER VI3 ;
  RECT 479.520 6.340 479.720 6.540 ;
  LAYER VI3 ;
  RECT 479.520 5.940 479.720 6.140 ;
  LAYER VI3 ;
  RECT 479.120 6.340 479.320 6.540 ;
  LAYER VI3 ;
  RECT 479.120 5.940 479.320 6.140 ;
  LAYER VI3 ;
  RECT 478.720 6.340 478.920 6.540 ;
  LAYER VI3 ;
  RECT 478.720 5.940 478.920 6.140 ;
  LAYER VI3 ;
  RECT 478.320 6.340 478.520 6.540 ;
  LAYER VI3 ;
  RECT 478.320 5.940 478.520 6.140 ;
  LAYER VI3 ;
  RECT 499.400 5.880 507.400 6.740 ;
  LAYER VI3 ;
  RECT 507.000 6.340 507.200 6.540 ;
  LAYER VI3 ;
  RECT 507.000 5.940 507.200 6.140 ;
  LAYER VI3 ;
  RECT 506.600 6.340 506.800 6.540 ;
  LAYER VI3 ;
  RECT 506.600 5.940 506.800 6.140 ;
  LAYER VI3 ;
  RECT 506.200 6.340 506.400 6.540 ;
  LAYER VI3 ;
  RECT 506.200 5.940 506.400 6.140 ;
  LAYER VI3 ;
  RECT 505.800 6.340 506.000 6.540 ;
  LAYER VI3 ;
  RECT 505.800 5.940 506.000 6.140 ;
  LAYER VI3 ;
  RECT 505.400 6.340 505.600 6.540 ;
  LAYER VI3 ;
  RECT 505.400 5.940 505.600 6.140 ;
  LAYER VI3 ;
  RECT 505.000 6.340 505.200 6.540 ;
  LAYER VI3 ;
  RECT 505.000 5.940 505.200 6.140 ;
  LAYER VI3 ;
  RECT 504.600 6.340 504.800 6.540 ;
  LAYER VI3 ;
  RECT 504.600 5.940 504.800 6.140 ;
  LAYER VI3 ;
  RECT 504.200 6.340 504.400 6.540 ;
  LAYER VI3 ;
  RECT 504.200 5.940 504.400 6.140 ;
  LAYER VI3 ;
  RECT 503.800 6.340 504.000 6.540 ;
  LAYER VI3 ;
  RECT 503.800 5.940 504.000 6.140 ;
  LAYER VI3 ;
  RECT 503.400 6.340 503.600 6.540 ;
  LAYER VI3 ;
  RECT 503.400 5.940 503.600 6.140 ;
  LAYER VI3 ;
  RECT 503.000 6.340 503.200 6.540 ;
  LAYER VI3 ;
  RECT 503.000 5.940 503.200 6.140 ;
  LAYER VI3 ;
  RECT 502.600 6.340 502.800 6.540 ;
  LAYER VI3 ;
  RECT 502.600 5.940 502.800 6.140 ;
  LAYER VI3 ;
  RECT 502.200 6.340 502.400 6.540 ;
  LAYER VI3 ;
  RECT 502.200 5.940 502.400 6.140 ;
  LAYER VI3 ;
  RECT 501.800 6.340 502.000 6.540 ;
  LAYER VI3 ;
  RECT 501.800 5.940 502.000 6.140 ;
  LAYER VI3 ;
  RECT 501.400 6.340 501.600 6.540 ;
  LAYER VI3 ;
  RECT 501.400 5.940 501.600 6.140 ;
  LAYER VI3 ;
  RECT 501.000 6.340 501.200 6.540 ;
  LAYER VI3 ;
  RECT 501.000 5.940 501.200 6.140 ;
  LAYER VI3 ;
  RECT 500.600 6.340 500.800 6.540 ;
  LAYER VI3 ;
  RECT 500.600 5.940 500.800 6.140 ;
  LAYER VI3 ;
  RECT 500.200 6.340 500.400 6.540 ;
  LAYER VI3 ;
  RECT 500.200 5.940 500.400 6.140 ;
  LAYER VI3 ;
  RECT 499.800 6.340 500.000 6.540 ;
  LAYER VI3 ;
  RECT 499.800 5.940 500.000 6.140 ;
  LAYER VI3 ;
  RECT 499.400 6.340 499.600 6.540 ;
  LAYER VI3 ;
  RECT 499.400 5.940 499.600 6.140 ;
  LAYER VI3 ;
  RECT 519.240 5.880 527.240 6.740 ;
  LAYER VI3 ;
  RECT 526.840 6.340 527.040 6.540 ;
  LAYER VI3 ;
  RECT 526.840 5.940 527.040 6.140 ;
  LAYER VI3 ;
  RECT 526.440 6.340 526.640 6.540 ;
  LAYER VI3 ;
  RECT 526.440 5.940 526.640 6.140 ;
  LAYER VI3 ;
  RECT 526.040 6.340 526.240 6.540 ;
  LAYER VI3 ;
  RECT 526.040 5.940 526.240 6.140 ;
  LAYER VI3 ;
  RECT 525.640 6.340 525.840 6.540 ;
  LAYER VI3 ;
  RECT 525.640 5.940 525.840 6.140 ;
  LAYER VI3 ;
  RECT 525.240 6.340 525.440 6.540 ;
  LAYER VI3 ;
  RECT 525.240 5.940 525.440 6.140 ;
  LAYER VI3 ;
  RECT 524.840 6.340 525.040 6.540 ;
  LAYER VI3 ;
  RECT 524.840 5.940 525.040 6.140 ;
  LAYER VI3 ;
  RECT 524.440 6.340 524.640 6.540 ;
  LAYER VI3 ;
  RECT 524.440 5.940 524.640 6.140 ;
  LAYER VI3 ;
  RECT 524.040 6.340 524.240 6.540 ;
  LAYER VI3 ;
  RECT 524.040 5.940 524.240 6.140 ;
  LAYER VI3 ;
  RECT 523.640 6.340 523.840 6.540 ;
  LAYER VI3 ;
  RECT 523.640 5.940 523.840 6.140 ;
  LAYER VI3 ;
  RECT 523.240 6.340 523.440 6.540 ;
  LAYER VI3 ;
  RECT 523.240 5.940 523.440 6.140 ;
  LAYER VI3 ;
  RECT 522.840 6.340 523.040 6.540 ;
  LAYER VI3 ;
  RECT 522.840 5.940 523.040 6.140 ;
  LAYER VI3 ;
  RECT 522.440 6.340 522.640 6.540 ;
  LAYER VI3 ;
  RECT 522.440 5.940 522.640 6.140 ;
  LAYER VI3 ;
  RECT 522.040 6.340 522.240 6.540 ;
  LAYER VI3 ;
  RECT 522.040 5.940 522.240 6.140 ;
  LAYER VI3 ;
  RECT 521.640 6.340 521.840 6.540 ;
  LAYER VI3 ;
  RECT 521.640 5.940 521.840 6.140 ;
  LAYER VI3 ;
  RECT 521.240 6.340 521.440 6.540 ;
  LAYER VI3 ;
  RECT 521.240 5.940 521.440 6.140 ;
  LAYER VI3 ;
  RECT 520.840 6.340 521.040 6.540 ;
  LAYER VI3 ;
  RECT 520.840 5.940 521.040 6.140 ;
  LAYER VI3 ;
  RECT 520.440 6.340 520.640 6.540 ;
  LAYER VI3 ;
  RECT 520.440 5.940 520.640 6.140 ;
  LAYER VI3 ;
  RECT 520.040 6.340 520.240 6.540 ;
  LAYER VI3 ;
  RECT 520.040 5.940 520.240 6.140 ;
  LAYER VI3 ;
  RECT 519.640 6.340 519.840 6.540 ;
  LAYER VI3 ;
  RECT 519.640 5.940 519.840 6.140 ;
  LAYER VI3 ;
  RECT 519.240 6.340 519.440 6.540 ;
  LAYER VI3 ;
  RECT 519.240 5.940 519.440 6.140 ;
  LAYER VI3 ;
  RECT 540.320 5.880 548.320 6.740 ;
  LAYER VI3 ;
  RECT 547.920 6.340 548.120 6.540 ;
  LAYER VI3 ;
  RECT 547.920 5.940 548.120 6.140 ;
  LAYER VI3 ;
  RECT 547.520 6.340 547.720 6.540 ;
  LAYER VI3 ;
  RECT 547.520 5.940 547.720 6.140 ;
  LAYER VI3 ;
  RECT 547.120 6.340 547.320 6.540 ;
  LAYER VI3 ;
  RECT 547.120 5.940 547.320 6.140 ;
  LAYER VI3 ;
  RECT 546.720 6.340 546.920 6.540 ;
  LAYER VI3 ;
  RECT 546.720 5.940 546.920 6.140 ;
  LAYER VI3 ;
  RECT 546.320 6.340 546.520 6.540 ;
  LAYER VI3 ;
  RECT 546.320 5.940 546.520 6.140 ;
  LAYER VI3 ;
  RECT 545.920 6.340 546.120 6.540 ;
  LAYER VI3 ;
  RECT 545.920 5.940 546.120 6.140 ;
  LAYER VI3 ;
  RECT 545.520 6.340 545.720 6.540 ;
  LAYER VI3 ;
  RECT 545.520 5.940 545.720 6.140 ;
  LAYER VI3 ;
  RECT 545.120 6.340 545.320 6.540 ;
  LAYER VI3 ;
  RECT 545.120 5.940 545.320 6.140 ;
  LAYER VI3 ;
  RECT 544.720 6.340 544.920 6.540 ;
  LAYER VI3 ;
  RECT 544.720 5.940 544.920 6.140 ;
  LAYER VI3 ;
  RECT 544.320 6.340 544.520 6.540 ;
  LAYER VI3 ;
  RECT 544.320 5.940 544.520 6.140 ;
  LAYER VI3 ;
  RECT 543.920 6.340 544.120 6.540 ;
  LAYER VI3 ;
  RECT 543.920 5.940 544.120 6.140 ;
  LAYER VI3 ;
  RECT 543.520 6.340 543.720 6.540 ;
  LAYER VI3 ;
  RECT 543.520 5.940 543.720 6.140 ;
  LAYER VI3 ;
  RECT 543.120 6.340 543.320 6.540 ;
  LAYER VI3 ;
  RECT 543.120 5.940 543.320 6.140 ;
  LAYER VI3 ;
  RECT 542.720 6.340 542.920 6.540 ;
  LAYER VI3 ;
  RECT 542.720 5.940 542.920 6.140 ;
  LAYER VI3 ;
  RECT 542.320 6.340 542.520 6.540 ;
  LAYER VI3 ;
  RECT 542.320 5.940 542.520 6.140 ;
  LAYER VI3 ;
  RECT 541.920 6.340 542.120 6.540 ;
  LAYER VI3 ;
  RECT 541.920 5.940 542.120 6.140 ;
  LAYER VI3 ;
  RECT 541.520 6.340 541.720 6.540 ;
  LAYER VI3 ;
  RECT 541.520 5.940 541.720 6.140 ;
  LAYER VI3 ;
  RECT 541.120 6.340 541.320 6.540 ;
  LAYER VI3 ;
  RECT 541.120 5.940 541.320 6.140 ;
  LAYER VI3 ;
  RECT 540.720 6.340 540.920 6.540 ;
  LAYER VI3 ;
  RECT 540.720 5.940 540.920 6.140 ;
  LAYER VI3 ;
  RECT 540.320 6.340 540.520 6.540 ;
  LAYER VI3 ;
  RECT 540.320 5.940 540.520 6.140 ;
  LAYER VI3 ;
  RECT 560.160 5.880 568.160 6.740 ;
  LAYER VI3 ;
  RECT 567.760 6.340 567.960 6.540 ;
  LAYER VI3 ;
  RECT 567.760 5.940 567.960 6.140 ;
  LAYER VI3 ;
  RECT 567.360 6.340 567.560 6.540 ;
  LAYER VI3 ;
  RECT 567.360 5.940 567.560 6.140 ;
  LAYER VI3 ;
  RECT 566.960 6.340 567.160 6.540 ;
  LAYER VI3 ;
  RECT 566.960 5.940 567.160 6.140 ;
  LAYER VI3 ;
  RECT 566.560 6.340 566.760 6.540 ;
  LAYER VI3 ;
  RECT 566.560 5.940 566.760 6.140 ;
  LAYER VI3 ;
  RECT 566.160 6.340 566.360 6.540 ;
  LAYER VI3 ;
  RECT 566.160 5.940 566.360 6.140 ;
  LAYER VI3 ;
  RECT 565.760 6.340 565.960 6.540 ;
  LAYER VI3 ;
  RECT 565.760 5.940 565.960 6.140 ;
  LAYER VI3 ;
  RECT 565.360 6.340 565.560 6.540 ;
  LAYER VI3 ;
  RECT 565.360 5.940 565.560 6.140 ;
  LAYER VI3 ;
  RECT 564.960 6.340 565.160 6.540 ;
  LAYER VI3 ;
  RECT 564.960 5.940 565.160 6.140 ;
  LAYER VI3 ;
  RECT 564.560 6.340 564.760 6.540 ;
  LAYER VI3 ;
  RECT 564.560 5.940 564.760 6.140 ;
  LAYER VI3 ;
  RECT 564.160 6.340 564.360 6.540 ;
  LAYER VI3 ;
  RECT 564.160 5.940 564.360 6.140 ;
  LAYER VI3 ;
  RECT 563.760 6.340 563.960 6.540 ;
  LAYER VI3 ;
  RECT 563.760 5.940 563.960 6.140 ;
  LAYER VI3 ;
  RECT 563.360 6.340 563.560 6.540 ;
  LAYER VI3 ;
  RECT 563.360 5.940 563.560 6.140 ;
  LAYER VI3 ;
  RECT 562.960 6.340 563.160 6.540 ;
  LAYER VI3 ;
  RECT 562.960 5.940 563.160 6.140 ;
  LAYER VI3 ;
  RECT 562.560 6.340 562.760 6.540 ;
  LAYER VI3 ;
  RECT 562.560 5.940 562.760 6.140 ;
  LAYER VI3 ;
  RECT 562.160 6.340 562.360 6.540 ;
  LAYER VI3 ;
  RECT 562.160 5.940 562.360 6.140 ;
  LAYER VI3 ;
  RECT 561.760 6.340 561.960 6.540 ;
  LAYER VI3 ;
  RECT 561.760 5.940 561.960 6.140 ;
  LAYER VI3 ;
  RECT 561.360 6.340 561.560 6.540 ;
  LAYER VI3 ;
  RECT 561.360 5.940 561.560 6.140 ;
  LAYER VI3 ;
  RECT 560.960 6.340 561.160 6.540 ;
  LAYER VI3 ;
  RECT 560.960 5.940 561.160 6.140 ;
  LAYER VI3 ;
  RECT 560.560 6.340 560.760 6.540 ;
  LAYER VI3 ;
  RECT 560.560 5.940 560.760 6.140 ;
  LAYER VI3 ;
  RECT 560.160 6.340 560.360 6.540 ;
  LAYER VI3 ;
  RECT 560.160 5.940 560.360 6.140 ;
  LAYER VI3 ;
  RECT 581.240 5.880 589.240 6.740 ;
  LAYER VI3 ;
  RECT 588.840 6.340 589.040 6.540 ;
  LAYER VI3 ;
  RECT 588.840 5.940 589.040 6.140 ;
  LAYER VI3 ;
  RECT 588.440 6.340 588.640 6.540 ;
  LAYER VI3 ;
  RECT 588.440 5.940 588.640 6.140 ;
  LAYER VI3 ;
  RECT 588.040 6.340 588.240 6.540 ;
  LAYER VI3 ;
  RECT 588.040 5.940 588.240 6.140 ;
  LAYER VI3 ;
  RECT 587.640 6.340 587.840 6.540 ;
  LAYER VI3 ;
  RECT 587.640 5.940 587.840 6.140 ;
  LAYER VI3 ;
  RECT 587.240 6.340 587.440 6.540 ;
  LAYER VI3 ;
  RECT 587.240 5.940 587.440 6.140 ;
  LAYER VI3 ;
  RECT 586.840 6.340 587.040 6.540 ;
  LAYER VI3 ;
  RECT 586.840 5.940 587.040 6.140 ;
  LAYER VI3 ;
  RECT 586.440 6.340 586.640 6.540 ;
  LAYER VI3 ;
  RECT 586.440 5.940 586.640 6.140 ;
  LAYER VI3 ;
  RECT 586.040 6.340 586.240 6.540 ;
  LAYER VI3 ;
  RECT 586.040 5.940 586.240 6.140 ;
  LAYER VI3 ;
  RECT 585.640 6.340 585.840 6.540 ;
  LAYER VI3 ;
  RECT 585.640 5.940 585.840 6.140 ;
  LAYER VI3 ;
  RECT 585.240 6.340 585.440 6.540 ;
  LAYER VI3 ;
  RECT 585.240 5.940 585.440 6.140 ;
  LAYER VI3 ;
  RECT 584.840 6.340 585.040 6.540 ;
  LAYER VI3 ;
  RECT 584.840 5.940 585.040 6.140 ;
  LAYER VI3 ;
  RECT 584.440 6.340 584.640 6.540 ;
  LAYER VI3 ;
  RECT 584.440 5.940 584.640 6.140 ;
  LAYER VI3 ;
  RECT 584.040 6.340 584.240 6.540 ;
  LAYER VI3 ;
  RECT 584.040 5.940 584.240 6.140 ;
  LAYER VI3 ;
  RECT 583.640 6.340 583.840 6.540 ;
  LAYER VI3 ;
  RECT 583.640 5.940 583.840 6.140 ;
  LAYER VI3 ;
  RECT 583.240 6.340 583.440 6.540 ;
  LAYER VI3 ;
  RECT 583.240 5.940 583.440 6.140 ;
  LAYER VI3 ;
  RECT 582.840 6.340 583.040 6.540 ;
  LAYER VI3 ;
  RECT 582.840 5.940 583.040 6.140 ;
  LAYER VI3 ;
  RECT 582.440 6.340 582.640 6.540 ;
  LAYER VI3 ;
  RECT 582.440 5.940 582.640 6.140 ;
  LAYER VI3 ;
  RECT 582.040 6.340 582.240 6.540 ;
  LAYER VI3 ;
  RECT 582.040 5.940 582.240 6.140 ;
  LAYER VI3 ;
  RECT 581.640 6.340 581.840 6.540 ;
  LAYER VI3 ;
  RECT 581.640 5.940 581.840 6.140 ;
  LAYER VI3 ;
  RECT 581.240 6.340 581.440 6.540 ;
  LAYER VI3 ;
  RECT 581.240 5.940 581.440 6.140 ;
  LAYER VI3 ;
  RECT 601.080 5.880 609.080 6.740 ;
  LAYER VI3 ;
  RECT 608.680 6.340 608.880 6.540 ;
  LAYER VI3 ;
  RECT 608.680 5.940 608.880 6.140 ;
  LAYER VI3 ;
  RECT 608.280 6.340 608.480 6.540 ;
  LAYER VI3 ;
  RECT 608.280 5.940 608.480 6.140 ;
  LAYER VI3 ;
  RECT 607.880 6.340 608.080 6.540 ;
  LAYER VI3 ;
  RECT 607.880 5.940 608.080 6.140 ;
  LAYER VI3 ;
  RECT 607.480 6.340 607.680 6.540 ;
  LAYER VI3 ;
  RECT 607.480 5.940 607.680 6.140 ;
  LAYER VI3 ;
  RECT 607.080 6.340 607.280 6.540 ;
  LAYER VI3 ;
  RECT 607.080 5.940 607.280 6.140 ;
  LAYER VI3 ;
  RECT 606.680 6.340 606.880 6.540 ;
  LAYER VI3 ;
  RECT 606.680 5.940 606.880 6.140 ;
  LAYER VI3 ;
  RECT 606.280 6.340 606.480 6.540 ;
  LAYER VI3 ;
  RECT 606.280 5.940 606.480 6.140 ;
  LAYER VI3 ;
  RECT 605.880 6.340 606.080 6.540 ;
  LAYER VI3 ;
  RECT 605.880 5.940 606.080 6.140 ;
  LAYER VI3 ;
  RECT 605.480 6.340 605.680 6.540 ;
  LAYER VI3 ;
  RECT 605.480 5.940 605.680 6.140 ;
  LAYER VI3 ;
  RECT 605.080 6.340 605.280 6.540 ;
  LAYER VI3 ;
  RECT 605.080 5.940 605.280 6.140 ;
  LAYER VI3 ;
  RECT 604.680 6.340 604.880 6.540 ;
  LAYER VI3 ;
  RECT 604.680 5.940 604.880 6.140 ;
  LAYER VI3 ;
  RECT 604.280 6.340 604.480 6.540 ;
  LAYER VI3 ;
  RECT 604.280 5.940 604.480 6.140 ;
  LAYER VI3 ;
  RECT 603.880 6.340 604.080 6.540 ;
  LAYER VI3 ;
  RECT 603.880 5.940 604.080 6.140 ;
  LAYER VI3 ;
  RECT 603.480 6.340 603.680 6.540 ;
  LAYER VI3 ;
  RECT 603.480 5.940 603.680 6.140 ;
  LAYER VI3 ;
  RECT 603.080 6.340 603.280 6.540 ;
  LAYER VI3 ;
  RECT 603.080 5.940 603.280 6.140 ;
  LAYER VI3 ;
  RECT 602.680 6.340 602.880 6.540 ;
  LAYER VI3 ;
  RECT 602.680 5.940 602.880 6.140 ;
  LAYER VI3 ;
  RECT 602.280 6.340 602.480 6.540 ;
  LAYER VI3 ;
  RECT 602.280 5.940 602.480 6.140 ;
  LAYER VI3 ;
  RECT 601.880 6.340 602.080 6.540 ;
  LAYER VI3 ;
  RECT 601.880 5.940 602.080 6.140 ;
  LAYER VI3 ;
  RECT 601.480 6.340 601.680 6.540 ;
  LAYER VI3 ;
  RECT 601.480 5.940 601.680 6.140 ;
  LAYER VI3 ;
  RECT 601.080 6.340 601.280 6.540 ;
  LAYER VI3 ;
  RECT 601.080 5.940 601.280 6.140 ;
  LAYER VI3 ;
  RECT 622.160 5.880 630.160 6.740 ;
  LAYER VI3 ;
  RECT 629.760 6.340 629.960 6.540 ;
  LAYER VI3 ;
  RECT 629.760 5.940 629.960 6.140 ;
  LAYER VI3 ;
  RECT 629.360 6.340 629.560 6.540 ;
  LAYER VI3 ;
  RECT 629.360 5.940 629.560 6.140 ;
  LAYER VI3 ;
  RECT 628.960 6.340 629.160 6.540 ;
  LAYER VI3 ;
  RECT 628.960 5.940 629.160 6.140 ;
  LAYER VI3 ;
  RECT 628.560 6.340 628.760 6.540 ;
  LAYER VI3 ;
  RECT 628.560 5.940 628.760 6.140 ;
  LAYER VI3 ;
  RECT 628.160 6.340 628.360 6.540 ;
  LAYER VI3 ;
  RECT 628.160 5.940 628.360 6.140 ;
  LAYER VI3 ;
  RECT 627.760 6.340 627.960 6.540 ;
  LAYER VI3 ;
  RECT 627.760 5.940 627.960 6.140 ;
  LAYER VI3 ;
  RECT 627.360 6.340 627.560 6.540 ;
  LAYER VI3 ;
  RECT 627.360 5.940 627.560 6.140 ;
  LAYER VI3 ;
  RECT 626.960 6.340 627.160 6.540 ;
  LAYER VI3 ;
  RECT 626.960 5.940 627.160 6.140 ;
  LAYER VI3 ;
  RECT 626.560 6.340 626.760 6.540 ;
  LAYER VI3 ;
  RECT 626.560 5.940 626.760 6.140 ;
  LAYER VI3 ;
  RECT 626.160 6.340 626.360 6.540 ;
  LAYER VI3 ;
  RECT 626.160 5.940 626.360 6.140 ;
  LAYER VI3 ;
  RECT 625.760 6.340 625.960 6.540 ;
  LAYER VI3 ;
  RECT 625.760 5.940 625.960 6.140 ;
  LAYER VI3 ;
  RECT 625.360 6.340 625.560 6.540 ;
  LAYER VI3 ;
  RECT 625.360 5.940 625.560 6.140 ;
  LAYER VI3 ;
  RECT 624.960 6.340 625.160 6.540 ;
  LAYER VI3 ;
  RECT 624.960 5.940 625.160 6.140 ;
  LAYER VI3 ;
  RECT 624.560 6.340 624.760 6.540 ;
  LAYER VI3 ;
  RECT 624.560 5.940 624.760 6.140 ;
  LAYER VI3 ;
  RECT 624.160 6.340 624.360 6.540 ;
  LAYER VI3 ;
  RECT 624.160 5.940 624.360 6.140 ;
  LAYER VI3 ;
  RECT 623.760 6.340 623.960 6.540 ;
  LAYER VI3 ;
  RECT 623.760 5.940 623.960 6.140 ;
  LAYER VI3 ;
  RECT 623.360 6.340 623.560 6.540 ;
  LAYER VI3 ;
  RECT 623.360 5.940 623.560 6.140 ;
  LAYER VI3 ;
  RECT 622.960 6.340 623.160 6.540 ;
  LAYER VI3 ;
  RECT 622.960 5.940 623.160 6.140 ;
  LAYER VI3 ;
  RECT 622.560 6.340 622.760 6.540 ;
  LAYER VI3 ;
  RECT 622.560 5.940 622.760 6.140 ;
  LAYER VI3 ;
  RECT 622.160 6.340 622.360 6.540 ;
  LAYER VI3 ;
  RECT 622.160 5.940 622.360 6.140 ;
  LAYER VI3 ;
  RECT 642.000 5.880 650.000 6.740 ;
  LAYER VI3 ;
  RECT 649.600 6.340 649.800 6.540 ;
  LAYER VI3 ;
  RECT 649.600 5.940 649.800 6.140 ;
  LAYER VI3 ;
  RECT 649.200 6.340 649.400 6.540 ;
  LAYER VI3 ;
  RECT 649.200 5.940 649.400 6.140 ;
  LAYER VI3 ;
  RECT 648.800 6.340 649.000 6.540 ;
  LAYER VI3 ;
  RECT 648.800 5.940 649.000 6.140 ;
  LAYER VI3 ;
  RECT 648.400 6.340 648.600 6.540 ;
  LAYER VI3 ;
  RECT 648.400 5.940 648.600 6.140 ;
  LAYER VI3 ;
  RECT 648.000 6.340 648.200 6.540 ;
  LAYER VI3 ;
  RECT 648.000 5.940 648.200 6.140 ;
  LAYER VI3 ;
  RECT 647.600 6.340 647.800 6.540 ;
  LAYER VI3 ;
  RECT 647.600 5.940 647.800 6.140 ;
  LAYER VI3 ;
  RECT 647.200 6.340 647.400 6.540 ;
  LAYER VI3 ;
  RECT 647.200 5.940 647.400 6.140 ;
  LAYER VI3 ;
  RECT 646.800 6.340 647.000 6.540 ;
  LAYER VI3 ;
  RECT 646.800 5.940 647.000 6.140 ;
  LAYER VI3 ;
  RECT 646.400 6.340 646.600 6.540 ;
  LAYER VI3 ;
  RECT 646.400 5.940 646.600 6.140 ;
  LAYER VI3 ;
  RECT 646.000 6.340 646.200 6.540 ;
  LAYER VI3 ;
  RECT 646.000 5.940 646.200 6.140 ;
  LAYER VI3 ;
  RECT 645.600 6.340 645.800 6.540 ;
  LAYER VI3 ;
  RECT 645.600 5.940 645.800 6.140 ;
  LAYER VI3 ;
  RECT 645.200 6.340 645.400 6.540 ;
  LAYER VI3 ;
  RECT 645.200 5.940 645.400 6.140 ;
  LAYER VI3 ;
  RECT 644.800 6.340 645.000 6.540 ;
  LAYER VI3 ;
  RECT 644.800 5.940 645.000 6.140 ;
  LAYER VI3 ;
  RECT 644.400 6.340 644.600 6.540 ;
  LAYER VI3 ;
  RECT 644.400 5.940 644.600 6.140 ;
  LAYER VI3 ;
  RECT 644.000 6.340 644.200 6.540 ;
  LAYER VI3 ;
  RECT 644.000 5.940 644.200 6.140 ;
  LAYER VI3 ;
  RECT 643.600 6.340 643.800 6.540 ;
  LAYER VI3 ;
  RECT 643.600 5.940 643.800 6.140 ;
  LAYER VI3 ;
  RECT 643.200 6.340 643.400 6.540 ;
  LAYER VI3 ;
  RECT 643.200 5.940 643.400 6.140 ;
  LAYER VI3 ;
  RECT 642.800 6.340 643.000 6.540 ;
  LAYER VI3 ;
  RECT 642.800 5.940 643.000 6.140 ;
  LAYER VI3 ;
  RECT 642.400 6.340 642.600 6.540 ;
  LAYER VI3 ;
  RECT 642.400 5.940 642.600 6.140 ;
  LAYER VI3 ;
  RECT 642.000 6.340 642.200 6.540 ;
  LAYER VI3 ;
  RECT 642.000 5.940 642.200 6.140 ;
  LAYER VI3 ;
  RECT 663.080 5.880 671.080 6.740 ;
  LAYER VI3 ;
  RECT 670.680 6.340 670.880 6.540 ;
  LAYER VI3 ;
  RECT 670.680 5.940 670.880 6.140 ;
  LAYER VI3 ;
  RECT 670.280 6.340 670.480 6.540 ;
  LAYER VI3 ;
  RECT 670.280 5.940 670.480 6.140 ;
  LAYER VI3 ;
  RECT 669.880 6.340 670.080 6.540 ;
  LAYER VI3 ;
  RECT 669.880 5.940 670.080 6.140 ;
  LAYER VI3 ;
  RECT 669.480 6.340 669.680 6.540 ;
  LAYER VI3 ;
  RECT 669.480 5.940 669.680 6.140 ;
  LAYER VI3 ;
  RECT 669.080 6.340 669.280 6.540 ;
  LAYER VI3 ;
  RECT 669.080 5.940 669.280 6.140 ;
  LAYER VI3 ;
  RECT 668.680 6.340 668.880 6.540 ;
  LAYER VI3 ;
  RECT 668.680 5.940 668.880 6.140 ;
  LAYER VI3 ;
  RECT 668.280 6.340 668.480 6.540 ;
  LAYER VI3 ;
  RECT 668.280 5.940 668.480 6.140 ;
  LAYER VI3 ;
  RECT 667.880 6.340 668.080 6.540 ;
  LAYER VI3 ;
  RECT 667.880 5.940 668.080 6.140 ;
  LAYER VI3 ;
  RECT 667.480 6.340 667.680 6.540 ;
  LAYER VI3 ;
  RECT 667.480 5.940 667.680 6.140 ;
  LAYER VI3 ;
  RECT 667.080 6.340 667.280 6.540 ;
  LAYER VI3 ;
  RECT 667.080 5.940 667.280 6.140 ;
  LAYER VI3 ;
  RECT 666.680 6.340 666.880 6.540 ;
  LAYER VI3 ;
  RECT 666.680 5.940 666.880 6.140 ;
  LAYER VI3 ;
  RECT 666.280 6.340 666.480 6.540 ;
  LAYER VI3 ;
  RECT 666.280 5.940 666.480 6.140 ;
  LAYER VI3 ;
  RECT 665.880 6.340 666.080 6.540 ;
  LAYER VI3 ;
  RECT 665.880 5.940 666.080 6.140 ;
  LAYER VI3 ;
  RECT 665.480 6.340 665.680 6.540 ;
  LAYER VI3 ;
  RECT 665.480 5.940 665.680 6.140 ;
  LAYER VI3 ;
  RECT 665.080 6.340 665.280 6.540 ;
  LAYER VI3 ;
  RECT 665.080 5.940 665.280 6.140 ;
  LAYER VI3 ;
  RECT 664.680 6.340 664.880 6.540 ;
  LAYER VI3 ;
  RECT 664.680 5.940 664.880 6.140 ;
  LAYER VI3 ;
  RECT 664.280 6.340 664.480 6.540 ;
  LAYER VI3 ;
  RECT 664.280 5.940 664.480 6.140 ;
  LAYER VI3 ;
  RECT 663.880 6.340 664.080 6.540 ;
  LAYER VI3 ;
  RECT 663.880 5.940 664.080 6.140 ;
  LAYER VI3 ;
  RECT 663.480 6.340 663.680 6.540 ;
  LAYER VI3 ;
  RECT 663.480 5.940 663.680 6.140 ;
  LAYER VI3 ;
  RECT 663.080 6.340 663.280 6.540 ;
  LAYER VI3 ;
  RECT 663.080 5.940 663.280 6.140 ;
  LAYER VI3 ;
  RECT 682.920 5.880 690.920 6.740 ;
  LAYER VI3 ;
  RECT 690.520 6.340 690.720 6.540 ;
  LAYER VI3 ;
  RECT 690.520 5.940 690.720 6.140 ;
  LAYER VI3 ;
  RECT 690.120 6.340 690.320 6.540 ;
  LAYER VI3 ;
  RECT 690.120 5.940 690.320 6.140 ;
  LAYER VI3 ;
  RECT 689.720 6.340 689.920 6.540 ;
  LAYER VI3 ;
  RECT 689.720 5.940 689.920 6.140 ;
  LAYER VI3 ;
  RECT 689.320 6.340 689.520 6.540 ;
  LAYER VI3 ;
  RECT 689.320 5.940 689.520 6.140 ;
  LAYER VI3 ;
  RECT 688.920 6.340 689.120 6.540 ;
  LAYER VI3 ;
  RECT 688.920 5.940 689.120 6.140 ;
  LAYER VI3 ;
  RECT 688.520 6.340 688.720 6.540 ;
  LAYER VI3 ;
  RECT 688.520 5.940 688.720 6.140 ;
  LAYER VI3 ;
  RECT 688.120 6.340 688.320 6.540 ;
  LAYER VI3 ;
  RECT 688.120 5.940 688.320 6.140 ;
  LAYER VI3 ;
  RECT 687.720 6.340 687.920 6.540 ;
  LAYER VI3 ;
  RECT 687.720 5.940 687.920 6.140 ;
  LAYER VI3 ;
  RECT 687.320 6.340 687.520 6.540 ;
  LAYER VI3 ;
  RECT 687.320 5.940 687.520 6.140 ;
  LAYER VI3 ;
  RECT 686.920 6.340 687.120 6.540 ;
  LAYER VI3 ;
  RECT 686.920 5.940 687.120 6.140 ;
  LAYER VI3 ;
  RECT 686.520 6.340 686.720 6.540 ;
  LAYER VI3 ;
  RECT 686.520 5.940 686.720 6.140 ;
  LAYER VI3 ;
  RECT 686.120 6.340 686.320 6.540 ;
  LAYER VI3 ;
  RECT 686.120 5.940 686.320 6.140 ;
  LAYER VI3 ;
  RECT 685.720 6.340 685.920 6.540 ;
  LAYER VI3 ;
  RECT 685.720 5.940 685.920 6.140 ;
  LAYER VI3 ;
  RECT 685.320 6.340 685.520 6.540 ;
  LAYER VI3 ;
  RECT 685.320 5.940 685.520 6.140 ;
  LAYER VI3 ;
  RECT 684.920 6.340 685.120 6.540 ;
  LAYER VI3 ;
  RECT 684.920 5.940 685.120 6.140 ;
  LAYER VI3 ;
  RECT 684.520 6.340 684.720 6.540 ;
  LAYER VI3 ;
  RECT 684.520 5.940 684.720 6.140 ;
  LAYER VI3 ;
  RECT 684.120 6.340 684.320 6.540 ;
  LAYER VI3 ;
  RECT 684.120 5.940 684.320 6.140 ;
  LAYER VI3 ;
  RECT 683.720 6.340 683.920 6.540 ;
  LAYER VI3 ;
  RECT 683.720 5.940 683.920 6.140 ;
  LAYER VI3 ;
  RECT 683.320 6.340 683.520 6.540 ;
  LAYER VI3 ;
  RECT 683.320 5.940 683.520 6.140 ;
  LAYER VI3 ;
  RECT 682.920 6.340 683.120 6.540 ;
  LAYER VI3 ;
  RECT 682.920 5.940 683.120 6.140 ;
  LAYER VI3 ;
  RECT 704.000 5.880 712.000 6.740 ;
  LAYER VI3 ;
  RECT 711.600 6.340 711.800 6.540 ;
  LAYER VI3 ;
  RECT 711.600 5.940 711.800 6.140 ;
  LAYER VI3 ;
  RECT 711.200 6.340 711.400 6.540 ;
  LAYER VI3 ;
  RECT 711.200 5.940 711.400 6.140 ;
  LAYER VI3 ;
  RECT 710.800 6.340 711.000 6.540 ;
  LAYER VI3 ;
  RECT 710.800 5.940 711.000 6.140 ;
  LAYER VI3 ;
  RECT 710.400 6.340 710.600 6.540 ;
  LAYER VI3 ;
  RECT 710.400 5.940 710.600 6.140 ;
  LAYER VI3 ;
  RECT 710.000 6.340 710.200 6.540 ;
  LAYER VI3 ;
  RECT 710.000 5.940 710.200 6.140 ;
  LAYER VI3 ;
  RECT 709.600 6.340 709.800 6.540 ;
  LAYER VI3 ;
  RECT 709.600 5.940 709.800 6.140 ;
  LAYER VI3 ;
  RECT 709.200 6.340 709.400 6.540 ;
  LAYER VI3 ;
  RECT 709.200 5.940 709.400 6.140 ;
  LAYER VI3 ;
  RECT 708.800 6.340 709.000 6.540 ;
  LAYER VI3 ;
  RECT 708.800 5.940 709.000 6.140 ;
  LAYER VI3 ;
  RECT 708.400 6.340 708.600 6.540 ;
  LAYER VI3 ;
  RECT 708.400 5.940 708.600 6.140 ;
  LAYER VI3 ;
  RECT 708.000 6.340 708.200 6.540 ;
  LAYER VI3 ;
  RECT 708.000 5.940 708.200 6.140 ;
  LAYER VI3 ;
  RECT 707.600 6.340 707.800 6.540 ;
  LAYER VI3 ;
  RECT 707.600 5.940 707.800 6.140 ;
  LAYER VI3 ;
  RECT 707.200 6.340 707.400 6.540 ;
  LAYER VI3 ;
  RECT 707.200 5.940 707.400 6.140 ;
  LAYER VI3 ;
  RECT 706.800 6.340 707.000 6.540 ;
  LAYER VI3 ;
  RECT 706.800 5.940 707.000 6.140 ;
  LAYER VI3 ;
  RECT 706.400 6.340 706.600 6.540 ;
  LAYER VI3 ;
  RECT 706.400 5.940 706.600 6.140 ;
  LAYER VI3 ;
  RECT 706.000 6.340 706.200 6.540 ;
  LAYER VI3 ;
  RECT 706.000 5.940 706.200 6.140 ;
  LAYER VI3 ;
  RECT 705.600 6.340 705.800 6.540 ;
  LAYER VI3 ;
  RECT 705.600 5.940 705.800 6.140 ;
  LAYER VI3 ;
  RECT 705.200 6.340 705.400 6.540 ;
  LAYER VI3 ;
  RECT 705.200 5.940 705.400 6.140 ;
  LAYER VI3 ;
  RECT 704.800 6.340 705.000 6.540 ;
  LAYER VI3 ;
  RECT 704.800 5.940 705.000 6.140 ;
  LAYER VI3 ;
  RECT 704.400 6.340 704.600 6.540 ;
  LAYER VI3 ;
  RECT 704.400 5.940 704.600 6.140 ;
  LAYER VI3 ;
  RECT 704.000 6.340 704.200 6.540 ;
  LAYER VI3 ;
  RECT 704.000 5.940 704.200 6.140 ;
  LAYER VI3 ;
  RECT 723.840 5.880 731.840 6.740 ;
  LAYER VI3 ;
  RECT 731.440 6.340 731.640 6.540 ;
  LAYER VI3 ;
  RECT 731.440 5.940 731.640 6.140 ;
  LAYER VI3 ;
  RECT 731.040 6.340 731.240 6.540 ;
  LAYER VI3 ;
  RECT 731.040 5.940 731.240 6.140 ;
  LAYER VI3 ;
  RECT 730.640 6.340 730.840 6.540 ;
  LAYER VI3 ;
  RECT 730.640 5.940 730.840 6.140 ;
  LAYER VI3 ;
  RECT 730.240 6.340 730.440 6.540 ;
  LAYER VI3 ;
  RECT 730.240 5.940 730.440 6.140 ;
  LAYER VI3 ;
  RECT 729.840 6.340 730.040 6.540 ;
  LAYER VI3 ;
  RECT 729.840 5.940 730.040 6.140 ;
  LAYER VI3 ;
  RECT 729.440 6.340 729.640 6.540 ;
  LAYER VI3 ;
  RECT 729.440 5.940 729.640 6.140 ;
  LAYER VI3 ;
  RECT 729.040 6.340 729.240 6.540 ;
  LAYER VI3 ;
  RECT 729.040 5.940 729.240 6.140 ;
  LAYER VI3 ;
  RECT 728.640 6.340 728.840 6.540 ;
  LAYER VI3 ;
  RECT 728.640 5.940 728.840 6.140 ;
  LAYER VI3 ;
  RECT 728.240 6.340 728.440 6.540 ;
  LAYER VI3 ;
  RECT 728.240 5.940 728.440 6.140 ;
  LAYER VI3 ;
  RECT 727.840 6.340 728.040 6.540 ;
  LAYER VI3 ;
  RECT 727.840 5.940 728.040 6.140 ;
  LAYER VI3 ;
  RECT 727.440 6.340 727.640 6.540 ;
  LAYER VI3 ;
  RECT 727.440 5.940 727.640 6.140 ;
  LAYER VI3 ;
  RECT 727.040 6.340 727.240 6.540 ;
  LAYER VI3 ;
  RECT 727.040 5.940 727.240 6.140 ;
  LAYER VI3 ;
  RECT 726.640 6.340 726.840 6.540 ;
  LAYER VI3 ;
  RECT 726.640 5.940 726.840 6.140 ;
  LAYER VI3 ;
  RECT 726.240 6.340 726.440 6.540 ;
  LAYER VI3 ;
  RECT 726.240 5.940 726.440 6.140 ;
  LAYER VI3 ;
  RECT 725.840 6.340 726.040 6.540 ;
  LAYER VI3 ;
  RECT 725.840 5.940 726.040 6.140 ;
  LAYER VI3 ;
  RECT 725.440 6.340 725.640 6.540 ;
  LAYER VI3 ;
  RECT 725.440 5.940 725.640 6.140 ;
  LAYER VI3 ;
  RECT 725.040 6.340 725.240 6.540 ;
  LAYER VI3 ;
  RECT 725.040 5.940 725.240 6.140 ;
  LAYER VI3 ;
  RECT 724.640 6.340 724.840 6.540 ;
  LAYER VI3 ;
  RECT 724.640 5.940 724.840 6.140 ;
  LAYER VI3 ;
  RECT 724.240 6.340 724.440 6.540 ;
  LAYER VI3 ;
  RECT 724.240 5.940 724.440 6.140 ;
  LAYER VI3 ;
  RECT 723.840 6.340 724.040 6.540 ;
  LAYER VI3 ;
  RECT 723.840 5.940 724.040 6.140 ;
  LAYER VI3 ;
  RECT 744.920 5.880 752.920 6.740 ;
  LAYER VI3 ;
  RECT 752.520 6.340 752.720 6.540 ;
  LAYER VI3 ;
  RECT 752.520 5.940 752.720 6.140 ;
  LAYER VI3 ;
  RECT 752.120 6.340 752.320 6.540 ;
  LAYER VI3 ;
  RECT 752.120 5.940 752.320 6.140 ;
  LAYER VI3 ;
  RECT 751.720 6.340 751.920 6.540 ;
  LAYER VI3 ;
  RECT 751.720 5.940 751.920 6.140 ;
  LAYER VI3 ;
  RECT 751.320 6.340 751.520 6.540 ;
  LAYER VI3 ;
  RECT 751.320 5.940 751.520 6.140 ;
  LAYER VI3 ;
  RECT 750.920 6.340 751.120 6.540 ;
  LAYER VI3 ;
  RECT 750.920 5.940 751.120 6.140 ;
  LAYER VI3 ;
  RECT 750.520 6.340 750.720 6.540 ;
  LAYER VI3 ;
  RECT 750.520 5.940 750.720 6.140 ;
  LAYER VI3 ;
  RECT 750.120 6.340 750.320 6.540 ;
  LAYER VI3 ;
  RECT 750.120 5.940 750.320 6.140 ;
  LAYER VI3 ;
  RECT 749.720 6.340 749.920 6.540 ;
  LAYER VI3 ;
  RECT 749.720 5.940 749.920 6.140 ;
  LAYER VI3 ;
  RECT 749.320 6.340 749.520 6.540 ;
  LAYER VI3 ;
  RECT 749.320 5.940 749.520 6.140 ;
  LAYER VI3 ;
  RECT 748.920 6.340 749.120 6.540 ;
  LAYER VI3 ;
  RECT 748.920 5.940 749.120 6.140 ;
  LAYER VI3 ;
  RECT 748.520 6.340 748.720 6.540 ;
  LAYER VI3 ;
  RECT 748.520 5.940 748.720 6.140 ;
  LAYER VI3 ;
  RECT 748.120 6.340 748.320 6.540 ;
  LAYER VI3 ;
  RECT 748.120 5.940 748.320 6.140 ;
  LAYER VI3 ;
  RECT 747.720 6.340 747.920 6.540 ;
  LAYER VI3 ;
  RECT 747.720 5.940 747.920 6.140 ;
  LAYER VI3 ;
  RECT 747.320 6.340 747.520 6.540 ;
  LAYER VI3 ;
  RECT 747.320 5.940 747.520 6.140 ;
  LAYER VI3 ;
  RECT 746.920 6.340 747.120 6.540 ;
  LAYER VI3 ;
  RECT 746.920 5.940 747.120 6.140 ;
  LAYER VI3 ;
  RECT 746.520 6.340 746.720 6.540 ;
  LAYER VI3 ;
  RECT 746.520 5.940 746.720 6.140 ;
  LAYER VI3 ;
  RECT 746.120 6.340 746.320 6.540 ;
  LAYER VI3 ;
  RECT 746.120 5.940 746.320 6.140 ;
  LAYER VI3 ;
  RECT 745.720 6.340 745.920 6.540 ;
  LAYER VI3 ;
  RECT 745.720 5.940 745.920 6.140 ;
  LAYER VI3 ;
  RECT 745.320 6.340 745.520 6.540 ;
  LAYER VI3 ;
  RECT 745.320 5.940 745.520 6.140 ;
  LAYER VI3 ;
  RECT 744.920 6.340 745.120 6.540 ;
  LAYER VI3 ;
  RECT 744.920 5.940 745.120 6.140 ;
  LAYER VI3 ;
  RECT 764.760 5.880 772.760 6.740 ;
  LAYER VI3 ;
  RECT 772.360 6.340 772.560 6.540 ;
  LAYER VI3 ;
  RECT 772.360 5.940 772.560 6.140 ;
  LAYER VI3 ;
  RECT 771.960 6.340 772.160 6.540 ;
  LAYER VI3 ;
  RECT 771.960 5.940 772.160 6.140 ;
  LAYER VI3 ;
  RECT 771.560 6.340 771.760 6.540 ;
  LAYER VI3 ;
  RECT 771.560 5.940 771.760 6.140 ;
  LAYER VI3 ;
  RECT 771.160 6.340 771.360 6.540 ;
  LAYER VI3 ;
  RECT 771.160 5.940 771.360 6.140 ;
  LAYER VI3 ;
  RECT 770.760 6.340 770.960 6.540 ;
  LAYER VI3 ;
  RECT 770.760 5.940 770.960 6.140 ;
  LAYER VI3 ;
  RECT 770.360 6.340 770.560 6.540 ;
  LAYER VI3 ;
  RECT 770.360 5.940 770.560 6.140 ;
  LAYER VI3 ;
  RECT 769.960 6.340 770.160 6.540 ;
  LAYER VI3 ;
  RECT 769.960 5.940 770.160 6.140 ;
  LAYER VI3 ;
  RECT 769.560 6.340 769.760 6.540 ;
  LAYER VI3 ;
  RECT 769.560 5.940 769.760 6.140 ;
  LAYER VI3 ;
  RECT 769.160 6.340 769.360 6.540 ;
  LAYER VI3 ;
  RECT 769.160 5.940 769.360 6.140 ;
  LAYER VI3 ;
  RECT 768.760 6.340 768.960 6.540 ;
  LAYER VI3 ;
  RECT 768.760 5.940 768.960 6.140 ;
  LAYER VI3 ;
  RECT 768.360 6.340 768.560 6.540 ;
  LAYER VI3 ;
  RECT 768.360 5.940 768.560 6.140 ;
  LAYER VI3 ;
  RECT 767.960 6.340 768.160 6.540 ;
  LAYER VI3 ;
  RECT 767.960 5.940 768.160 6.140 ;
  LAYER VI3 ;
  RECT 767.560 6.340 767.760 6.540 ;
  LAYER VI3 ;
  RECT 767.560 5.940 767.760 6.140 ;
  LAYER VI3 ;
  RECT 767.160 6.340 767.360 6.540 ;
  LAYER VI3 ;
  RECT 767.160 5.940 767.360 6.140 ;
  LAYER VI3 ;
  RECT 766.760 6.340 766.960 6.540 ;
  LAYER VI3 ;
  RECT 766.760 5.940 766.960 6.140 ;
  LAYER VI3 ;
  RECT 766.360 6.340 766.560 6.540 ;
  LAYER VI3 ;
  RECT 766.360 5.940 766.560 6.140 ;
  LAYER VI3 ;
  RECT 765.960 6.340 766.160 6.540 ;
  LAYER VI3 ;
  RECT 765.960 5.940 766.160 6.140 ;
  LAYER VI3 ;
  RECT 765.560 6.340 765.760 6.540 ;
  LAYER VI3 ;
  RECT 765.560 5.940 765.760 6.140 ;
  LAYER VI3 ;
  RECT 765.160 6.340 765.360 6.540 ;
  LAYER VI3 ;
  RECT 765.160 5.940 765.360 6.140 ;
  LAYER VI3 ;
  RECT 764.760 6.340 764.960 6.540 ;
  LAYER VI3 ;
  RECT 764.760 5.940 764.960 6.140 ;
  LAYER VI3 ;
  RECT 785.840 5.880 793.840 6.740 ;
  LAYER VI3 ;
  RECT 793.440 6.340 793.640 6.540 ;
  LAYER VI3 ;
  RECT 793.440 5.940 793.640 6.140 ;
  LAYER VI3 ;
  RECT 793.040 6.340 793.240 6.540 ;
  LAYER VI3 ;
  RECT 793.040 5.940 793.240 6.140 ;
  LAYER VI3 ;
  RECT 792.640 6.340 792.840 6.540 ;
  LAYER VI3 ;
  RECT 792.640 5.940 792.840 6.140 ;
  LAYER VI3 ;
  RECT 792.240 6.340 792.440 6.540 ;
  LAYER VI3 ;
  RECT 792.240 5.940 792.440 6.140 ;
  LAYER VI3 ;
  RECT 791.840 6.340 792.040 6.540 ;
  LAYER VI3 ;
  RECT 791.840 5.940 792.040 6.140 ;
  LAYER VI3 ;
  RECT 791.440 6.340 791.640 6.540 ;
  LAYER VI3 ;
  RECT 791.440 5.940 791.640 6.140 ;
  LAYER VI3 ;
  RECT 791.040 6.340 791.240 6.540 ;
  LAYER VI3 ;
  RECT 791.040 5.940 791.240 6.140 ;
  LAYER VI3 ;
  RECT 790.640 6.340 790.840 6.540 ;
  LAYER VI3 ;
  RECT 790.640 5.940 790.840 6.140 ;
  LAYER VI3 ;
  RECT 790.240 6.340 790.440 6.540 ;
  LAYER VI3 ;
  RECT 790.240 5.940 790.440 6.140 ;
  LAYER VI3 ;
  RECT 789.840 6.340 790.040 6.540 ;
  LAYER VI3 ;
  RECT 789.840 5.940 790.040 6.140 ;
  LAYER VI3 ;
  RECT 789.440 6.340 789.640 6.540 ;
  LAYER VI3 ;
  RECT 789.440 5.940 789.640 6.140 ;
  LAYER VI3 ;
  RECT 789.040 6.340 789.240 6.540 ;
  LAYER VI3 ;
  RECT 789.040 5.940 789.240 6.140 ;
  LAYER VI3 ;
  RECT 788.640 6.340 788.840 6.540 ;
  LAYER VI3 ;
  RECT 788.640 5.940 788.840 6.140 ;
  LAYER VI3 ;
  RECT 788.240 6.340 788.440 6.540 ;
  LAYER VI3 ;
  RECT 788.240 5.940 788.440 6.140 ;
  LAYER VI3 ;
  RECT 787.840 6.340 788.040 6.540 ;
  LAYER VI3 ;
  RECT 787.840 5.940 788.040 6.140 ;
  LAYER VI3 ;
  RECT 787.440 6.340 787.640 6.540 ;
  LAYER VI3 ;
  RECT 787.440 5.940 787.640 6.140 ;
  LAYER VI3 ;
  RECT 787.040 6.340 787.240 6.540 ;
  LAYER VI3 ;
  RECT 787.040 5.940 787.240 6.140 ;
  LAYER VI3 ;
  RECT 786.640 6.340 786.840 6.540 ;
  LAYER VI3 ;
  RECT 786.640 5.940 786.840 6.140 ;
  LAYER VI3 ;
  RECT 786.240 6.340 786.440 6.540 ;
  LAYER VI3 ;
  RECT 786.240 5.940 786.440 6.140 ;
  LAYER VI3 ;
  RECT 785.840 6.340 786.040 6.540 ;
  LAYER VI3 ;
  RECT 785.840 5.940 786.040 6.140 ;
  LAYER VI3 ;
  RECT 805.680 5.880 813.680 6.740 ;
  LAYER VI3 ;
  RECT 813.280 6.340 813.480 6.540 ;
  LAYER VI3 ;
  RECT 813.280 5.940 813.480 6.140 ;
  LAYER VI3 ;
  RECT 812.880 6.340 813.080 6.540 ;
  LAYER VI3 ;
  RECT 812.880 5.940 813.080 6.140 ;
  LAYER VI3 ;
  RECT 812.480 6.340 812.680 6.540 ;
  LAYER VI3 ;
  RECT 812.480 5.940 812.680 6.140 ;
  LAYER VI3 ;
  RECT 812.080 6.340 812.280 6.540 ;
  LAYER VI3 ;
  RECT 812.080 5.940 812.280 6.140 ;
  LAYER VI3 ;
  RECT 811.680 6.340 811.880 6.540 ;
  LAYER VI3 ;
  RECT 811.680 5.940 811.880 6.140 ;
  LAYER VI3 ;
  RECT 811.280 6.340 811.480 6.540 ;
  LAYER VI3 ;
  RECT 811.280 5.940 811.480 6.140 ;
  LAYER VI3 ;
  RECT 810.880 6.340 811.080 6.540 ;
  LAYER VI3 ;
  RECT 810.880 5.940 811.080 6.140 ;
  LAYER VI3 ;
  RECT 810.480 6.340 810.680 6.540 ;
  LAYER VI3 ;
  RECT 810.480 5.940 810.680 6.140 ;
  LAYER VI3 ;
  RECT 810.080 6.340 810.280 6.540 ;
  LAYER VI3 ;
  RECT 810.080 5.940 810.280 6.140 ;
  LAYER VI3 ;
  RECT 809.680 6.340 809.880 6.540 ;
  LAYER VI3 ;
  RECT 809.680 5.940 809.880 6.140 ;
  LAYER VI3 ;
  RECT 809.280 6.340 809.480 6.540 ;
  LAYER VI3 ;
  RECT 809.280 5.940 809.480 6.140 ;
  LAYER VI3 ;
  RECT 808.880 6.340 809.080 6.540 ;
  LAYER VI3 ;
  RECT 808.880 5.940 809.080 6.140 ;
  LAYER VI3 ;
  RECT 808.480 6.340 808.680 6.540 ;
  LAYER VI3 ;
  RECT 808.480 5.940 808.680 6.140 ;
  LAYER VI3 ;
  RECT 808.080 6.340 808.280 6.540 ;
  LAYER VI3 ;
  RECT 808.080 5.940 808.280 6.140 ;
  LAYER VI3 ;
  RECT 807.680 6.340 807.880 6.540 ;
  LAYER VI3 ;
  RECT 807.680 5.940 807.880 6.140 ;
  LAYER VI3 ;
  RECT 807.280 6.340 807.480 6.540 ;
  LAYER VI3 ;
  RECT 807.280 5.940 807.480 6.140 ;
  LAYER VI3 ;
  RECT 806.880 6.340 807.080 6.540 ;
  LAYER VI3 ;
  RECT 806.880 5.940 807.080 6.140 ;
  LAYER VI3 ;
  RECT 806.480 6.340 806.680 6.540 ;
  LAYER VI3 ;
  RECT 806.480 5.940 806.680 6.140 ;
  LAYER VI3 ;
  RECT 806.080 6.340 806.280 6.540 ;
  LAYER VI3 ;
  RECT 806.080 5.940 806.280 6.140 ;
  LAYER VI3 ;
  RECT 805.680 6.340 805.880 6.540 ;
  LAYER VI3 ;
  RECT 805.680 5.940 805.880 6.140 ;
  LAYER VI3 ;
  RECT 826.760 5.880 834.760 6.740 ;
  LAYER VI3 ;
  RECT 834.360 6.340 834.560 6.540 ;
  LAYER VI3 ;
  RECT 834.360 5.940 834.560 6.140 ;
  LAYER VI3 ;
  RECT 833.960 6.340 834.160 6.540 ;
  LAYER VI3 ;
  RECT 833.960 5.940 834.160 6.140 ;
  LAYER VI3 ;
  RECT 833.560 6.340 833.760 6.540 ;
  LAYER VI3 ;
  RECT 833.560 5.940 833.760 6.140 ;
  LAYER VI3 ;
  RECT 833.160 6.340 833.360 6.540 ;
  LAYER VI3 ;
  RECT 833.160 5.940 833.360 6.140 ;
  LAYER VI3 ;
  RECT 832.760 6.340 832.960 6.540 ;
  LAYER VI3 ;
  RECT 832.760 5.940 832.960 6.140 ;
  LAYER VI3 ;
  RECT 832.360 6.340 832.560 6.540 ;
  LAYER VI3 ;
  RECT 832.360 5.940 832.560 6.140 ;
  LAYER VI3 ;
  RECT 831.960 6.340 832.160 6.540 ;
  LAYER VI3 ;
  RECT 831.960 5.940 832.160 6.140 ;
  LAYER VI3 ;
  RECT 831.560 6.340 831.760 6.540 ;
  LAYER VI3 ;
  RECT 831.560 5.940 831.760 6.140 ;
  LAYER VI3 ;
  RECT 831.160 6.340 831.360 6.540 ;
  LAYER VI3 ;
  RECT 831.160 5.940 831.360 6.140 ;
  LAYER VI3 ;
  RECT 830.760 6.340 830.960 6.540 ;
  LAYER VI3 ;
  RECT 830.760 5.940 830.960 6.140 ;
  LAYER VI3 ;
  RECT 830.360 6.340 830.560 6.540 ;
  LAYER VI3 ;
  RECT 830.360 5.940 830.560 6.140 ;
  LAYER VI3 ;
  RECT 829.960 6.340 830.160 6.540 ;
  LAYER VI3 ;
  RECT 829.960 5.940 830.160 6.140 ;
  LAYER VI3 ;
  RECT 829.560 6.340 829.760 6.540 ;
  LAYER VI3 ;
  RECT 829.560 5.940 829.760 6.140 ;
  LAYER VI3 ;
  RECT 829.160 6.340 829.360 6.540 ;
  LAYER VI3 ;
  RECT 829.160 5.940 829.360 6.140 ;
  LAYER VI3 ;
  RECT 828.760 6.340 828.960 6.540 ;
  LAYER VI3 ;
  RECT 828.760 5.940 828.960 6.140 ;
  LAYER VI3 ;
  RECT 828.360 6.340 828.560 6.540 ;
  LAYER VI3 ;
  RECT 828.360 5.940 828.560 6.140 ;
  LAYER VI3 ;
  RECT 827.960 6.340 828.160 6.540 ;
  LAYER VI3 ;
  RECT 827.960 5.940 828.160 6.140 ;
  LAYER VI3 ;
  RECT 827.560 6.340 827.760 6.540 ;
  LAYER VI3 ;
  RECT 827.560 5.940 827.760 6.140 ;
  LAYER VI3 ;
  RECT 827.160 6.340 827.360 6.540 ;
  LAYER VI3 ;
  RECT 827.160 5.940 827.360 6.140 ;
  LAYER VI3 ;
  RECT 826.760 6.340 826.960 6.540 ;
  LAYER VI3 ;
  RECT 826.760 5.940 826.960 6.140 ;
  LAYER VI3 ;
  RECT 846.600 5.880 854.600 6.740 ;
  LAYER VI3 ;
  RECT 854.200 6.340 854.400 6.540 ;
  LAYER VI3 ;
  RECT 854.200 5.940 854.400 6.140 ;
  LAYER VI3 ;
  RECT 853.800 6.340 854.000 6.540 ;
  LAYER VI3 ;
  RECT 853.800 5.940 854.000 6.140 ;
  LAYER VI3 ;
  RECT 853.400 6.340 853.600 6.540 ;
  LAYER VI3 ;
  RECT 853.400 5.940 853.600 6.140 ;
  LAYER VI3 ;
  RECT 853.000 6.340 853.200 6.540 ;
  LAYER VI3 ;
  RECT 853.000 5.940 853.200 6.140 ;
  LAYER VI3 ;
  RECT 852.600 6.340 852.800 6.540 ;
  LAYER VI3 ;
  RECT 852.600 5.940 852.800 6.140 ;
  LAYER VI3 ;
  RECT 852.200 6.340 852.400 6.540 ;
  LAYER VI3 ;
  RECT 852.200 5.940 852.400 6.140 ;
  LAYER VI3 ;
  RECT 851.800 6.340 852.000 6.540 ;
  LAYER VI3 ;
  RECT 851.800 5.940 852.000 6.140 ;
  LAYER VI3 ;
  RECT 851.400 6.340 851.600 6.540 ;
  LAYER VI3 ;
  RECT 851.400 5.940 851.600 6.140 ;
  LAYER VI3 ;
  RECT 851.000 6.340 851.200 6.540 ;
  LAYER VI3 ;
  RECT 851.000 5.940 851.200 6.140 ;
  LAYER VI3 ;
  RECT 850.600 6.340 850.800 6.540 ;
  LAYER VI3 ;
  RECT 850.600 5.940 850.800 6.140 ;
  LAYER VI3 ;
  RECT 850.200 6.340 850.400 6.540 ;
  LAYER VI3 ;
  RECT 850.200 5.940 850.400 6.140 ;
  LAYER VI3 ;
  RECT 849.800 6.340 850.000 6.540 ;
  LAYER VI3 ;
  RECT 849.800 5.940 850.000 6.140 ;
  LAYER VI3 ;
  RECT 849.400 6.340 849.600 6.540 ;
  LAYER VI3 ;
  RECT 849.400 5.940 849.600 6.140 ;
  LAYER VI3 ;
  RECT 849.000 6.340 849.200 6.540 ;
  LAYER VI3 ;
  RECT 849.000 5.940 849.200 6.140 ;
  LAYER VI3 ;
  RECT 848.600 6.340 848.800 6.540 ;
  LAYER VI3 ;
  RECT 848.600 5.940 848.800 6.140 ;
  LAYER VI3 ;
  RECT 848.200 6.340 848.400 6.540 ;
  LAYER VI3 ;
  RECT 848.200 5.940 848.400 6.140 ;
  LAYER VI3 ;
  RECT 847.800 6.340 848.000 6.540 ;
  LAYER VI3 ;
  RECT 847.800 5.940 848.000 6.140 ;
  LAYER VI3 ;
  RECT 847.400 6.340 847.600 6.540 ;
  LAYER VI3 ;
  RECT 847.400 5.940 847.600 6.140 ;
  LAYER VI3 ;
  RECT 847.000 6.340 847.200 6.540 ;
  LAYER VI3 ;
  RECT 847.000 5.940 847.200 6.140 ;
  LAYER VI3 ;
  RECT 846.600 6.340 846.800 6.540 ;
  LAYER VI3 ;
  RECT 846.600 5.940 846.800 6.140 ;
  LAYER VI3 ;
  RECT 867.680 5.880 875.680 6.740 ;
  LAYER VI3 ;
  RECT 875.280 6.340 875.480 6.540 ;
  LAYER VI3 ;
  RECT 875.280 5.940 875.480 6.140 ;
  LAYER VI3 ;
  RECT 874.880 6.340 875.080 6.540 ;
  LAYER VI3 ;
  RECT 874.880 5.940 875.080 6.140 ;
  LAYER VI3 ;
  RECT 874.480 6.340 874.680 6.540 ;
  LAYER VI3 ;
  RECT 874.480 5.940 874.680 6.140 ;
  LAYER VI3 ;
  RECT 874.080 6.340 874.280 6.540 ;
  LAYER VI3 ;
  RECT 874.080 5.940 874.280 6.140 ;
  LAYER VI3 ;
  RECT 873.680 6.340 873.880 6.540 ;
  LAYER VI3 ;
  RECT 873.680 5.940 873.880 6.140 ;
  LAYER VI3 ;
  RECT 873.280 6.340 873.480 6.540 ;
  LAYER VI3 ;
  RECT 873.280 5.940 873.480 6.140 ;
  LAYER VI3 ;
  RECT 872.880 6.340 873.080 6.540 ;
  LAYER VI3 ;
  RECT 872.880 5.940 873.080 6.140 ;
  LAYER VI3 ;
  RECT 872.480 6.340 872.680 6.540 ;
  LAYER VI3 ;
  RECT 872.480 5.940 872.680 6.140 ;
  LAYER VI3 ;
  RECT 872.080 6.340 872.280 6.540 ;
  LAYER VI3 ;
  RECT 872.080 5.940 872.280 6.140 ;
  LAYER VI3 ;
  RECT 871.680 6.340 871.880 6.540 ;
  LAYER VI3 ;
  RECT 871.680 5.940 871.880 6.140 ;
  LAYER VI3 ;
  RECT 871.280 6.340 871.480 6.540 ;
  LAYER VI3 ;
  RECT 871.280 5.940 871.480 6.140 ;
  LAYER VI3 ;
  RECT 870.880 6.340 871.080 6.540 ;
  LAYER VI3 ;
  RECT 870.880 5.940 871.080 6.140 ;
  LAYER VI3 ;
  RECT 870.480 6.340 870.680 6.540 ;
  LAYER VI3 ;
  RECT 870.480 5.940 870.680 6.140 ;
  LAYER VI3 ;
  RECT 870.080 6.340 870.280 6.540 ;
  LAYER VI3 ;
  RECT 870.080 5.940 870.280 6.140 ;
  LAYER VI3 ;
  RECT 869.680 6.340 869.880 6.540 ;
  LAYER VI3 ;
  RECT 869.680 5.940 869.880 6.140 ;
  LAYER VI3 ;
  RECT 869.280 6.340 869.480 6.540 ;
  LAYER VI3 ;
  RECT 869.280 5.940 869.480 6.140 ;
  LAYER VI3 ;
  RECT 868.880 6.340 869.080 6.540 ;
  LAYER VI3 ;
  RECT 868.880 5.940 869.080 6.140 ;
  LAYER VI3 ;
  RECT 868.480 6.340 868.680 6.540 ;
  LAYER VI3 ;
  RECT 868.480 5.940 868.680 6.140 ;
  LAYER VI3 ;
  RECT 868.080 6.340 868.280 6.540 ;
  LAYER VI3 ;
  RECT 868.080 5.940 868.280 6.140 ;
  LAYER VI3 ;
  RECT 867.680 6.340 867.880 6.540 ;
  LAYER VI3 ;
  RECT 867.680 5.940 867.880 6.140 ;
  LAYER VI3 ;
  RECT 887.520 5.880 895.520 6.740 ;
  LAYER VI3 ;
  RECT 895.120 6.340 895.320 6.540 ;
  LAYER VI3 ;
  RECT 895.120 5.940 895.320 6.140 ;
  LAYER VI3 ;
  RECT 894.720 6.340 894.920 6.540 ;
  LAYER VI3 ;
  RECT 894.720 5.940 894.920 6.140 ;
  LAYER VI3 ;
  RECT 894.320 6.340 894.520 6.540 ;
  LAYER VI3 ;
  RECT 894.320 5.940 894.520 6.140 ;
  LAYER VI3 ;
  RECT 893.920 6.340 894.120 6.540 ;
  LAYER VI3 ;
  RECT 893.920 5.940 894.120 6.140 ;
  LAYER VI3 ;
  RECT 893.520 6.340 893.720 6.540 ;
  LAYER VI3 ;
  RECT 893.520 5.940 893.720 6.140 ;
  LAYER VI3 ;
  RECT 893.120 6.340 893.320 6.540 ;
  LAYER VI3 ;
  RECT 893.120 5.940 893.320 6.140 ;
  LAYER VI3 ;
  RECT 892.720 6.340 892.920 6.540 ;
  LAYER VI3 ;
  RECT 892.720 5.940 892.920 6.140 ;
  LAYER VI3 ;
  RECT 892.320 6.340 892.520 6.540 ;
  LAYER VI3 ;
  RECT 892.320 5.940 892.520 6.140 ;
  LAYER VI3 ;
  RECT 891.920 6.340 892.120 6.540 ;
  LAYER VI3 ;
  RECT 891.920 5.940 892.120 6.140 ;
  LAYER VI3 ;
  RECT 891.520 6.340 891.720 6.540 ;
  LAYER VI3 ;
  RECT 891.520 5.940 891.720 6.140 ;
  LAYER VI3 ;
  RECT 891.120 6.340 891.320 6.540 ;
  LAYER VI3 ;
  RECT 891.120 5.940 891.320 6.140 ;
  LAYER VI3 ;
  RECT 890.720 6.340 890.920 6.540 ;
  LAYER VI3 ;
  RECT 890.720 5.940 890.920 6.140 ;
  LAYER VI3 ;
  RECT 890.320 6.340 890.520 6.540 ;
  LAYER VI3 ;
  RECT 890.320 5.940 890.520 6.140 ;
  LAYER VI3 ;
  RECT 889.920 6.340 890.120 6.540 ;
  LAYER VI3 ;
  RECT 889.920 5.940 890.120 6.140 ;
  LAYER VI3 ;
  RECT 889.520 6.340 889.720 6.540 ;
  LAYER VI3 ;
  RECT 889.520 5.940 889.720 6.140 ;
  LAYER VI3 ;
  RECT 889.120 6.340 889.320 6.540 ;
  LAYER VI3 ;
  RECT 889.120 5.940 889.320 6.140 ;
  LAYER VI3 ;
  RECT 888.720 6.340 888.920 6.540 ;
  LAYER VI3 ;
  RECT 888.720 5.940 888.920 6.140 ;
  LAYER VI3 ;
  RECT 888.320 6.340 888.520 6.540 ;
  LAYER VI3 ;
  RECT 888.320 5.940 888.520 6.140 ;
  LAYER VI3 ;
  RECT 887.920 6.340 888.120 6.540 ;
  LAYER VI3 ;
  RECT 887.920 5.940 888.120 6.140 ;
  LAYER VI3 ;
  RECT 887.520 6.340 887.720 6.540 ;
  LAYER VI3 ;
  RECT 887.520 5.940 887.720 6.140 ;
  LAYER VI3 ;
  RECT 908.600 5.880 916.600 6.740 ;
  LAYER VI3 ;
  RECT 916.200 6.340 916.400 6.540 ;
  LAYER VI3 ;
  RECT 916.200 5.940 916.400 6.140 ;
  LAYER VI3 ;
  RECT 915.800 6.340 916.000 6.540 ;
  LAYER VI3 ;
  RECT 915.800 5.940 916.000 6.140 ;
  LAYER VI3 ;
  RECT 915.400 6.340 915.600 6.540 ;
  LAYER VI3 ;
  RECT 915.400 5.940 915.600 6.140 ;
  LAYER VI3 ;
  RECT 915.000 6.340 915.200 6.540 ;
  LAYER VI3 ;
  RECT 915.000 5.940 915.200 6.140 ;
  LAYER VI3 ;
  RECT 914.600 6.340 914.800 6.540 ;
  LAYER VI3 ;
  RECT 914.600 5.940 914.800 6.140 ;
  LAYER VI3 ;
  RECT 914.200 6.340 914.400 6.540 ;
  LAYER VI3 ;
  RECT 914.200 5.940 914.400 6.140 ;
  LAYER VI3 ;
  RECT 913.800 6.340 914.000 6.540 ;
  LAYER VI3 ;
  RECT 913.800 5.940 914.000 6.140 ;
  LAYER VI3 ;
  RECT 913.400 6.340 913.600 6.540 ;
  LAYER VI3 ;
  RECT 913.400 5.940 913.600 6.140 ;
  LAYER VI3 ;
  RECT 913.000 6.340 913.200 6.540 ;
  LAYER VI3 ;
  RECT 913.000 5.940 913.200 6.140 ;
  LAYER VI3 ;
  RECT 912.600 6.340 912.800 6.540 ;
  LAYER VI3 ;
  RECT 912.600 5.940 912.800 6.140 ;
  LAYER VI3 ;
  RECT 912.200 6.340 912.400 6.540 ;
  LAYER VI3 ;
  RECT 912.200 5.940 912.400 6.140 ;
  LAYER VI3 ;
  RECT 911.800 6.340 912.000 6.540 ;
  LAYER VI3 ;
  RECT 911.800 5.940 912.000 6.140 ;
  LAYER VI3 ;
  RECT 911.400 6.340 911.600 6.540 ;
  LAYER VI3 ;
  RECT 911.400 5.940 911.600 6.140 ;
  LAYER VI3 ;
  RECT 911.000 6.340 911.200 6.540 ;
  LAYER VI3 ;
  RECT 911.000 5.940 911.200 6.140 ;
  LAYER VI3 ;
  RECT 910.600 6.340 910.800 6.540 ;
  LAYER VI3 ;
  RECT 910.600 5.940 910.800 6.140 ;
  LAYER VI3 ;
  RECT 910.200 6.340 910.400 6.540 ;
  LAYER VI3 ;
  RECT 910.200 5.940 910.400 6.140 ;
  LAYER VI3 ;
  RECT 909.800 6.340 910.000 6.540 ;
  LAYER VI3 ;
  RECT 909.800 5.940 910.000 6.140 ;
  LAYER VI3 ;
  RECT 909.400 6.340 909.600 6.540 ;
  LAYER VI3 ;
  RECT 909.400 5.940 909.600 6.140 ;
  LAYER VI3 ;
  RECT 909.000 6.340 909.200 6.540 ;
  LAYER VI3 ;
  RECT 909.000 5.940 909.200 6.140 ;
  LAYER VI3 ;
  RECT 908.600 6.340 908.800 6.540 ;
  LAYER VI3 ;
  RECT 908.600 5.940 908.800 6.140 ;
  LAYER VI3 ;
  RECT 928.440 5.880 936.440 6.740 ;
  LAYER VI3 ;
  RECT 936.040 6.340 936.240 6.540 ;
  LAYER VI3 ;
  RECT 936.040 5.940 936.240 6.140 ;
  LAYER VI3 ;
  RECT 935.640 6.340 935.840 6.540 ;
  LAYER VI3 ;
  RECT 935.640 5.940 935.840 6.140 ;
  LAYER VI3 ;
  RECT 935.240 6.340 935.440 6.540 ;
  LAYER VI3 ;
  RECT 935.240 5.940 935.440 6.140 ;
  LAYER VI3 ;
  RECT 934.840 6.340 935.040 6.540 ;
  LAYER VI3 ;
  RECT 934.840 5.940 935.040 6.140 ;
  LAYER VI3 ;
  RECT 934.440 6.340 934.640 6.540 ;
  LAYER VI3 ;
  RECT 934.440 5.940 934.640 6.140 ;
  LAYER VI3 ;
  RECT 934.040 6.340 934.240 6.540 ;
  LAYER VI3 ;
  RECT 934.040 5.940 934.240 6.140 ;
  LAYER VI3 ;
  RECT 933.640 6.340 933.840 6.540 ;
  LAYER VI3 ;
  RECT 933.640 5.940 933.840 6.140 ;
  LAYER VI3 ;
  RECT 933.240 6.340 933.440 6.540 ;
  LAYER VI3 ;
  RECT 933.240 5.940 933.440 6.140 ;
  LAYER VI3 ;
  RECT 932.840 6.340 933.040 6.540 ;
  LAYER VI3 ;
  RECT 932.840 5.940 933.040 6.140 ;
  LAYER VI3 ;
  RECT 932.440 6.340 932.640 6.540 ;
  LAYER VI3 ;
  RECT 932.440 5.940 932.640 6.140 ;
  LAYER VI3 ;
  RECT 932.040 6.340 932.240 6.540 ;
  LAYER VI3 ;
  RECT 932.040 5.940 932.240 6.140 ;
  LAYER VI3 ;
  RECT 931.640 6.340 931.840 6.540 ;
  LAYER VI3 ;
  RECT 931.640 5.940 931.840 6.140 ;
  LAYER VI3 ;
  RECT 931.240 6.340 931.440 6.540 ;
  LAYER VI3 ;
  RECT 931.240 5.940 931.440 6.140 ;
  LAYER VI3 ;
  RECT 930.840 6.340 931.040 6.540 ;
  LAYER VI3 ;
  RECT 930.840 5.940 931.040 6.140 ;
  LAYER VI3 ;
  RECT 930.440 6.340 930.640 6.540 ;
  LAYER VI3 ;
  RECT 930.440 5.940 930.640 6.140 ;
  LAYER VI3 ;
  RECT 930.040 6.340 930.240 6.540 ;
  LAYER VI3 ;
  RECT 930.040 5.940 930.240 6.140 ;
  LAYER VI3 ;
  RECT 929.640 6.340 929.840 6.540 ;
  LAYER VI3 ;
  RECT 929.640 5.940 929.840 6.140 ;
  LAYER VI3 ;
  RECT 929.240 6.340 929.440 6.540 ;
  LAYER VI3 ;
  RECT 929.240 5.940 929.440 6.140 ;
  LAYER VI3 ;
  RECT 928.840 6.340 929.040 6.540 ;
  LAYER VI3 ;
  RECT 928.840 5.940 929.040 6.140 ;
  LAYER VI3 ;
  RECT 928.440 6.340 928.640 6.540 ;
  LAYER VI3 ;
  RECT 928.440 5.940 928.640 6.140 ;
  LAYER VI3 ;
  RECT 949.520 5.880 957.520 6.740 ;
  LAYER VI3 ;
  RECT 957.120 6.340 957.320 6.540 ;
  LAYER VI3 ;
  RECT 957.120 5.940 957.320 6.140 ;
  LAYER VI3 ;
  RECT 956.720 6.340 956.920 6.540 ;
  LAYER VI3 ;
  RECT 956.720 5.940 956.920 6.140 ;
  LAYER VI3 ;
  RECT 956.320 6.340 956.520 6.540 ;
  LAYER VI3 ;
  RECT 956.320 5.940 956.520 6.140 ;
  LAYER VI3 ;
  RECT 955.920 6.340 956.120 6.540 ;
  LAYER VI3 ;
  RECT 955.920 5.940 956.120 6.140 ;
  LAYER VI3 ;
  RECT 955.520 6.340 955.720 6.540 ;
  LAYER VI3 ;
  RECT 955.520 5.940 955.720 6.140 ;
  LAYER VI3 ;
  RECT 955.120 6.340 955.320 6.540 ;
  LAYER VI3 ;
  RECT 955.120 5.940 955.320 6.140 ;
  LAYER VI3 ;
  RECT 954.720 6.340 954.920 6.540 ;
  LAYER VI3 ;
  RECT 954.720 5.940 954.920 6.140 ;
  LAYER VI3 ;
  RECT 954.320 6.340 954.520 6.540 ;
  LAYER VI3 ;
  RECT 954.320 5.940 954.520 6.140 ;
  LAYER VI3 ;
  RECT 953.920 6.340 954.120 6.540 ;
  LAYER VI3 ;
  RECT 953.920 5.940 954.120 6.140 ;
  LAYER VI3 ;
  RECT 953.520 6.340 953.720 6.540 ;
  LAYER VI3 ;
  RECT 953.520 5.940 953.720 6.140 ;
  LAYER VI3 ;
  RECT 953.120 6.340 953.320 6.540 ;
  LAYER VI3 ;
  RECT 953.120 5.940 953.320 6.140 ;
  LAYER VI3 ;
  RECT 952.720 6.340 952.920 6.540 ;
  LAYER VI3 ;
  RECT 952.720 5.940 952.920 6.140 ;
  LAYER VI3 ;
  RECT 952.320 6.340 952.520 6.540 ;
  LAYER VI3 ;
  RECT 952.320 5.940 952.520 6.140 ;
  LAYER VI3 ;
  RECT 951.920 6.340 952.120 6.540 ;
  LAYER VI3 ;
  RECT 951.920 5.940 952.120 6.140 ;
  LAYER VI3 ;
  RECT 951.520 6.340 951.720 6.540 ;
  LAYER VI3 ;
  RECT 951.520 5.940 951.720 6.140 ;
  LAYER VI3 ;
  RECT 951.120 6.340 951.320 6.540 ;
  LAYER VI3 ;
  RECT 951.120 5.940 951.320 6.140 ;
  LAYER VI3 ;
  RECT 950.720 6.340 950.920 6.540 ;
  LAYER VI3 ;
  RECT 950.720 5.940 950.920 6.140 ;
  LAYER VI3 ;
  RECT 950.320 6.340 950.520 6.540 ;
  LAYER VI3 ;
  RECT 950.320 5.940 950.520 6.140 ;
  LAYER VI3 ;
  RECT 949.920 6.340 950.120 6.540 ;
  LAYER VI3 ;
  RECT 949.920 5.940 950.120 6.140 ;
  LAYER VI3 ;
  RECT 949.520 6.340 949.720 6.540 ;
  LAYER VI3 ;
  RECT 949.520 5.940 949.720 6.140 ;
  LAYER VI3 ;
  RECT 969.360 5.880 977.360 6.740 ;
  LAYER VI3 ;
  RECT 976.960 6.340 977.160 6.540 ;
  LAYER VI3 ;
  RECT 976.960 5.940 977.160 6.140 ;
  LAYER VI3 ;
  RECT 976.560 6.340 976.760 6.540 ;
  LAYER VI3 ;
  RECT 976.560 5.940 976.760 6.140 ;
  LAYER VI3 ;
  RECT 976.160 6.340 976.360 6.540 ;
  LAYER VI3 ;
  RECT 976.160 5.940 976.360 6.140 ;
  LAYER VI3 ;
  RECT 975.760 6.340 975.960 6.540 ;
  LAYER VI3 ;
  RECT 975.760 5.940 975.960 6.140 ;
  LAYER VI3 ;
  RECT 975.360 6.340 975.560 6.540 ;
  LAYER VI3 ;
  RECT 975.360 5.940 975.560 6.140 ;
  LAYER VI3 ;
  RECT 974.960 6.340 975.160 6.540 ;
  LAYER VI3 ;
  RECT 974.960 5.940 975.160 6.140 ;
  LAYER VI3 ;
  RECT 974.560 6.340 974.760 6.540 ;
  LAYER VI3 ;
  RECT 974.560 5.940 974.760 6.140 ;
  LAYER VI3 ;
  RECT 974.160 6.340 974.360 6.540 ;
  LAYER VI3 ;
  RECT 974.160 5.940 974.360 6.140 ;
  LAYER VI3 ;
  RECT 973.760 6.340 973.960 6.540 ;
  LAYER VI3 ;
  RECT 973.760 5.940 973.960 6.140 ;
  LAYER VI3 ;
  RECT 973.360 6.340 973.560 6.540 ;
  LAYER VI3 ;
  RECT 973.360 5.940 973.560 6.140 ;
  LAYER VI3 ;
  RECT 972.960 6.340 973.160 6.540 ;
  LAYER VI3 ;
  RECT 972.960 5.940 973.160 6.140 ;
  LAYER VI3 ;
  RECT 972.560 6.340 972.760 6.540 ;
  LAYER VI3 ;
  RECT 972.560 5.940 972.760 6.140 ;
  LAYER VI3 ;
  RECT 972.160 6.340 972.360 6.540 ;
  LAYER VI3 ;
  RECT 972.160 5.940 972.360 6.140 ;
  LAYER VI3 ;
  RECT 971.760 6.340 971.960 6.540 ;
  LAYER VI3 ;
  RECT 971.760 5.940 971.960 6.140 ;
  LAYER VI3 ;
  RECT 971.360 6.340 971.560 6.540 ;
  LAYER VI3 ;
  RECT 971.360 5.940 971.560 6.140 ;
  LAYER VI3 ;
  RECT 970.960 6.340 971.160 6.540 ;
  LAYER VI3 ;
  RECT 970.960 5.940 971.160 6.140 ;
  LAYER VI3 ;
  RECT 970.560 6.340 970.760 6.540 ;
  LAYER VI3 ;
  RECT 970.560 5.940 970.760 6.140 ;
  LAYER VI3 ;
  RECT 970.160 6.340 970.360 6.540 ;
  LAYER VI3 ;
  RECT 970.160 5.940 970.360 6.140 ;
  LAYER VI3 ;
  RECT 969.760 6.340 969.960 6.540 ;
  LAYER VI3 ;
  RECT 969.760 5.940 969.960 6.140 ;
  LAYER VI3 ;
  RECT 969.360 6.340 969.560 6.540 ;
  LAYER VI3 ;
  RECT 969.360 5.940 969.560 6.140 ;
  LAYER VI3 ;
  RECT 990.440 5.880 998.440 6.740 ;
  LAYER VI3 ;
  RECT 998.040 6.340 998.240 6.540 ;
  LAYER VI3 ;
  RECT 998.040 5.940 998.240 6.140 ;
  LAYER VI3 ;
  RECT 997.640 6.340 997.840 6.540 ;
  LAYER VI3 ;
  RECT 997.640 5.940 997.840 6.140 ;
  LAYER VI3 ;
  RECT 997.240 6.340 997.440 6.540 ;
  LAYER VI3 ;
  RECT 997.240 5.940 997.440 6.140 ;
  LAYER VI3 ;
  RECT 996.840 6.340 997.040 6.540 ;
  LAYER VI3 ;
  RECT 996.840 5.940 997.040 6.140 ;
  LAYER VI3 ;
  RECT 996.440 6.340 996.640 6.540 ;
  LAYER VI3 ;
  RECT 996.440 5.940 996.640 6.140 ;
  LAYER VI3 ;
  RECT 996.040 6.340 996.240 6.540 ;
  LAYER VI3 ;
  RECT 996.040 5.940 996.240 6.140 ;
  LAYER VI3 ;
  RECT 995.640 6.340 995.840 6.540 ;
  LAYER VI3 ;
  RECT 995.640 5.940 995.840 6.140 ;
  LAYER VI3 ;
  RECT 995.240 6.340 995.440 6.540 ;
  LAYER VI3 ;
  RECT 995.240 5.940 995.440 6.140 ;
  LAYER VI3 ;
  RECT 994.840 6.340 995.040 6.540 ;
  LAYER VI3 ;
  RECT 994.840 5.940 995.040 6.140 ;
  LAYER VI3 ;
  RECT 994.440 6.340 994.640 6.540 ;
  LAYER VI3 ;
  RECT 994.440 5.940 994.640 6.140 ;
  LAYER VI3 ;
  RECT 994.040 6.340 994.240 6.540 ;
  LAYER VI3 ;
  RECT 994.040 5.940 994.240 6.140 ;
  LAYER VI3 ;
  RECT 993.640 6.340 993.840 6.540 ;
  LAYER VI3 ;
  RECT 993.640 5.940 993.840 6.140 ;
  LAYER VI3 ;
  RECT 993.240 6.340 993.440 6.540 ;
  LAYER VI3 ;
  RECT 993.240 5.940 993.440 6.140 ;
  LAYER VI3 ;
  RECT 992.840 6.340 993.040 6.540 ;
  LAYER VI3 ;
  RECT 992.840 5.940 993.040 6.140 ;
  LAYER VI3 ;
  RECT 992.440 6.340 992.640 6.540 ;
  LAYER VI3 ;
  RECT 992.440 5.940 992.640 6.140 ;
  LAYER VI3 ;
  RECT 992.040 6.340 992.240 6.540 ;
  LAYER VI3 ;
  RECT 992.040 5.940 992.240 6.140 ;
  LAYER VI3 ;
  RECT 991.640 6.340 991.840 6.540 ;
  LAYER VI3 ;
  RECT 991.640 5.940 991.840 6.140 ;
  LAYER VI3 ;
  RECT 991.240 6.340 991.440 6.540 ;
  LAYER VI3 ;
  RECT 991.240 5.940 991.440 6.140 ;
  LAYER VI3 ;
  RECT 990.840 6.340 991.040 6.540 ;
  LAYER VI3 ;
  RECT 990.840 5.940 991.040 6.140 ;
  LAYER VI3 ;
  RECT 990.440 6.340 990.640 6.540 ;
  LAYER VI3 ;
  RECT 990.440 5.940 990.640 6.140 ;
  LAYER VI3 ;
  RECT 1010.280 5.880 1018.280 6.740 ;
  LAYER VI3 ;
  RECT 1017.880 6.340 1018.080 6.540 ;
  LAYER VI3 ;
  RECT 1017.880 5.940 1018.080 6.140 ;
  LAYER VI3 ;
  RECT 1017.480 6.340 1017.680 6.540 ;
  LAYER VI3 ;
  RECT 1017.480 5.940 1017.680 6.140 ;
  LAYER VI3 ;
  RECT 1017.080 6.340 1017.280 6.540 ;
  LAYER VI3 ;
  RECT 1017.080 5.940 1017.280 6.140 ;
  LAYER VI3 ;
  RECT 1016.680 6.340 1016.880 6.540 ;
  LAYER VI3 ;
  RECT 1016.680 5.940 1016.880 6.140 ;
  LAYER VI3 ;
  RECT 1016.280 6.340 1016.480 6.540 ;
  LAYER VI3 ;
  RECT 1016.280 5.940 1016.480 6.140 ;
  LAYER VI3 ;
  RECT 1015.880 6.340 1016.080 6.540 ;
  LAYER VI3 ;
  RECT 1015.880 5.940 1016.080 6.140 ;
  LAYER VI3 ;
  RECT 1015.480 6.340 1015.680 6.540 ;
  LAYER VI3 ;
  RECT 1015.480 5.940 1015.680 6.140 ;
  LAYER VI3 ;
  RECT 1015.080 6.340 1015.280 6.540 ;
  LAYER VI3 ;
  RECT 1015.080 5.940 1015.280 6.140 ;
  LAYER VI3 ;
  RECT 1014.680 6.340 1014.880 6.540 ;
  LAYER VI3 ;
  RECT 1014.680 5.940 1014.880 6.140 ;
  LAYER VI3 ;
  RECT 1014.280 6.340 1014.480 6.540 ;
  LAYER VI3 ;
  RECT 1014.280 5.940 1014.480 6.140 ;
  LAYER VI3 ;
  RECT 1013.880 6.340 1014.080 6.540 ;
  LAYER VI3 ;
  RECT 1013.880 5.940 1014.080 6.140 ;
  LAYER VI3 ;
  RECT 1013.480 6.340 1013.680 6.540 ;
  LAYER VI3 ;
  RECT 1013.480 5.940 1013.680 6.140 ;
  LAYER VI3 ;
  RECT 1013.080 6.340 1013.280 6.540 ;
  LAYER VI3 ;
  RECT 1013.080 5.940 1013.280 6.140 ;
  LAYER VI3 ;
  RECT 1012.680 6.340 1012.880 6.540 ;
  LAYER VI3 ;
  RECT 1012.680 5.940 1012.880 6.140 ;
  LAYER VI3 ;
  RECT 1012.280 6.340 1012.480 6.540 ;
  LAYER VI3 ;
  RECT 1012.280 5.940 1012.480 6.140 ;
  LAYER VI3 ;
  RECT 1011.880 6.340 1012.080 6.540 ;
  LAYER VI3 ;
  RECT 1011.880 5.940 1012.080 6.140 ;
  LAYER VI3 ;
  RECT 1011.480 6.340 1011.680 6.540 ;
  LAYER VI3 ;
  RECT 1011.480 5.940 1011.680 6.140 ;
  LAYER VI3 ;
  RECT 1011.080 6.340 1011.280 6.540 ;
  LAYER VI3 ;
  RECT 1011.080 5.940 1011.280 6.140 ;
  LAYER VI3 ;
  RECT 1010.680 6.340 1010.880 6.540 ;
  LAYER VI3 ;
  RECT 1010.680 5.940 1010.880 6.140 ;
  LAYER VI3 ;
  RECT 1010.280 6.340 1010.480 6.540 ;
  LAYER VI3 ;
  RECT 1010.280 5.940 1010.480 6.140 ;
  LAYER VI3 ;
  RECT 1031.360 5.880 1039.360 6.740 ;
  LAYER VI3 ;
  RECT 1038.960 6.340 1039.160 6.540 ;
  LAYER VI3 ;
  RECT 1038.960 5.940 1039.160 6.140 ;
  LAYER VI3 ;
  RECT 1038.560 6.340 1038.760 6.540 ;
  LAYER VI3 ;
  RECT 1038.560 5.940 1038.760 6.140 ;
  LAYER VI3 ;
  RECT 1038.160 6.340 1038.360 6.540 ;
  LAYER VI3 ;
  RECT 1038.160 5.940 1038.360 6.140 ;
  LAYER VI3 ;
  RECT 1037.760 6.340 1037.960 6.540 ;
  LAYER VI3 ;
  RECT 1037.760 5.940 1037.960 6.140 ;
  LAYER VI3 ;
  RECT 1037.360 6.340 1037.560 6.540 ;
  LAYER VI3 ;
  RECT 1037.360 5.940 1037.560 6.140 ;
  LAYER VI3 ;
  RECT 1036.960 6.340 1037.160 6.540 ;
  LAYER VI3 ;
  RECT 1036.960 5.940 1037.160 6.140 ;
  LAYER VI3 ;
  RECT 1036.560 6.340 1036.760 6.540 ;
  LAYER VI3 ;
  RECT 1036.560 5.940 1036.760 6.140 ;
  LAYER VI3 ;
  RECT 1036.160 6.340 1036.360 6.540 ;
  LAYER VI3 ;
  RECT 1036.160 5.940 1036.360 6.140 ;
  LAYER VI3 ;
  RECT 1035.760 6.340 1035.960 6.540 ;
  LAYER VI3 ;
  RECT 1035.760 5.940 1035.960 6.140 ;
  LAYER VI3 ;
  RECT 1035.360 6.340 1035.560 6.540 ;
  LAYER VI3 ;
  RECT 1035.360 5.940 1035.560 6.140 ;
  LAYER VI3 ;
  RECT 1034.960 6.340 1035.160 6.540 ;
  LAYER VI3 ;
  RECT 1034.960 5.940 1035.160 6.140 ;
  LAYER VI3 ;
  RECT 1034.560 6.340 1034.760 6.540 ;
  LAYER VI3 ;
  RECT 1034.560 5.940 1034.760 6.140 ;
  LAYER VI3 ;
  RECT 1034.160 6.340 1034.360 6.540 ;
  LAYER VI3 ;
  RECT 1034.160 5.940 1034.360 6.140 ;
  LAYER VI3 ;
  RECT 1033.760 6.340 1033.960 6.540 ;
  LAYER VI3 ;
  RECT 1033.760 5.940 1033.960 6.140 ;
  LAYER VI3 ;
  RECT 1033.360 6.340 1033.560 6.540 ;
  LAYER VI3 ;
  RECT 1033.360 5.940 1033.560 6.140 ;
  LAYER VI3 ;
  RECT 1032.960 6.340 1033.160 6.540 ;
  LAYER VI3 ;
  RECT 1032.960 5.940 1033.160 6.140 ;
  LAYER VI3 ;
  RECT 1032.560 6.340 1032.760 6.540 ;
  LAYER VI3 ;
  RECT 1032.560 5.940 1032.760 6.140 ;
  LAYER VI3 ;
  RECT 1032.160 6.340 1032.360 6.540 ;
  LAYER VI3 ;
  RECT 1032.160 5.940 1032.360 6.140 ;
  LAYER VI3 ;
  RECT 1031.760 6.340 1031.960 6.540 ;
  LAYER VI3 ;
  RECT 1031.760 5.940 1031.960 6.140 ;
  LAYER VI3 ;
  RECT 1031.360 6.340 1031.560 6.540 ;
  LAYER VI3 ;
  RECT 1031.360 5.940 1031.560 6.140 ;
  LAYER VI3 ;
  RECT 1051.200 5.880 1059.200 6.740 ;
  LAYER VI3 ;
  RECT 1058.800 6.340 1059.000 6.540 ;
  LAYER VI3 ;
  RECT 1058.800 5.940 1059.000 6.140 ;
  LAYER VI3 ;
  RECT 1058.400 6.340 1058.600 6.540 ;
  LAYER VI3 ;
  RECT 1058.400 5.940 1058.600 6.140 ;
  LAYER VI3 ;
  RECT 1058.000 6.340 1058.200 6.540 ;
  LAYER VI3 ;
  RECT 1058.000 5.940 1058.200 6.140 ;
  LAYER VI3 ;
  RECT 1057.600 6.340 1057.800 6.540 ;
  LAYER VI3 ;
  RECT 1057.600 5.940 1057.800 6.140 ;
  LAYER VI3 ;
  RECT 1057.200 6.340 1057.400 6.540 ;
  LAYER VI3 ;
  RECT 1057.200 5.940 1057.400 6.140 ;
  LAYER VI3 ;
  RECT 1056.800 6.340 1057.000 6.540 ;
  LAYER VI3 ;
  RECT 1056.800 5.940 1057.000 6.140 ;
  LAYER VI3 ;
  RECT 1056.400 6.340 1056.600 6.540 ;
  LAYER VI3 ;
  RECT 1056.400 5.940 1056.600 6.140 ;
  LAYER VI3 ;
  RECT 1056.000 6.340 1056.200 6.540 ;
  LAYER VI3 ;
  RECT 1056.000 5.940 1056.200 6.140 ;
  LAYER VI3 ;
  RECT 1055.600 6.340 1055.800 6.540 ;
  LAYER VI3 ;
  RECT 1055.600 5.940 1055.800 6.140 ;
  LAYER VI3 ;
  RECT 1055.200 6.340 1055.400 6.540 ;
  LAYER VI3 ;
  RECT 1055.200 5.940 1055.400 6.140 ;
  LAYER VI3 ;
  RECT 1054.800 6.340 1055.000 6.540 ;
  LAYER VI3 ;
  RECT 1054.800 5.940 1055.000 6.140 ;
  LAYER VI3 ;
  RECT 1054.400 6.340 1054.600 6.540 ;
  LAYER VI3 ;
  RECT 1054.400 5.940 1054.600 6.140 ;
  LAYER VI3 ;
  RECT 1054.000 6.340 1054.200 6.540 ;
  LAYER VI3 ;
  RECT 1054.000 5.940 1054.200 6.140 ;
  LAYER VI3 ;
  RECT 1053.600 6.340 1053.800 6.540 ;
  LAYER VI3 ;
  RECT 1053.600 5.940 1053.800 6.140 ;
  LAYER VI3 ;
  RECT 1053.200 6.340 1053.400 6.540 ;
  LAYER VI3 ;
  RECT 1053.200 5.940 1053.400 6.140 ;
  LAYER VI3 ;
  RECT 1052.800 6.340 1053.000 6.540 ;
  LAYER VI3 ;
  RECT 1052.800 5.940 1053.000 6.140 ;
  LAYER VI3 ;
  RECT 1052.400 6.340 1052.600 6.540 ;
  LAYER VI3 ;
  RECT 1052.400 5.940 1052.600 6.140 ;
  LAYER VI3 ;
  RECT 1052.000 6.340 1052.200 6.540 ;
  LAYER VI3 ;
  RECT 1052.000 5.940 1052.200 6.140 ;
  LAYER VI3 ;
  RECT 1051.600 6.340 1051.800 6.540 ;
  LAYER VI3 ;
  RECT 1051.600 5.940 1051.800 6.140 ;
  LAYER VI3 ;
  RECT 1051.200 6.340 1051.400 6.540 ;
  LAYER VI3 ;
  RECT 1051.200 5.940 1051.400 6.140 ;
  LAYER VI3 ;
  RECT 1072.280 5.880 1080.280 6.740 ;
  LAYER VI3 ;
  RECT 1079.880 6.340 1080.080 6.540 ;
  LAYER VI3 ;
  RECT 1079.880 5.940 1080.080 6.140 ;
  LAYER VI3 ;
  RECT 1079.480 6.340 1079.680 6.540 ;
  LAYER VI3 ;
  RECT 1079.480 5.940 1079.680 6.140 ;
  LAYER VI3 ;
  RECT 1079.080 6.340 1079.280 6.540 ;
  LAYER VI3 ;
  RECT 1079.080 5.940 1079.280 6.140 ;
  LAYER VI3 ;
  RECT 1078.680 6.340 1078.880 6.540 ;
  LAYER VI3 ;
  RECT 1078.680 5.940 1078.880 6.140 ;
  LAYER VI3 ;
  RECT 1078.280 6.340 1078.480 6.540 ;
  LAYER VI3 ;
  RECT 1078.280 5.940 1078.480 6.140 ;
  LAYER VI3 ;
  RECT 1077.880 6.340 1078.080 6.540 ;
  LAYER VI3 ;
  RECT 1077.880 5.940 1078.080 6.140 ;
  LAYER VI3 ;
  RECT 1077.480 6.340 1077.680 6.540 ;
  LAYER VI3 ;
  RECT 1077.480 5.940 1077.680 6.140 ;
  LAYER VI3 ;
  RECT 1077.080 6.340 1077.280 6.540 ;
  LAYER VI3 ;
  RECT 1077.080 5.940 1077.280 6.140 ;
  LAYER VI3 ;
  RECT 1076.680 6.340 1076.880 6.540 ;
  LAYER VI3 ;
  RECT 1076.680 5.940 1076.880 6.140 ;
  LAYER VI3 ;
  RECT 1076.280 6.340 1076.480 6.540 ;
  LAYER VI3 ;
  RECT 1076.280 5.940 1076.480 6.140 ;
  LAYER VI3 ;
  RECT 1075.880 6.340 1076.080 6.540 ;
  LAYER VI3 ;
  RECT 1075.880 5.940 1076.080 6.140 ;
  LAYER VI3 ;
  RECT 1075.480 6.340 1075.680 6.540 ;
  LAYER VI3 ;
  RECT 1075.480 5.940 1075.680 6.140 ;
  LAYER VI3 ;
  RECT 1075.080 6.340 1075.280 6.540 ;
  LAYER VI3 ;
  RECT 1075.080 5.940 1075.280 6.140 ;
  LAYER VI3 ;
  RECT 1074.680 6.340 1074.880 6.540 ;
  LAYER VI3 ;
  RECT 1074.680 5.940 1074.880 6.140 ;
  LAYER VI3 ;
  RECT 1074.280 6.340 1074.480 6.540 ;
  LAYER VI3 ;
  RECT 1074.280 5.940 1074.480 6.140 ;
  LAYER VI3 ;
  RECT 1073.880 6.340 1074.080 6.540 ;
  LAYER VI3 ;
  RECT 1073.880 5.940 1074.080 6.140 ;
  LAYER VI3 ;
  RECT 1073.480 6.340 1073.680 6.540 ;
  LAYER VI3 ;
  RECT 1073.480 5.940 1073.680 6.140 ;
  LAYER VI3 ;
  RECT 1073.080 6.340 1073.280 6.540 ;
  LAYER VI3 ;
  RECT 1073.080 5.940 1073.280 6.140 ;
  LAYER VI3 ;
  RECT 1072.680 6.340 1072.880 6.540 ;
  LAYER VI3 ;
  RECT 1072.680 5.940 1072.880 6.140 ;
  LAYER VI3 ;
  RECT 1072.280 6.340 1072.480 6.540 ;
  LAYER VI3 ;
  RECT 1072.280 5.940 1072.480 6.140 ;
  LAYER VI3 ;
  RECT 1092.120 5.880 1100.120 6.740 ;
  LAYER VI3 ;
  RECT 1099.720 6.340 1099.920 6.540 ;
  LAYER VI3 ;
  RECT 1099.720 5.940 1099.920 6.140 ;
  LAYER VI3 ;
  RECT 1099.320 6.340 1099.520 6.540 ;
  LAYER VI3 ;
  RECT 1099.320 5.940 1099.520 6.140 ;
  LAYER VI3 ;
  RECT 1098.920 6.340 1099.120 6.540 ;
  LAYER VI3 ;
  RECT 1098.920 5.940 1099.120 6.140 ;
  LAYER VI3 ;
  RECT 1098.520 6.340 1098.720 6.540 ;
  LAYER VI3 ;
  RECT 1098.520 5.940 1098.720 6.140 ;
  LAYER VI3 ;
  RECT 1098.120 6.340 1098.320 6.540 ;
  LAYER VI3 ;
  RECT 1098.120 5.940 1098.320 6.140 ;
  LAYER VI3 ;
  RECT 1097.720 6.340 1097.920 6.540 ;
  LAYER VI3 ;
  RECT 1097.720 5.940 1097.920 6.140 ;
  LAYER VI3 ;
  RECT 1097.320 6.340 1097.520 6.540 ;
  LAYER VI3 ;
  RECT 1097.320 5.940 1097.520 6.140 ;
  LAYER VI3 ;
  RECT 1096.920 6.340 1097.120 6.540 ;
  LAYER VI3 ;
  RECT 1096.920 5.940 1097.120 6.140 ;
  LAYER VI3 ;
  RECT 1096.520 6.340 1096.720 6.540 ;
  LAYER VI3 ;
  RECT 1096.520 5.940 1096.720 6.140 ;
  LAYER VI3 ;
  RECT 1096.120 6.340 1096.320 6.540 ;
  LAYER VI3 ;
  RECT 1096.120 5.940 1096.320 6.140 ;
  LAYER VI3 ;
  RECT 1095.720 6.340 1095.920 6.540 ;
  LAYER VI3 ;
  RECT 1095.720 5.940 1095.920 6.140 ;
  LAYER VI3 ;
  RECT 1095.320 6.340 1095.520 6.540 ;
  LAYER VI3 ;
  RECT 1095.320 5.940 1095.520 6.140 ;
  LAYER VI3 ;
  RECT 1094.920 6.340 1095.120 6.540 ;
  LAYER VI3 ;
  RECT 1094.920 5.940 1095.120 6.140 ;
  LAYER VI3 ;
  RECT 1094.520 6.340 1094.720 6.540 ;
  LAYER VI3 ;
  RECT 1094.520 5.940 1094.720 6.140 ;
  LAYER VI3 ;
  RECT 1094.120 6.340 1094.320 6.540 ;
  LAYER VI3 ;
  RECT 1094.120 5.940 1094.320 6.140 ;
  LAYER VI3 ;
  RECT 1093.720 6.340 1093.920 6.540 ;
  LAYER VI3 ;
  RECT 1093.720 5.940 1093.920 6.140 ;
  LAYER VI3 ;
  RECT 1093.320 6.340 1093.520 6.540 ;
  LAYER VI3 ;
  RECT 1093.320 5.940 1093.520 6.140 ;
  LAYER VI3 ;
  RECT 1092.920 6.340 1093.120 6.540 ;
  LAYER VI3 ;
  RECT 1092.920 5.940 1093.120 6.140 ;
  LAYER VI3 ;
  RECT 1092.520 6.340 1092.720 6.540 ;
  LAYER VI3 ;
  RECT 1092.520 5.940 1092.720 6.140 ;
  LAYER VI3 ;
  RECT 1092.120 6.340 1092.320 6.540 ;
  LAYER VI3 ;
  RECT 1092.120 5.940 1092.320 6.140 ;
  LAYER VI3 ;
  RECT 1113.200 5.880 1121.200 6.740 ;
  LAYER VI3 ;
  RECT 1120.800 6.340 1121.000 6.540 ;
  LAYER VI3 ;
  RECT 1120.800 5.940 1121.000 6.140 ;
  LAYER VI3 ;
  RECT 1120.400 6.340 1120.600 6.540 ;
  LAYER VI3 ;
  RECT 1120.400 5.940 1120.600 6.140 ;
  LAYER VI3 ;
  RECT 1120.000 6.340 1120.200 6.540 ;
  LAYER VI3 ;
  RECT 1120.000 5.940 1120.200 6.140 ;
  LAYER VI3 ;
  RECT 1119.600 6.340 1119.800 6.540 ;
  LAYER VI3 ;
  RECT 1119.600 5.940 1119.800 6.140 ;
  LAYER VI3 ;
  RECT 1119.200 6.340 1119.400 6.540 ;
  LAYER VI3 ;
  RECT 1119.200 5.940 1119.400 6.140 ;
  LAYER VI3 ;
  RECT 1118.800 6.340 1119.000 6.540 ;
  LAYER VI3 ;
  RECT 1118.800 5.940 1119.000 6.140 ;
  LAYER VI3 ;
  RECT 1118.400 6.340 1118.600 6.540 ;
  LAYER VI3 ;
  RECT 1118.400 5.940 1118.600 6.140 ;
  LAYER VI3 ;
  RECT 1118.000 6.340 1118.200 6.540 ;
  LAYER VI3 ;
  RECT 1118.000 5.940 1118.200 6.140 ;
  LAYER VI3 ;
  RECT 1117.600 6.340 1117.800 6.540 ;
  LAYER VI3 ;
  RECT 1117.600 5.940 1117.800 6.140 ;
  LAYER VI3 ;
  RECT 1117.200 6.340 1117.400 6.540 ;
  LAYER VI3 ;
  RECT 1117.200 5.940 1117.400 6.140 ;
  LAYER VI3 ;
  RECT 1116.800 6.340 1117.000 6.540 ;
  LAYER VI3 ;
  RECT 1116.800 5.940 1117.000 6.140 ;
  LAYER VI3 ;
  RECT 1116.400 6.340 1116.600 6.540 ;
  LAYER VI3 ;
  RECT 1116.400 5.940 1116.600 6.140 ;
  LAYER VI3 ;
  RECT 1116.000 6.340 1116.200 6.540 ;
  LAYER VI3 ;
  RECT 1116.000 5.940 1116.200 6.140 ;
  LAYER VI3 ;
  RECT 1115.600 6.340 1115.800 6.540 ;
  LAYER VI3 ;
  RECT 1115.600 5.940 1115.800 6.140 ;
  LAYER VI3 ;
  RECT 1115.200 6.340 1115.400 6.540 ;
  LAYER VI3 ;
  RECT 1115.200 5.940 1115.400 6.140 ;
  LAYER VI3 ;
  RECT 1114.800 6.340 1115.000 6.540 ;
  LAYER VI3 ;
  RECT 1114.800 5.940 1115.000 6.140 ;
  LAYER VI3 ;
  RECT 1114.400 6.340 1114.600 6.540 ;
  LAYER VI3 ;
  RECT 1114.400 5.940 1114.600 6.140 ;
  LAYER VI3 ;
  RECT 1114.000 6.340 1114.200 6.540 ;
  LAYER VI3 ;
  RECT 1114.000 5.940 1114.200 6.140 ;
  LAYER VI3 ;
  RECT 1113.600 6.340 1113.800 6.540 ;
  LAYER VI3 ;
  RECT 1113.600 5.940 1113.800 6.140 ;
  LAYER VI3 ;
  RECT 1113.200 6.340 1113.400 6.540 ;
  LAYER VI3 ;
  RECT 1113.200 5.940 1113.400 6.140 ;
  LAYER VI3 ;
  RECT 1133.040 5.880 1141.040 6.740 ;
  LAYER VI3 ;
  RECT 1140.640 6.340 1140.840 6.540 ;
  LAYER VI3 ;
  RECT 1140.640 5.940 1140.840 6.140 ;
  LAYER VI3 ;
  RECT 1140.240 6.340 1140.440 6.540 ;
  LAYER VI3 ;
  RECT 1140.240 5.940 1140.440 6.140 ;
  LAYER VI3 ;
  RECT 1139.840 6.340 1140.040 6.540 ;
  LAYER VI3 ;
  RECT 1139.840 5.940 1140.040 6.140 ;
  LAYER VI3 ;
  RECT 1139.440 6.340 1139.640 6.540 ;
  LAYER VI3 ;
  RECT 1139.440 5.940 1139.640 6.140 ;
  LAYER VI3 ;
  RECT 1139.040 6.340 1139.240 6.540 ;
  LAYER VI3 ;
  RECT 1139.040 5.940 1139.240 6.140 ;
  LAYER VI3 ;
  RECT 1138.640 6.340 1138.840 6.540 ;
  LAYER VI3 ;
  RECT 1138.640 5.940 1138.840 6.140 ;
  LAYER VI3 ;
  RECT 1138.240 6.340 1138.440 6.540 ;
  LAYER VI3 ;
  RECT 1138.240 5.940 1138.440 6.140 ;
  LAYER VI3 ;
  RECT 1137.840 6.340 1138.040 6.540 ;
  LAYER VI3 ;
  RECT 1137.840 5.940 1138.040 6.140 ;
  LAYER VI3 ;
  RECT 1137.440 6.340 1137.640 6.540 ;
  LAYER VI3 ;
  RECT 1137.440 5.940 1137.640 6.140 ;
  LAYER VI3 ;
  RECT 1137.040 6.340 1137.240 6.540 ;
  LAYER VI3 ;
  RECT 1137.040 5.940 1137.240 6.140 ;
  LAYER VI3 ;
  RECT 1136.640 6.340 1136.840 6.540 ;
  LAYER VI3 ;
  RECT 1136.640 5.940 1136.840 6.140 ;
  LAYER VI3 ;
  RECT 1136.240 6.340 1136.440 6.540 ;
  LAYER VI3 ;
  RECT 1136.240 5.940 1136.440 6.140 ;
  LAYER VI3 ;
  RECT 1135.840 6.340 1136.040 6.540 ;
  LAYER VI3 ;
  RECT 1135.840 5.940 1136.040 6.140 ;
  LAYER VI3 ;
  RECT 1135.440 6.340 1135.640 6.540 ;
  LAYER VI3 ;
  RECT 1135.440 5.940 1135.640 6.140 ;
  LAYER VI3 ;
  RECT 1135.040 6.340 1135.240 6.540 ;
  LAYER VI3 ;
  RECT 1135.040 5.940 1135.240 6.140 ;
  LAYER VI3 ;
  RECT 1134.640 6.340 1134.840 6.540 ;
  LAYER VI3 ;
  RECT 1134.640 5.940 1134.840 6.140 ;
  LAYER VI3 ;
  RECT 1134.240 6.340 1134.440 6.540 ;
  LAYER VI3 ;
  RECT 1134.240 5.940 1134.440 6.140 ;
  LAYER VI3 ;
  RECT 1133.840 6.340 1134.040 6.540 ;
  LAYER VI3 ;
  RECT 1133.840 5.940 1134.040 6.140 ;
  LAYER VI3 ;
  RECT 1133.440 6.340 1133.640 6.540 ;
  LAYER VI3 ;
  RECT 1133.440 5.940 1133.640 6.140 ;
  LAYER VI3 ;
  RECT 1133.040 6.340 1133.240 6.540 ;
  LAYER VI3 ;
  RECT 1133.040 5.940 1133.240 6.140 ;
  LAYER VI3 ;
  RECT 1154.120 5.880 1162.120 6.740 ;
  LAYER VI3 ;
  RECT 1161.720 6.340 1161.920 6.540 ;
  LAYER VI3 ;
  RECT 1161.720 5.940 1161.920 6.140 ;
  LAYER VI3 ;
  RECT 1161.320 6.340 1161.520 6.540 ;
  LAYER VI3 ;
  RECT 1161.320 5.940 1161.520 6.140 ;
  LAYER VI3 ;
  RECT 1160.920 6.340 1161.120 6.540 ;
  LAYER VI3 ;
  RECT 1160.920 5.940 1161.120 6.140 ;
  LAYER VI3 ;
  RECT 1160.520 6.340 1160.720 6.540 ;
  LAYER VI3 ;
  RECT 1160.520 5.940 1160.720 6.140 ;
  LAYER VI3 ;
  RECT 1160.120 6.340 1160.320 6.540 ;
  LAYER VI3 ;
  RECT 1160.120 5.940 1160.320 6.140 ;
  LAYER VI3 ;
  RECT 1159.720 6.340 1159.920 6.540 ;
  LAYER VI3 ;
  RECT 1159.720 5.940 1159.920 6.140 ;
  LAYER VI3 ;
  RECT 1159.320 6.340 1159.520 6.540 ;
  LAYER VI3 ;
  RECT 1159.320 5.940 1159.520 6.140 ;
  LAYER VI3 ;
  RECT 1158.920 6.340 1159.120 6.540 ;
  LAYER VI3 ;
  RECT 1158.920 5.940 1159.120 6.140 ;
  LAYER VI3 ;
  RECT 1158.520 6.340 1158.720 6.540 ;
  LAYER VI3 ;
  RECT 1158.520 5.940 1158.720 6.140 ;
  LAYER VI3 ;
  RECT 1158.120 6.340 1158.320 6.540 ;
  LAYER VI3 ;
  RECT 1158.120 5.940 1158.320 6.140 ;
  LAYER VI3 ;
  RECT 1157.720 6.340 1157.920 6.540 ;
  LAYER VI3 ;
  RECT 1157.720 5.940 1157.920 6.140 ;
  LAYER VI3 ;
  RECT 1157.320 6.340 1157.520 6.540 ;
  LAYER VI3 ;
  RECT 1157.320 5.940 1157.520 6.140 ;
  LAYER VI3 ;
  RECT 1156.920 6.340 1157.120 6.540 ;
  LAYER VI3 ;
  RECT 1156.920 5.940 1157.120 6.140 ;
  LAYER VI3 ;
  RECT 1156.520 6.340 1156.720 6.540 ;
  LAYER VI3 ;
  RECT 1156.520 5.940 1156.720 6.140 ;
  LAYER VI3 ;
  RECT 1156.120 6.340 1156.320 6.540 ;
  LAYER VI3 ;
  RECT 1156.120 5.940 1156.320 6.140 ;
  LAYER VI3 ;
  RECT 1155.720 6.340 1155.920 6.540 ;
  LAYER VI3 ;
  RECT 1155.720 5.940 1155.920 6.140 ;
  LAYER VI3 ;
  RECT 1155.320 6.340 1155.520 6.540 ;
  LAYER VI3 ;
  RECT 1155.320 5.940 1155.520 6.140 ;
  LAYER VI3 ;
  RECT 1154.920 6.340 1155.120 6.540 ;
  LAYER VI3 ;
  RECT 1154.920 5.940 1155.120 6.140 ;
  LAYER VI3 ;
  RECT 1154.520 6.340 1154.720 6.540 ;
  LAYER VI3 ;
  RECT 1154.520 5.940 1154.720 6.140 ;
  LAYER VI3 ;
  RECT 1154.120 6.340 1154.320 6.540 ;
  LAYER VI3 ;
  RECT 1154.120 5.940 1154.320 6.140 ;
  LAYER VI3 ;
  RECT 1173.960 5.880 1181.960 6.740 ;
  LAYER VI3 ;
  RECT 1181.560 6.340 1181.760 6.540 ;
  LAYER VI3 ;
  RECT 1181.560 5.940 1181.760 6.140 ;
  LAYER VI3 ;
  RECT 1181.160 6.340 1181.360 6.540 ;
  LAYER VI3 ;
  RECT 1181.160 5.940 1181.360 6.140 ;
  LAYER VI3 ;
  RECT 1180.760 6.340 1180.960 6.540 ;
  LAYER VI3 ;
  RECT 1180.760 5.940 1180.960 6.140 ;
  LAYER VI3 ;
  RECT 1180.360 6.340 1180.560 6.540 ;
  LAYER VI3 ;
  RECT 1180.360 5.940 1180.560 6.140 ;
  LAYER VI3 ;
  RECT 1179.960 6.340 1180.160 6.540 ;
  LAYER VI3 ;
  RECT 1179.960 5.940 1180.160 6.140 ;
  LAYER VI3 ;
  RECT 1179.560 6.340 1179.760 6.540 ;
  LAYER VI3 ;
  RECT 1179.560 5.940 1179.760 6.140 ;
  LAYER VI3 ;
  RECT 1179.160 6.340 1179.360 6.540 ;
  LAYER VI3 ;
  RECT 1179.160 5.940 1179.360 6.140 ;
  LAYER VI3 ;
  RECT 1178.760 6.340 1178.960 6.540 ;
  LAYER VI3 ;
  RECT 1178.760 5.940 1178.960 6.140 ;
  LAYER VI3 ;
  RECT 1178.360 6.340 1178.560 6.540 ;
  LAYER VI3 ;
  RECT 1178.360 5.940 1178.560 6.140 ;
  LAYER VI3 ;
  RECT 1177.960 6.340 1178.160 6.540 ;
  LAYER VI3 ;
  RECT 1177.960 5.940 1178.160 6.140 ;
  LAYER VI3 ;
  RECT 1177.560 6.340 1177.760 6.540 ;
  LAYER VI3 ;
  RECT 1177.560 5.940 1177.760 6.140 ;
  LAYER VI3 ;
  RECT 1177.160 6.340 1177.360 6.540 ;
  LAYER VI3 ;
  RECT 1177.160 5.940 1177.360 6.140 ;
  LAYER VI3 ;
  RECT 1176.760 6.340 1176.960 6.540 ;
  LAYER VI3 ;
  RECT 1176.760 5.940 1176.960 6.140 ;
  LAYER VI3 ;
  RECT 1176.360 6.340 1176.560 6.540 ;
  LAYER VI3 ;
  RECT 1176.360 5.940 1176.560 6.140 ;
  LAYER VI3 ;
  RECT 1175.960 6.340 1176.160 6.540 ;
  LAYER VI3 ;
  RECT 1175.960 5.940 1176.160 6.140 ;
  LAYER VI3 ;
  RECT 1175.560 6.340 1175.760 6.540 ;
  LAYER VI3 ;
  RECT 1175.560 5.940 1175.760 6.140 ;
  LAYER VI3 ;
  RECT 1175.160 6.340 1175.360 6.540 ;
  LAYER VI3 ;
  RECT 1175.160 5.940 1175.360 6.140 ;
  LAYER VI3 ;
  RECT 1174.760 6.340 1174.960 6.540 ;
  LAYER VI3 ;
  RECT 1174.760 5.940 1174.960 6.140 ;
  LAYER VI3 ;
  RECT 1174.360 6.340 1174.560 6.540 ;
  LAYER VI3 ;
  RECT 1174.360 5.940 1174.560 6.140 ;
  LAYER VI3 ;
  RECT 1173.960 6.340 1174.160 6.540 ;
  LAYER VI3 ;
  RECT 1173.960 5.940 1174.160 6.140 ;
  LAYER VI3 ;
  RECT 1195.040 5.880 1203.040 6.740 ;
  LAYER VI3 ;
  RECT 1202.640 6.340 1202.840 6.540 ;
  LAYER VI3 ;
  RECT 1202.640 5.940 1202.840 6.140 ;
  LAYER VI3 ;
  RECT 1202.240 6.340 1202.440 6.540 ;
  LAYER VI3 ;
  RECT 1202.240 5.940 1202.440 6.140 ;
  LAYER VI3 ;
  RECT 1201.840 6.340 1202.040 6.540 ;
  LAYER VI3 ;
  RECT 1201.840 5.940 1202.040 6.140 ;
  LAYER VI3 ;
  RECT 1201.440 6.340 1201.640 6.540 ;
  LAYER VI3 ;
  RECT 1201.440 5.940 1201.640 6.140 ;
  LAYER VI3 ;
  RECT 1201.040 6.340 1201.240 6.540 ;
  LAYER VI3 ;
  RECT 1201.040 5.940 1201.240 6.140 ;
  LAYER VI3 ;
  RECT 1200.640 6.340 1200.840 6.540 ;
  LAYER VI3 ;
  RECT 1200.640 5.940 1200.840 6.140 ;
  LAYER VI3 ;
  RECT 1200.240 6.340 1200.440 6.540 ;
  LAYER VI3 ;
  RECT 1200.240 5.940 1200.440 6.140 ;
  LAYER VI3 ;
  RECT 1199.840 6.340 1200.040 6.540 ;
  LAYER VI3 ;
  RECT 1199.840 5.940 1200.040 6.140 ;
  LAYER VI3 ;
  RECT 1199.440 6.340 1199.640 6.540 ;
  LAYER VI3 ;
  RECT 1199.440 5.940 1199.640 6.140 ;
  LAYER VI3 ;
  RECT 1199.040 6.340 1199.240 6.540 ;
  LAYER VI3 ;
  RECT 1199.040 5.940 1199.240 6.140 ;
  LAYER VI3 ;
  RECT 1198.640 6.340 1198.840 6.540 ;
  LAYER VI3 ;
  RECT 1198.640 5.940 1198.840 6.140 ;
  LAYER VI3 ;
  RECT 1198.240 6.340 1198.440 6.540 ;
  LAYER VI3 ;
  RECT 1198.240 5.940 1198.440 6.140 ;
  LAYER VI3 ;
  RECT 1197.840 6.340 1198.040 6.540 ;
  LAYER VI3 ;
  RECT 1197.840 5.940 1198.040 6.140 ;
  LAYER VI3 ;
  RECT 1197.440 6.340 1197.640 6.540 ;
  LAYER VI3 ;
  RECT 1197.440 5.940 1197.640 6.140 ;
  LAYER VI3 ;
  RECT 1197.040 6.340 1197.240 6.540 ;
  LAYER VI3 ;
  RECT 1197.040 5.940 1197.240 6.140 ;
  LAYER VI3 ;
  RECT 1196.640 6.340 1196.840 6.540 ;
  LAYER VI3 ;
  RECT 1196.640 5.940 1196.840 6.140 ;
  LAYER VI3 ;
  RECT 1196.240 6.340 1196.440 6.540 ;
  LAYER VI3 ;
  RECT 1196.240 5.940 1196.440 6.140 ;
  LAYER VI3 ;
  RECT 1195.840 6.340 1196.040 6.540 ;
  LAYER VI3 ;
  RECT 1195.840 5.940 1196.040 6.140 ;
  LAYER VI3 ;
  RECT 1195.440 6.340 1195.640 6.540 ;
  LAYER VI3 ;
  RECT 1195.440 5.940 1195.640 6.140 ;
  LAYER VI3 ;
  RECT 1195.040 6.340 1195.240 6.540 ;
  LAYER VI3 ;
  RECT 1195.040 5.940 1195.240 6.140 ;
  LAYER VI3 ;
  RECT 1214.880 5.880 1222.880 6.740 ;
  LAYER VI3 ;
  RECT 1222.480 6.340 1222.680 6.540 ;
  LAYER VI3 ;
  RECT 1222.480 5.940 1222.680 6.140 ;
  LAYER VI3 ;
  RECT 1222.080 6.340 1222.280 6.540 ;
  LAYER VI3 ;
  RECT 1222.080 5.940 1222.280 6.140 ;
  LAYER VI3 ;
  RECT 1221.680 6.340 1221.880 6.540 ;
  LAYER VI3 ;
  RECT 1221.680 5.940 1221.880 6.140 ;
  LAYER VI3 ;
  RECT 1221.280 6.340 1221.480 6.540 ;
  LAYER VI3 ;
  RECT 1221.280 5.940 1221.480 6.140 ;
  LAYER VI3 ;
  RECT 1220.880 6.340 1221.080 6.540 ;
  LAYER VI3 ;
  RECT 1220.880 5.940 1221.080 6.140 ;
  LAYER VI3 ;
  RECT 1220.480 6.340 1220.680 6.540 ;
  LAYER VI3 ;
  RECT 1220.480 5.940 1220.680 6.140 ;
  LAYER VI3 ;
  RECT 1220.080 6.340 1220.280 6.540 ;
  LAYER VI3 ;
  RECT 1220.080 5.940 1220.280 6.140 ;
  LAYER VI3 ;
  RECT 1219.680 6.340 1219.880 6.540 ;
  LAYER VI3 ;
  RECT 1219.680 5.940 1219.880 6.140 ;
  LAYER VI3 ;
  RECT 1219.280 6.340 1219.480 6.540 ;
  LAYER VI3 ;
  RECT 1219.280 5.940 1219.480 6.140 ;
  LAYER VI3 ;
  RECT 1218.880 6.340 1219.080 6.540 ;
  LAYER VI3 ;
  RECT 1218.880 5.940 1219.080 6.140 ;
  LAYER VI3 ;
  RECT 1218.480 6.340 1218.680 6.540 ;
  LAYER VI3 ;
  RECT 1218.480 5.940 1218.680 6.140 ;
  LAYER VI3 ;
  RECT 1218.080 6.340 1218.280 6.540 ;
  LAYER VI3 ;
  RECT 1218.080 5.940 1218.280 6.140 ;
  LAYER VI3 ;
  RECT 1217.680 6.340 1217.880 6.540 ;
  LAYER VI3 ;
  RECT 1217.680 5.940 1217.880 6.140 ;
  LAYER VI3 ;
  RECT 1217.280 6.340 1217.480 6.540 ;
  LAYER VI3 ;
  RECT 1217.280 5.940 1217.480 6.140 ;
  LAYER VI3 ;
  RECT 1216.880 6.340 1217.080 6.540 ;
  LAYER VI3 ;
  RECT 1216.880 5.940 1217.080 6.140 ;
  LAYER VI3 ;
  RECT 1216.480 6.340 1216.680 6.540 ;
  LAYER VI3 ;
  RECT 1216.480 5.940 1216.680 6.140 ;
  LAYER VI3 ;
  RECT 1216.080 6.340 1216.280 6.540 ;
  LAYER VI3 ;
  RECT 1216.080 5.940 1216.280 6.140 ;
  LAYER VI3 ;
  RECT 1215.680 6.340 1215.880 6.540 ;
  LAYER VI3 ;
  RECT 1215.680 5.940 1215.880 6.140 ;
  LAYER VI3 ;
  RECT 1215.280 6.340 1215.480 6.540 ;
  LAYER VI3 ;
  RECT 1215.280 5.940 1215.480 6.140 ;
  LAYER VI3 ;
  RECT 1214.880 6.340 1215.080 6.540 ;
  LAYER VI3 ;
  RECT 1214.880 5.940 1215.080 6.140 ;
  LAYER VI3 ;
  RECT 1235.960 5.880 1243.960 6.740 ;
  LAYER VI3 ;
  RECT 1243.560 6.340 1243.760 6.540 ;
  LAYER VI3 ;
  RECT 1243.560 5.940 1243.760 6.140 ;
  LAYER VI3 ;
  RECT 1243.160 6.340 1243.360 6.540 ;
  LAYER VI3 ;
  RECT 1243.160 5.940 1243.360 6.140 ;
  LAYER VI3 ;
  RECT 1242.760 6.340 1242.960 6.540 ;
  LAYER VI3 ;
  RECT 1242.760 5.940 1242.960 6.140 ;
  LAYER VI3 ;
  RECT 1242.360 6.340 1242.560 6.540 ;
  LAYER VI3 ;
  RECT 1242.360 5.940 1242.560 6.140 ;
  LAYER VI3 ;
  RECT 1241.960 6.340 1242.160 6.540 ;
  LAYER VI3 ;
  RECT 1241.960 5.940 1242.160 6.140 ;
  LAYER VI3 ;
  RECT 1241.560 6.340 1241.760 6.540 ;
  LAYER VI3 ;
  RECT 1241.560 5.940 1241.760 6.140 ;
  LAYER VI3 ;
  RECT 1241.160 6.340 1241.360 6.540 ;
  LAYER VI3 ;
  RECT 1241.160 5.940 1241.360 6.140 ;
  LAYER VI3 ;
  RECT 1240.760 6.340 1240.960 6.540 ;
  LAYER VI3 ;
  RECT 1240.760 5.940 1240.960 6.140 ;
  LAYER VI3 ;
  RECT 1240.360 6.340 1240.560 6.540 ;
  LAYER VI3 ;
  RECT 1240.360 5.940 1240.560 6.140 ;
  LAYER VI3 ;
  RECT 1239.960 6.340 1240.160 6.540 ;
  LAYER VI3 ;
  RECT 1239.960 5.940 1240.160 6.140 ;
  LAYER VI3 ;
  RECT 1239.560 6.340 1239.760 6.540 ;
  LAYER VI3 ;
  RECT 1239.560 5.940 1239.760 6.140 ;
  LAYER VI3 ;
  RECT 1239.160 6.340 1239.360 6.540 ;
  LAYER VI3 ;
  RECT 1239.160 5.940 1239.360 6.140 ;
  LAYER VI3 ;
  RECT 1238.760 6.340 1238.960 6.540 ;
  LAYER VI3 ;
  RECT 1238.760 5.940 1238.960 6.140 ;
  LAYER VI3 ;
  RECT 1238.360 6.340 1238.560 6.540 ;
  LAYER VI3 ;
  RECT 1238.360 5.940 1238.560 6.140 ;
  LAYER VI3 ;
  RECT 1237.960 6.340 1238.160 6.540 ;
  LAYER VI3 ;
  RECT 1237.960 5.940 1238.160 6.140 ;
  LAYER VI3 ;
  RECT 1237.560 6.340 1237.760 6.540 ;
  LAYER VI3 ;
  RECT 1237.560 5.940 1237.760 6.140 ;
  LAYER VI3 ;
  RECT 1237.160 6.340 1237.360 6.540 ;
  LAYER VI3 ;
  RECT 1237.160 5.940 1237.360 6.140 ;
  LAYER VI3 ;
  RECT 1236.760 6.340 1236.960 6.540 ;
  LAYER VI3 ;
  RECT 1236.760 5.940 1236.960 6.140 ;
  LAYER VI3 ;
  RECT 1236.360 6.340 1236.560 6.540 ;
  LAYER VI3 ;
  RECT 1236.360 5.940 1236.560 6.140 ;
  LAYER VI3 ;
  RECT 1235.960 6.340 1236.160 6.540 ;
  LAYER VI3 ;
  RECT 1235.960 5.940 1236.160 6.140 ;
  LAYER VI3 ;
  RECT 1255.800 5.880 1263.800 6.740 ;
  LAYER VI3 ;
  RECT 1263.400 6.340 1263.600 6.540 ;
  LAYER VI3 ;
  RECT 1263.400 5.940 1263.600 6.140 ;
  LAYER VI3 ;
  RECT 1263.000 6.340 1263.200 6.540 ;
  LAYER VI3 ;
  RECT 1263.000 5.940 1263.200 6.140 ;
  LAYER VI3 ;
  RECT 1262.600 6.340 1262.800 6.540 ;
  LAYER VI3 ;
  RECT 1262.600 5.940 1262.800 6.140 ;
  LAYER VI3 ;
  RECT 1262.200 6.340 1262.400 6.540 ;
  LAYER VI3 ;
  RECT 1262.200 5.940 1262.400 6.140 ;
  LAYER VI3 ;
  RECT 1261.800 6.340 1262.000 6.540 ;
  LAYER VI3 ;
  RECT 1261.800 5.940 1262.000 6.140 ;
  LAYER VI3 ;
  RECT 1261.400 6.340 1261.600 6.540 ;
  LAYER VI3 ;
  RECT 1261.400 5.940 1261.600 6.140 ;
  LAYER VI3 ;
  RECT 1261.000 6.340 1261.200 6.540 ;
  LAYER VI3 ;
  RECT 1261.000 5.940 1261.200 6.140 ;
  LAYER VI3 ;
  RECT 1260.600 6.340 1260.800 6.540 ;
  LAYER VI3 ;
  RECT 1260.600 5.940 1260.800 6.140 ;
  LAYER VI3 ;
  RECT 1260.200 6.340 1260.400 6.540 ;
  LAYER VI3 ;
  RECT 1260.200 5.940 1260.400 6.140 ;
  LAYER VI3 ;
  RECT 1259.800 6.340 1260.000 6.540 ;
  LAYER VI3 ;
  RECT 1259.800 5.940 1260.000 6.140 ;
  LAYER VI3 ;
  RECT 1259.400 6.340 1259.600 6.540 ;
  LAYER VI3 ;
  RECT 1259.400 5.940 1259.600 6.140 ;
  LAYER VI3 ;
  RECT 1259.000 6.340 1259.200 6.540 ;
  LAYER VI3 ;
  RECT 1259.000 5.940 1259.200 6.140 ;
  LAYER VI3 ;
  RECT 1258.600 6.340 1258.800 6.540 ;
  LAYER VI3 ;
  RECT 1258.600 5.940 1258.800 6.140 ;
  LAYER VI3 ;
  RECT 1258.200 6.340 1258.400 6.540 ;
  LAYER VI3 ;
  RECT 1258.200 5.940 1258.400 6.140 ;
  LAYER VI3 ;
  RECT 1257.800 6.340 1258.000 6.540 ;
  LAYER VI3 ;
  RECT 1257.800 5.940 1258.000 6.140 ;
  LAYER VI3 ;
  RECT 1257.400 6.340 1257.600 6.540 ;
  LAYER VI3 ;
  RECT 1257.400 5.940 1257.600 6.140 ;
  LAYER VI3 ;
  RECT 1257.000 6.340 1257.200 6.540 ;
  LAYER VI3 ;
  RECT 1257.000 5.940 1257.200 6.140 ;
  LAYER VI3 ;
  RECT 1256.600 6.340 1256.800 6.540 ;
  LAYER VI3 ;
  RECT 1256.600 5.940 1256.800 6.140 ;
  LAYER VI3 ;
  RECT 1256.200 6.340 1256.400 6.540 ;
  LAYER VI3 ;
  RECT 1256.200 5.940 1256.400 6.140 ;
  LAYER VI3 ;
  RECT 1255.800 6.340 1256.000 6.540 ;
  LAYER VI3 ;
  RECT 1255.800 5.940 1256.000 6.140 ;
  LAYER VI3 ;
  RECT 1276.880 5.880 1284.880 6.740 ;
  LAYER VI3 ;
  RECT 1284.480 6.340 1284.680 6.540 ;
  LAYER VI3 ;
  RECT 1284.480 5.940 1284.680 6.140 ;
  LAYER VI3 ;
  RECT 1284.080 6.340 1284.280 6.540 ;
  LAYER VI3 ;
  RECT 1284.080 5.940 1284.280 6.140 ;
  LAYER VI3 ;
  RECT 1283.680 6.340 1283.880 6.540 ;
  LAYER VI3 ;
  RECT 1283.680 5.940 1283.880 6.140 ;
  LAYER VI3 ;
  RECT 1283.280 6.340 1283.480 6.540 ;
  LAYER VI3 ;
  RECT 1283.280 5.940 1283.480 6.140 ;
  LAYER VI3 ;
  RECT 1282.880 6.340 1283.080 6.540 ;
  LAYER VI3 ;
  RECT 1282.880 5.940 1283.080 6.140 ;
  LAYER VI3 ;
  RECT 1282.480 6.340 1282.680 6.540 ;
  LAYER VI3 ;
  RECT 1282.480 5.940 1282.680 6.140 ;
  LAYER VI3 ;
  RECT 1282.080 6.340 1282.280 6.540 ;
  LAYER VI3 ;
  RECT 1282.080 5.940 1282.280 6.140 ;
  LAYER VI3 ;
  RECT 1281.680 6.340 1281.880 6.540 ;
  LAYER VI3 ;
  RECT 1281.680 5.940 1281.880 6.140 ;
  LAYER VI3 ;
  RECT 1281.280 6.340 1281.480 6.540 ;
  LAYER VI3 ;
  RECT 1281.280 5.940 1281.480 6.140 ;
  LAYER VI3 ;
  RECT 1280.880 6.340 1281.080 6.540 ;
  LAYER VI3 ;
  RECT 1280.880 5.940 1281.080 6.140 ;
  LAYER VI3 ;
  RECT 1280.480 6.340 1280.680 6.540 ;
  LAYER VI3 ;
  RECT 1280.480 5.940 1280.680 6.140 ;
  LAYER VI3 ;
  RECT 1280.080 6.340 1280.280 6.540 ;
  LAYER VI3 ;
  RECT 1280.080 5.940 1280.280 6.140 ;
  LAYER VI3 ;
  RECT 1279.680 6.340 1279.880 6.540 ;
  LAYER VI3 ;
  RECT 1279.680 5.940 1279.880 6.140 ;
  LAYER VI3 ;
  RECT 1279.280 6.340 1279.480 6.540 ;
  LAYER VI3 ;
  RECT 1279.280 5.940 1279.480 6.140 ;
  LAYER VI3 ;
  RECT 1278.880 6.340 1279.080 6.540 ;
  LAYER VI3 ;
  RECT 1278.880 5.940 1279.080 6.140 ;
  LAYER VI3 ;
  RECT 1278.480 6.340 1278.680 6.540 ;
  LAYER VI3 ;
  RECT 1278.480 5.940 1278.680 6.140 ;
  LAYER VI3 ;
  RECT 1278.080 6.340 1278.280 6.540 ;
  LAYER VI3 ;
  RECT 1278.080 5.940 1278.280 6.140 ;
  LAYER VI3 ;
  RECT 1277.680 6.340 1277.880 6.540 ;
  LAYER VI3 ;
  RECT 1277.680 5.940 1277.880 6.140 ;
  LAYER VI3 ;
  RECT 1277.280 6.340 1277.480 6.540 ;
  LAYER VI3 ;
  RECT 1277.280 5.940 1277.480 6.140 ;
  LAYER VI3 ;
  RECT 1276.880 6.340 1277.080 6.540 ;
  LAYER VI3 ;
  RECT 1276.880 5.940 1277.080 6.140 ;
  LAYER VI3 ;
  RECT 1296.720 5.880 1304.720 6.740 ;
  LAYER VI3 ;
  RECT 1304.320 6.340 1304.520 6.540 ;
  LAYER VI3 ;
  RECT 1304.320 5.940 1304.520 6.140 ;
  LAYER VI3 ;
  RECT 1303.920 6.340 1304.120 6.540 ;
  LAYER VI3 ;
  RECT 1303.920 5.940 1304.120 6.140 ;
  LAYER VI3 ;
  RECT 1303.520 6.340 1303.720 6.540 ;
  LAYER VI3 ;
  RECT 1303.520 5.940 1303.720 6.140 ;
  LAYER VI3 ;
  RECT 1303.120 6.340 1303.320 6.540 ;
  LAYER VI3 ;
  RECT 1303.120 5.940 1303.320 6.140 ;
  LAYER VI3 ;
  RECT 1302.720 6.340 1302.920 6.540 ;
  LAYER VI3 ;
  RECT 1302.720 5.940 1302.920 6.140 ;
  LAYER VI3 ;
  RECT 1302.320 6.340 1302.520 6.540 ;
  LAYER VI3 ;
  RECT 1302.320 5.940 1302.520 6.140 ;
  LAYER VI3 ;
  RECT 1301.920 6.340 1302.120 6.540 ;
  LAYER VI3 ;
  RECT 1301.920 5.940 1302.120 6.140 ;
  LAYER VI3 ;
  RECT 1301.520 6.340 1301.720 6.540 ;
  LAYER VI3 ;
  RECT 1301.520 5.940 1301.720 6.140 ;
  LAYER VI3 ;
  RECT 1301.120 6.340 1301.320 6.540 ;
  LAYER VI3 ;
  RECT 1301.120 5.940 1301.320 6.140 ;
  LAYER VI3 ;
  RECT 1300.720 6.340 1300.920 6.540 ;
  LAYER VI3 ;
  RECT 1300.720 5.940 1300.920 6.140 ;
  LAYER VI3 ;
  RECT 1300.320 6.340 1300.520 6.540 ;
  LAYER VI3 ;
  RECT 1300.320 5.940 1300.520 6.140 ;
  LAYER VI3 ;
  RECT 1299.920 6.340 1300.120 6.540 ;
  LAYER VI3 ;
  RECT 1299.920 5.940 1300.120 6.140 ;
  LAYER VI3 ;
  RECT 1299.520 6.340 1299.720 6.540 ;
  LAYER VI3 ;
  RECT 1299.520 5.940 1299.720 6.140 ;
  LAYER VI3 ;
  RECT 1299.120 6.340 1299.320 6.540 ;
  LAYER VI3 ;
  RECT 1299.120 5.940 1299.320 6.140 ;
  LAYER VI3 ;
  RECT 1298.720 6.340 1298.920 6.540 ;
  LAYER VI3 ;
  RECT 1298.720 5.940 1298.920 6.140 ;
  LAYER VI3 ;
  RECT 1298.320 6.340 1298.520 6.540 ;
  LAYER VI3 ;
  RECT 1298.320 5.940 1298.520 6.140 ;
  LAYER VI3 ;
  RECT 1297.920 6.340 1298.120 6.540 ;
  LAYER VI3 ;
  RECT 1297.920 5.940 1298.120 6.140 ;
  LAYER VI3 ;
  RECT 1297.520 6.340 1297.720 6.540 ;
  LAYER VI3 ;
  RECT 1297.520 5.940 1297.720 6.140 ;
  LAYER VI3 ;
  RECT 1297.120 6.340 1297.320 6.540 ;
  LAYER VI3 ;
  RECT 1297.120 5.940 1297.320 6.140 ;
  LAYER VI3 ;
  RECT 1296.720 6.340 1296.920 6.540 ;
  LAYER VI3 ;
  RECT 1296.720 5.940 1296.920 6.140 ;
  LAYER VI3 ;
  RECT 2687.800 559.940 2688.660 560.320 ;
  LAYER VI3 ;
  RECT 2688.200 560.000 2688.400 560.200 ;
  LAYER VI3 ;
  RECT 2687.800 560.000 2688.000 560.200 ;
  LAYER VI2 ;
  RECT 2687.800 559.940 2688.660 560.320 ;
  LAYER VI2 ;
  RECT 2688.200 560.000 2688.400 560.200 ;
  LAYER VI2 ;
  RECT 2687.800 560.000 2688.000 560.200 ;
  LAYER VI3 ;
  RECT 2687.800 552.020 2688.660 552.300 ;
  LAYER VI3 ;
  RECT 2688.260 552.020 2688.460 552.220 ;
  LAYER VI3 ;
  RECT 2687.860 552.020 2688.060 552.220 ;
  LAYER VI2 ;
  RECT 2687.800 552.020 2688.660 552.300 ;
  LAYER VI2 ;
  RECT 2688.260 552.020 2688.460 552.220 ;
  LAYER VI2 ;
  RECT 2687.860 552.020 2688.060 552.220 ;
  LAYER VI3 ;
  RECT 2687.800 548.340 2688.660 548.620 ;
  LAYER VI3 ;
  RECT 2688.260 548.340 2688.460 548.540 ;
  LAYER VI3 ;
  RECT 2687.860 548.340 2688.060 548.540 ;
  LAYER VI2 ;
  RECT 2687.800 548.340 2688.660 548.620 ;
  LAYER VI2 ;
  RECT 2688.260 548.340 2688.460 548.540 ;
  LAYER VI2 ;
  RECT 2687.860 548.340 2688.060 548.540 ;
  LAYER VI3 ;
  RECT 2687.800 544.660 2688.660 544.940 ;
  LAYER VI3 ;
  RECT 2688.260 544.660 2688.460 544.860 ;
  LAYER VI3 ;
  RECT 2687.860 544.660 2688.060 544.860 ;
  LAYER VI2 ;
  RECT 2687.800 544.660 2688.660 544.940 ;
  LAYER VI2 ;
  RECT 2688.260 544.660 2688.460 544.860 ;
  LAYER VI2 ;
  RECT 2687.860 544.660 2688.060 544.860 ;
  LAYER VI3 ;
  RECT 2687.800 540.980 2688.660 541.260 ;
  LAYER VI3 ;
  RECT 2688.260 540.980 2688.460 541.180 ;
  LAYER VI3 ;
  RECT 2687.860 540.980 2688.060 541.180 ;
  LAYER VI2 ;
  RECT 2687.800 540.980 2688.660 541.260 ;
  LAYER VI2 ;
  RECT 2688.260 540.980 2688.460 541.180 ;
  LAYER VI2 ;
  RECT 2687.860 540.980 2688.060 541.180 ;
  LAYER VI3 ;
  RECT 2687.800 537.300 2688.660 537.580 ;
  LAYER VI3 ;
  RECT 2688.260 537.300 2688.460 537.500 ;
  LAYER VI3 ;
  RECT 2687.860 537.300 2688.060 537.500 ;
  LAYER VI2 ;
  RECT 2687.800 537.300 2688.660 537.580 ;
  LAYER VI2 ;
  RECT 2688.260 537.300 2688.460 537.500 ;
  LAYER VI2 ;
  RECT 2687.860 537.300 2688.060 537.500 ;
  LAYER VI3 ;
  RECT 2687.800 533.620 2688.660 533.900 ;
  LAYER VI3 ;
  RECT 2688.260 533.620 2688.460 533.820 ;
  LAYER VI3 ;
  RECT 2687.860 533.620 2688.060 533.820 ;
  LAYER VI2 ;
  RECT 2687.800 533.620 2688.660 533.900 ;
  LAYER VI2 ;
  RECT 2688.260 533.620 2688.460 533.820 ;
  LAYER VI2 ;
  RECT 2687.860 533.620 2688.060 533.820 ;
  LAYER VI3 ;
  RECT 2687.800 529.940 2688.660 530.220 ;
  LAYER VI3 ;
  RECT 2688.260 529.940 2688.460 530.140 ;
  LAYER VI3 ;
  RECT 2687.860 529.940 2688.060 530.140 ;
  LAYER VI2 ;
  RECT 2687.800 529.940 2688.660 530.220 ;
  LAYER VI2 ;
  RECT 2688.260 529.940 2688.460 530.140 ;
  LAYER VI2 ;
  RECT 2687.860 529.940 2688.060 530.140 ;
  LAYER VI3 ;
  RECT 2687.800 526.260 2688.660 526.540 ;
  LAYER VI3 ;
  RECT 2688.260 526.260 2688.460 526.460 ;
  LAYER VI3 ;
  RECT 2687.860 526.260 2688.060 526.460 ;
  LAYER VI2 ;
  RECT 2687.800 526.260 2688.660 526.540 ;
  LAYER VI2 ;
  RECT 2688.260 526.260 2688.460 526.460 ;
  LAYER VI2 ;
  RECT 2687.860 526.260 2688.060 526.460 ;
  LAYER VI3 ;
  RECT 2687.800 522.580 2688.660 522.860 ;
  LAYER VI3 ;
  RECT 2688.260 522.580 2688.460 522.780 ;
  LAYER VI3 ;
  RECT 2687.860 522.580 2688.060 522.780 ;
  LAYER VI2 ;
  RECT 2687.800 522.580 2688.660 522.860 ;
  LAYER VI2 ;
  RECT 2688.260 522.580 2688.460 522.780 ;
  LAYER VI2 ;
  RECT 2687.860 522.580 2688.060 522.780 ;
  LAYER VI3 ;
  RECT 2687.800 518.900 2688.660 519.180 ;
  LAYER VI3 ;
  RECT 2688.260 518.900 2688.460 519.100 ;
  LAYER VI3 ;
  RECT 2687.860 518.900 2688.060 519.100 ;
  LAYER VI2 ;
  RECT 2687.800 518.900 2688.660 519.180 ;
  LAYER VI2 ;
  RECT 2688.260 518.900 2688.460 519.100 ;
  LAYER VI2 ;
  RECT 2687.860 518.900 2688.060 519.100 ;
  LAYER VI3 ;
  RECT 2687.800 515.220 2688.660 515.500 ;
  LAYER VI3 ;
  RECT 2688.260 515.220 2688.460 515.420 ;
  LAYER VI3 ;
  RECT 2687.860 515.220 2688.060 515.420 ;
  LAYER VI2 ;
  RECT 2687.800 515.220 2688.660 515.500 ;
  LAYER VI2 ;
  RECT 2688.260 515.220 2688.460 515.420 ;
  LAYER VI2 ;
  RECT 2687.860 515.220 2688.060 515.420 ;
  LAYER VI3 ;
  RECT 2687.800 511.540 2688.660 511.820 ;
  LAYER VI3 ;
  RECT 2688.260 511.540 2688.460 511.740 ;
  LAYER VI3 ;
  RECT 2687.860 511.540 2688.060 511.740 ;
  LAYER VI2 ;
  RECT 2687.800 511.540 2688.660 511.820 ;
  LAYER VI2 ;
  RECT 2688.260 511.540 2688.460 511.740 ;
  LAYER VI2 ;
  RECT 2687.860 511.540 2688.060 511.740 ;
  LAYER VI3 ;
  RECT 2687.800 507.860 2688.660 508.140 ;
  LAYER VI3 ;
  RECT 2688.260 507.860 2688.460 508.060 ;
  LAYER VI3 ;
  RECT 2687.860 507.860 2688.060 508.060 ;
  LAYER VI2 ;
  RECT 2687.800 507.860 2688.660 508.140 ;
  LAYER VI2 ;
  RECT 2688.260 507.860 2688.460 508.060 ;
  LAYER VI2 ;
  RECT 2687.860 507.860 2688.060 508.060 ;
  LAYER VI3 ;
  RECT 2687.800 504.180 2688.660 504.460 ;
  LAYER VI3 ;
  RECT 2688.260 504.180 2688.460 504.380 ;
  LAYER VI3 ;
  RECT 2687.860 504.180 2688.060 504.380 ;
  LAYER VI2 ;
  RECT 2687.800 504.180 2688.660 504.460 ;
  LAYER VI2 ;
  RECT 2688.260 504.180 2688.460 504.380 ;
  LAYER VI2 ;
  RECT 2687.860 504.180 2688.060 504.380 ;
  LAYER VI3 ;
  RECT 2687.800 500.500 2688.660 500.780 ;
  LAYER VI3 ;
  RECT 2688.260 500.500 2688.460 500.700 ;
  LAYER VI3 ;
  RECT 2687.860 500.500 2688.060 500.700 ;
  LAYER VI2 ;
  RECT 2687.800 500.500 2688.660 500.780 ;
  LAYER VI2 ;
  RECT 2688.260 500.500 2688.460 500.700 ;
  LAYER VI2 ;
  RECT 2687.860 500.500 2688.060 500.700 ;
  LAYER VI3 ;
  RECT 2687.800 496.820 2688.660 497.100 ;
  LAYER VI3 ;
  RECT 2688.260 496.820 2688.460 497.020 ;
  LAYER VI3 ;
  RECT 2687.860 496.820 2688.060 497.020 ;
  LAYER VI2 ;
  RECT 2687.800 496.820 2688.660 497.100 ;
  LAYER VI2 ;
  RECT 2688.260 496.820 2688.460 497.020 ;
  LAYER VI2 ;
  RECT 2687.860 496.820 2688.060 497.020 ;
  LAYER VI3 ;
  RECT 2687.800 493.140 2688.660 493.420 ;
  LAYER VI3 ;
  RECT 2688.260 493.140 2688.460 493.340 ;
  LAYER VI3 ;
  RECT 2687.860 493.140 2688.060 493.340 ;
  LAYER VI2 ;
  RECT 2687.800 493.140 2688.660 493.420 ;
  LAYER VI2 ;
  RECT 2688.260 493.140 2688.460 493.340 ;
  LAYER VI2 ;
  RECT 2687.860 493.140 2688.060 493.340 ;
  LAYER VI3 ;
  RECT 2687.800 489.460 2688.660 489.740 ;
  LAYER VI3 ;
  RECT 2688.260 489.460 2688.460 489.660 ;
  LAYER VI3 ;
  RECT 2687.860 489.460 2688.060 489.660 ;
  LAYER VI2 ;
  RECT 2687.800 489.460 2688.660 489.740 ;
  LAYER VI2 ;
  RECT 2688.260 489.460 2688.460 489.660 ;
  LAYER VI2 ;
  RECT 2687.860 489.460 2688.060 489.660 ;
  LAYER VI3 ;
  RECT 2687.800 485.780 2688.660 486.060 ;
  LAYER VI3 ;
  RECT 2688.260 485.780 2688.460 485.980 ;
  LAYER VI3 ;
  RECT 2687.860 485.780 2688.060 485.980 ;
  LAYER VI2 ;
  RECT 2687.800 485.780 2688.660 486.060 ;
  LAYER VI2 ;
  RECT 2688.260 485.780 2688.460 485.980 ;
  LAYER VI2 ;
  RECT 2687.860 485.780 2688.060 485.980 ;
  LAYER VI3 ;
  RECT 2687.800 482.100 2688.660 482.380 ;
  LAYER VI3 ;
  RECT 2688.260 482.100 2688.460 482.300 ;
  LAYER VI3 ;
  RECT 2687.860 482.100 2688.060 482.300 ;
  LAYER VI2 ;
  RECT 2687.800 482.100 2688.660 482.380 ;
  LAYER VI2 ;
  RECT 2688.260 482.100 2688.460 482.300 ;
  LAYER VI2 ;
  RECT 2687.860 482.100 2688.060 482.300 ;
  LAYER VI3 ;
  RECT 2687.800 478.420 2688.660 478.700 ;
  LAYER VI3 ;
  RECT 2688.260 478.420 2688.460 478.620 ;
  LAYER VI3 ;
  RECT 2687.860 478.420 2688.060 478.620 ;
  LAYER VI2 ;
  RECT 2687.800 478.420 2688.660 478.700 ;
  LAYER VI2 ;
  RECT 2688.260 478.420 2688.460 478.620 ;
  LAYER VI2 ;
  RECT 2687.860 478.420 2688.060 478.620 ;
  LAYER VI3 ;
  RECT 2687.800 474.740 2688.660 475.020 ;
  LAYER VI3 ;
  RECT 2688.260 474.740 2688.460 474.940 ;
  LAYER VI3 ;
  RECT 2687.860 474.740 2688.060 474.940 ;
  LAYER VI2 ;
  RECT 2687.800 474.740 2688.660 475.020 ;
  LAYER VI2 ;
  RECT 2688.260 474.740 2688.460 474.940 ;
  LAYER VI2 ;
  RECT 2687.860 474.740 2688.060 474.940 ;
  LAYER VI3 ;
  RECT 2687.800 471.060 2688.660 471.340 ;
  LAYER VI3 ;
  RECT 2688.260 471.060 2688.460 471.260 ;
  LAYER VI3 ;
  RECT 2687.860 471.060 2688.060 471.260 ;
  LAYER VI2 ;
  RECT 2687.800 471.060 2688.660 471.340 ;
  LAYER VI2 ;
  RECT 2688.260 471.060 2688.460 471.260 ;
  LAYER VI2 ;
  RECT 2687.860 471.060 2688.060 471.260 ;
  LAYER VI3 ;
  RECT 2687.800 467.380 2688.660 467.660 ;
  LAYER VI3 ;
  RECT 2688.260 467.380 2688.460 467.580 ;
  LAYER VI3 ;
  RECT 2687.860 467.380 2688.060 467.580 ;
  LAYER VI2 ;
  RECT 2687.800 467.380 2688.660 467.660 ;
  LAYER VI2 ;
  RECT 2688.260 467.380 2688.460 467.580 ;
  LAYER VI2 ;
  RECT 2687.860 467.380 2688.060 467.580 ;
  LAYER VI3 ;
  RECT 2687.800 463.700 2688.660 463.980 ;
  LAYER VI3 ;
  RECT 2688.260 463.700 2688.460 463.900 ;
  LAYER VI3 ;
  RECT 2687.860 463.700 2688.060 463.900 ;
  LAYER VI2 ;
  RECT 2687.800 463.700 2688.660 463.980 ;
  LAYER VI2 ;
  RECT 2688.260 463.700 2688.460 463.900 ;
  LAYER VI2 ;
  RECT 2687.860 463.700 2688.060 463.900 ;
  LAYER VI3 ;
  RECT 2687.800 460.020 2688.660 460.300 ;
  LAYER VI3 ;
  RECT 2688.260 460.020 2688.460 460.220 ;
  LAYER VI3 ;
  RECT 2687.860 460.020 2688.060 460.220 ;
  LAYER VI2 ;
  RECT 2687.800 460.020 2688.660 460.300 ;
  LAYER VI2 ;
  RECT 2688.260 460.020 2688.460 460.220 ;
  LAYER VI2 ;
  RECT 2687.860 460.020 2688.060 460.220 ;
  LAYER VI3 ;
  RECT 2687.800 456.340 2688.660 456.620 ;
  LAYER VI3 ;
  RECT 2688.260 456.340 2688.460 456.540 ;
  LAYER VI3 ;
  RECT 2687.860 456.340 2688.060 456.540 ;
  LAYER VI2 ;
  RECT 2687.800 456.340 2688.660 456.620 ;
  LAYER VI2 ;
  RECT 2688.260 456.340 2688.460 456.540 ;
  LAYER VI2 ;
  RECT 2687.860 456.340 2688.060 456.540 ;
  LAYER VI3 ;
  RECT 2687.800 452.660 2688.660 452.940 ;
  LAYER VI3 ;
  RECT 2688.260 452.660 2688.460 452.860 ;
  LAYER VI3 ;
  RECT 2687.860 452.660 2688.060 452.860 ;
  LAYER VI2 ;
  RECT 2687.800 452.660 2688.660 452.940 ;
  LAYER VI2 ;
  RECT 2688.260 452.660 2688.460 452.860 ;
  LAYER VI2 ;
  RECT 2687.860 452.660 2688.060 452.860 ;
  LAYER VI3 ;
  RECT 2687.800 448.980 2688.660 449.260 ;
  LAYER VI3 ;
  RECT 2688.260 448.980 2688.460 449.180 ;
  LAYER VI3 ;
  RECT 2687.860 448.980 2688.060 449.180 ;
  LAYER VI2 ;
  RECT 2687.800 448.980 2688.660 449.260 ;
  LAYER VI2 ;
  RECT 2688.260 448.980 2688.460 449.180 ;
  LAYER VI2 ;
  RECT 2687.860 448.980 2688.060 449.180 ;
  LAYER VI3 ;
  RECT 2687.800 445.300 2688.660 445.580 ;
  LAYER VI3 ;
  RECT 2688.260 445.300 2688.460 445.500 ;
  LAYER VI3 ;
  RECT 2687.860 445.300 2688.060 445.500 ;
  LAYER VI2 ;
  RECT 2687.800 445.300 2688.660 445.580 ;
  LAYER VI2 ;
  RECT 2688.260 445.300 2688.460 445.500 ;
  LAYER VI2 ;
  RECT 2687.860 445.300 2688.060 445.500 ;
  LAYER VI3 ;
  RECT 2687.800 441.620 2688.660 441.900 ;
  LAYER VI3 ;
  RECT 2688.260 441.620 2688.460 441.820 ;
  LAYER VI3 ;
  RECT 2687.860 441.620 2688.060 441.820 ;
  LAYER VI2 ;
  RECT 2687.800 441.620 2688.660 441.900 ;
  LAYER VI2 ;
  RECT 2688.260 441.620 2688.460 441.820 ;
  LAYER VI2 ;
  RECT 2687.860 441.620 2688.060 441.820 ;
  LAYER VI3 ;
  RECT 2687.800 437.940 2688.660 438.220 ;
  LAYER VI3 ;
  RECT 2688.260 437.940 2688.460 438.140 ;
  LAYER VI3 ;
  RECT 2687.860 437.940 2688.060 438.140 ;
  LAYER VI2 ;
  RECT 2687.800 437.940 2688.660 438.220 ;
  LAYER VI2 ;
  RECT 2688.260 437.940 2688.460 438.140 ;
  LAYER VI2 ;
  RECT 2687.860 437.940 2688.060 438.140 ;
  LAYER VI3 ;
  RECT 2687.800 434.260 2688.660 434.540 ;
  LAYER VI3 ;
  RECT 2688.260 434.260 2688.460 434.460 ;
  LAYER VI3 ;
  RECT 2687.860 434.260 2688.060 434.460 ;
  LAYER VI2 ;
  RECT 2687.800 434.260 2688.660 434.540 ;
  LAYER VI2 ;
  RECT 2688.260 434.260 2688.460 434.460 ;
  LAYER VI2 ;
  RECT 2687.860 434.260 2688.060 434.460 ;
  LAYER VI3 ;
  RECT 2687.800 430.580 2688.660 430.860 ;
  LAYER VI3 ;
  RECT 2688.260 430.580 2688.460 430.780 ;
  LAYER VI3 ;
  RECT 2687.860 430.580 2688.060 430.780 ;
  LAYER VI2 ;
  RECT 2687.800 430.580 2688.660 430.860 ;
  LAYER VI2 ;
  RECT 2688.260 430.580 2688.460 430.780 ;
  LAYER VI2 ;
  RECT 2687.860 430.580 2688.060 430.780 ;
  LAYER VI3 ;
  RECT 2687.800 426.900 2688.660 427.180 ;
  LAYER VI3 ;
  RECT 2688.260 426.900 2688.460 427.100 ;
  LAYER VI3 ;
  RECT 2687.860 426.900 2688.060 427.100 ;
  LAYER VI2 ;
  RECT 2687.800 426.900 2688.660 427.180 ;
  LAYER VI2 ;
  RECT 2688.260 426.900 2688.460 427.100 ;
  LAYER VI2 ;
  RECT 2687.860 426.900 2688.060 427.100 ;
  LAYER VI3 ;
  RECT 2687.800 423.220 2688.660 423.500 ;
  LAYER VI3 ;
  RECT 2688.260 423.220 2688.460 423.420 ;
  LAYER VI3 ;
  RECT 2687.860 423.220 2688.060 423.420 ;
  LAYER VI2 ;
  RECT 2687.800 423.220 2688.660 423.500 ;
  LAYER VI2 ;
  RECT 2688.260 423.220 2688.460 423.420 ;
  LAYER VI2 ;
  RECT 2687.860 423.220 2688.060 423.420 ;
  LAYER VI3 ;
  RECT 2687.800 419.540 2688.660 419.820 ;
  LAYER VI3 ;
  RECT 2688.260 419.540 2688.460 419.740 ;
  LAYER VI3 ;
  RECT 2687.860 419.540 2688.060 419.740 ;
  LAYER VI2 ;
  RECT 2687.800 419.540 2688.660 419.820 ;
  LAYER VI2 ;
  RECT 2688.260 419.540 2688.460 419.740 ;
  LAYER VI2 ;
  RECT 2687.860 419.540 2688.060 419.740 ;
  LAYER VI3 ;
  RECT 2687.800 415.860 2688.660 416.140 ;
  LAYER VI3 ;
  RECT 2688.260 415.860 2688.460 416.060 ;
  LAYER VI3 ;
  RECT 2687.860 415.860 2688.060 416.060 ;
  LAYER VI2 ;
  RECT 2687.800 415.860 2688.660 416.140 ;
  LAYER VI2 ;
  RECT 2688.260 415.860 2688.460 416.060 ;
  LAYER VI2 ;
  RECT 2687.860 415.860 2688.060 416.060 ;
  LAYER VI3 ;
  RECT 2687.800 412.180 2688.660 412.460 ;
  LAYER VI3 ;
  RECT 2688.260 412.180 2688.460 412.380 ;
  LAYER VI3 ;
  RECT 2687.860 412.180 2688.060 412.380 ;
  LAYER VI2 ;
  RECT 2687.800 412.180 2688.660 412.460 ;
  LAYER VI2 ;
  RECT 2688.260 412.180 2688.460 412.380 ;
  LAYER VI2 ;
  RECT 2687.860 412.180 2688.060 412.380 ;
  LAYER VI3 ;
  RECT 2687.800 408.500 2688.660 408.780 ;
  LAYER VI3 ;
  RECT 2688.260 408.500 2688.460 408.700 ;
  LAYER VI3 ;
  RECT 2687.860 408.500 2688.060 408.700 ;
  LAYER VI2 ;
  RECT 2687.800 408.500 2688.660 408.780 ;
  LAYER VI2 ;
  RECT 2688.260 408.500 2688.460 408.700 ;
  LAYER VI2 ;
  RECT 2687.860 408.500 2688.060 408.700 ;
  LAYER VI3 ;
  RECT 2687.800 404.820 2688.660 405.100 ;
  LAYER VI3 ;
  RECT 2688.260 404.820 2688.460 405.020 ;
  LAYER VI3 ;
  RECT 2687.860 404.820 2688.060 405.020 ;
  LAYER VI2 ;
  RECT 2687.800 404.820 2688.660 405.100 ;
  LAYER VI2 ;
  RECT 2688.260 404.820 2688.460 405.020 ;
  LAYER VI2 ;
  RECT 2687.860 404.820 2688.060 405.020 ;
  LAYER VI3 ;
  RECT 2687.800 401.140 2688.660 401.420 ;
  LAYER VI3 ;
  RECT 2688.260 401.140 2688.460 401.340 ;
  LAYER VI3 ;
  RECT 2687.860 401.140 2688.060 401.340 ;
  LAYER VI2 ;
  RECT 2687.800 401.140 2688.660 401.420 ;
  LAYER VI2 ;
  RECT 2688.260 401.140 2688.460 401.340 ;
  LAYER VI2 ;
  RECT 2687.860 401.140 2688.060 401.340 ;
  LAYER VI3 ;
  RECT 2687.800 397.460 2688.660 397.740 ;
  LAYER VI3 ;
  RECT 2688.260 397.460 2688.460 397.660 ;
  LAYER VI3 ;
  RECT 2687.860 397.460 2688.060 397.660 ;
  LAYER VI2 ;
  RECT 2687.800 397.460 2688.660 397.740 ;
  LAYER VI2 ;
  RECT 2688.260 397.460 2688.460 397.660 ;
  LAYER VI2 ;
  RECT 2687.860 397.460 2688.060 397.660 ;
  LAYER VI3 ;
  RECT 2687.800 393.780 2688.660 394.060 ;
  LAYER VI3 ;
  RECT 2688.260 393.780 2688.460 393.980 ;
  LAYER VI3 ;
  RECT 2687.860 393.780 2688.060 393.980 ;
  LAYER VI2 ;
  RECT 2687.800 393.780 2688.660 394.060 ;
  LAYER VI2 ;
  RECT 2688.260 393.780 2688.460 393.980 ;
  LAYER VI2 ;
  RECT 2687.860 393.780 2688.060 393.980 ;
  LAYER VI3 ;
  RECT 2687.800 390.100 2688.660 390.380 ;
  LAYER VI3 ;
  RECT 2688.260 390.100 2688.460 390.300 ;
  LAYER VI3 ;
  RECT 2687.860 390.100 2688.060 390.300 ;
  LAYER VI2 ;
  RECT 2687.800 390.100 2688.660 390.380 ;
  LAYER VI2 ;
  RECT 2688.260 390.100 2688.460 390.300 ;
  LAYER VI2 ;
  RECT 2687.860 390.100 2688.060 390.300 ;
  LAYER VI3 ;
  RECT 2687.800 386.420 2688.660 386.700 ;
  LAYER VI3 ;
  RECT 2688.260 386.420 2688.460 386.620 ;
  LAYER VI3 ;
  RECT 2687.860 386.420 2688.060 386.620 ;
  LAYER VI2 ;
  RECT 2687.800 386.420 2688.660 386.700 ;
  LAYER VI2 ;
  RECT 2688.260 386.420 2688.460 386.620 ;
  LAYER VI2 ;
  RECT 2687.860 386.420 2688.060 386.620 ;
  LAYER VI3 ;
  RECT 2687.800 382.740 2688.660 383.020 ;
  LAYER VI3 ;
  RECT 2688.260 382.740 2688.460 382.940 ;
  LAYER VI3 ;
  RECT 2687.860 382.740 2688.060 382.940 ;
  LAYER VI2 ;
  RECT 2687.800 382.740 2688.660 383.020 ;
  LAYER VI2 ;
  RECT 2688.260 382.740 2688.460 382.940 ;
  LAYER VI2 ;
  RECT 2687.860 382.740 2688.060 382.940 ;
  LAYER VI3 ;
  RECT 2687.800 379.060 2688.660 379.340 ;
  LAYER VI3 ;
  RECT 2688.260 379.060 2688.460 379.260 ;
  LAYER VI3 ;
  RECT 2687.860 379.060 2688.060 379.260 ;
  LAYER VI2 ;
  RECT 2687.800 379.060 2688.660 379.340 ;
  LAYER VI2 ;
  RECT 2688.260 379.060 2688.460 379.260 ;
  LAYER VI2 ;
  RECT 2687.860 379.060 2688.060 379.260 ;
  LAYER VI3 ;
  RECT 2687.800 375.380 2688.660 375.660 ;
  LAYER VI3 ;
  RECT 2688.260 375.380 2688.460 375.580 ;
  LAYER VI3 ;
  RECT 2687.860 375.380 2688.060 375.580 ;
  LAYER VI2 ;
  RECT 2687.800 375.380 2688.660 375.660 ;
  LAYER VI2 ;
  RECT 2688.260 375.380 2688.460 375.580 ;
  LAYER VI2 ;
  RECT 2687.860 375.380 2688.060 375.580 ;
  LAYER VI3 ;
  RECT 2687.800 371.700 2688.660 371.980 ;
  LAYER VI3 ;
  RECT 2688.260 371.700 2688.460 371.900 ;
  LAYER VI3 ;
  RECT 2687.860 371.700 2688.060 371.900 ;
  LAYER VI2 ;
  RECT 2687.800 371.700 2688.660 371.980 ;
  LAYER VI2 ;
  RECT 2688.260 371.700 2688.460 371.900 ;
  LAYER VI2 ;
  RECT 2687.860 371.700 2688.060 371.900 ;
  LAYER VI3 ;
  RECT 2687.800 368.020 2688.660 368.300 ;
  LAYER VI3 ;
  RECT 2688.260 368.020 2688.460 368.220 ;
  LAYER VI3 ;
  RECT 2687.860 368.020 2688.060 368.220 ;
  LAYER VI2 ;
  RECT 2687.800 368.020 2688.660 368.300 ;
  LAYER VI2 ;
  RECT 2688.260 368.020 2688.460 368.220 ;
  LAYER VI2 ;
  RECT 2687.860 368.020 2688.060 368.220 ;
  LAYER VI3 ;
  RECT 2687.800 364.340 2688.660 364.620 ;
  LAYER VI3 ;
  RECT 2688.260 364.340 2688.460 364.540 ;
  LAYER VI3 ;
  RECT 2687.860 364.340 2688.060 364.540 ;
  LAYER VI2 ;
  RECT 2687.800 364.340 2688.660 364.620 ;
  LAYER VI2 ;
  RECT 2688.260 364.340 2688.460 364.540 ;
  LAYER VI2 ;
  RECT 2687.860 364.340 2688.060 364.540 ;
  LAYER VI3 ;
  RECT 2687.800 360.660 2688.660 360.940 ;
  LAYER VI3 ;
  RECT 2688.260 360.660 2688.460 360.860 ;
  LAYER VI3 ;
  RECT 2687.860 360.660 2688.060 360.860 ;
  LAYER VI2 ;
  RECT 2687.800 360.660 2688.660 360.940 ;
  LAYER VI2 ;
  RECT 2688.260 360.660 2688.460 360.860 ;
  LAYER VI2 ;
  RECT 2687.860 360.660 2688.060 360.860 ;
  LAYER VI3 ;
  RECT 2687.800 356.980 2688.660 357.260 ;
  LAYER VI3 ;
  RECT 2688.260 356.980 2688.460 357.180 ;
  LAYER VI3 ;
  RECT 2687.860 356.980 2688.060 357.180 ;
  LAYER VI2 ;
  RECT 2687.800 356.980 2688.660 357.260 ;
  LAYER VI2 ;
  RECT 2688.260 356.980 2688.460 357.180 ;
  LAYER VI2 ;
  RECT 2687.860 356.980 2688.060 357.180 ;
  LAYER VI3 ;
  RECT 2687.800 353.300 2688.660 353.580 ;
  LAYER VI3 ;
  RECT 2688.260 353.300 2688.460 353.500 ;
  LAYER VI3 ;
  RECT 2687.860 353.300 2688.060 353.500 ;
  LAYER VI2 ;
  RECT 2687.800 353.300 2688.660 353.580 ;
  LAYER VI2 ;
  RECT 2688.260 353.300 2688.460 353.500 ;
  LAYER VI2 ;
  RECT 2687.860 353.300 2688.060 353.500 ;
  LAYER VI3 ;
  RECT 2687.800 349.620 2688.660 349.900 ;
  LAYER VI3 ;
  RECT 2688.260 349.620 2688.460 349.820 ;
  LAYER VI3 ;
  RECT 2687.860 349.620 2688.060 349.820 ;
  LAYER VI2 ;
  RECT 2687.800 349.620 2688.660 349.900 ;
  LAYER VI2 ;
  RECT 2688.260 349.620 2688.460 349.820 ;
  LAYER VI2 ;
  RECT 2687.860 349.620 2688.060 349.820 ;
  LAYER VI3 ;
  RECT 2687.800 345.940 2688.660 346.220 ;
  LAYER VI3 ;
  RECT 2688.260 345.940 2688.460 346.140 ;
  LAYER VI3 ;
  RECT 2687.860 345.940 2688.060 346.140 ;
  LAYER VI2 ;
  RECT 2687.800 345.940 2688.660 346.220 ;
  LAYER VI2 ;
  RECT 2688.260 345.940 2688.460 346.140 ;
  LAYER VI2 ;
  RECT 2687.860 345.940 2688.060 346.140 ;
  LAYER VI3 ;
  RECT 2687.800 342.260 2688.660 342.540 ;
  LAYER VI3 ;
  RECT 2688.260 342.260 2688.460 342.460 ;
  LAYER VI3 ;
  RECT 2687.860 342.260 2688.060 342.460 ;
  LAYER VI2 ;
  RECT 2687.800 342.260 2688.660 342.540 ;
  LAYER VI2 ;
  RECT 2688.260 342.260 2688.460 342.460 ;
  LAYER VI2 ;
  RECT 2687.860 342.260 2688.060 342.460 ;
  LAYER VI3 ;
  RECT 2687.800 338.580 2688.660 338.860 ;
  LAYER VI3 ;
  RECT 2688.260 338.580 2688.460 338.780 ;
  LAYER VI3 ;
  RECT 2687.860 338.580 2688.060 338.780 ;
  LAYER VI2 ;
  RECT 2687.800 338.580 2688.660 338.860 ;
  LAYER VI2 ;
  RECT 2688.260 338.580 2688.460 338.780 ;
  LAYER VI2 ;
  RECT 2687.860 338.580 2688.060 338.780 ;
  LAYER VI3 ;
  RECT 2687.800 334.900 2688.660 335.180 ;
  LAYER VI3 ;
  RECT 2688.260 334.900 2688.460 335.100 ;
  LAYER VI3 ;
  RECT 2687.860 334.900 2688.060 335.100 ;
  LAYER VI2 ;
  RECT 2687.800 334.900 2688.660 335.180 ;
  LAYER VI2 ;
  RECT 2688.260 334.900 2688.460 335.100 ;
  LAYER VI2 ;
  RECT 2687.860 334.900 2688.060 335.100 ;
  LAYER VI3 ;
  RECT 2687.800 331.220 2688.660 331.500 ;
  LAYER VI3 ;
  RECT 2688.260 331.220 2688.460 331.420 ;
  LAYER VI3 ;
  RECT 2687.860 331.220 2688.060 331.420 ;
  LAYER VI2 ;
  RECT 2687.800 331.220 2688.660 331.500 ;
  LAYER VI2 ;
  RECT 2688.260 331.220 2688.460 331.420 ;
  LAYER VI2 ;
  RECT 2687.860 331.220 2688.060 331.420 ;
  LAYER VI3 ;
  RECT 2687.800 327.540 2688.660 327.820 ;
  LAYER VI3 ;
  RECT 2688.260 327.540 2688.460 327.740 ;
  LAYER VI3 ;
  RECT 2687.860 327.540 2688.060 327.740 ;
  LAYER VI2 ;
  RECT 2687.800 327.540 2688.660 327.820 ;
  LAYER VI2 ;
  RECT 2688.260 327.540 2688.460 327.740 ;
  LAYER VI2 ;
  RECT 2687.860 327.540 2688.060 327.740 ;
  LAYER VI3 ;
  RECT 2687.800 323.860 2688.660 324.140 ;
  LAYER VI3 ;
  RECT 2688.260 323.860 2688.460 324.060 ;
  LAYER VI3 ;
  RECT 2687.860 323.860 2688.060 324.060 ;
  LAYER VI2 ;
  RECT 2687.800 323.860 2688.660 324.140 ;
  LAYER VI2 ;
  RECT 2688.260 323.860 2688.460 324.060 ;
  LAYER VI2 ;
  RECT 2687.860 323.860 2688.060 324.060 ;
  LAYER VI3 ;
  RECT 2687.800 320.180 2688.660 320.460 ;
  LAYER VI3 ;
  RECT 2688.260 320.180 2688.460 320.380 ;
  LAYER VI3 ;
  RECT 2687.860 320.180 2688.060 320.380 ;
  LAYER VI2 ;
  RECT 2687.800 320.180 2688.660 320.460 ;
  LAYER VI2 ;
  RECT 2688.260 320.180 2688.460 320.380 ;
  LAYER VI2 ;
  RECT 2687.860 320.180 2688.060 320.380 ;
  LAYER VI3 ;
  RECT 2687.800 316.500 2688.660 316.780 ;
  LAYER VI3 ;
  RECT 2688.260 316.500 2688.460 316.700 ;
  LAYER VI3 ;
  RECT 2687.860 316.500 2688.060 316.700 ;
  LAYER VI2 ;
  RECT 2687.800 316.500 2688.660 316.780 ;
  LAYER VI2 ;
  RECT 2688.260 316.500 2688.460 316.700 ;
  LAYER VI2 ;
  RECT 2687.860 316.500 2688.060 316.700 ;
  LAYER VI3 ;
  RECT 2687.800 312.820 2688.660 313.100 ;
  LAYER VI3 ;
  RECT 2688.260 312.820 2688.460 313.020 ;
  LAYER VI3 ;
  RECT 2687.860 312.820 2688.060 313.020 ;
  LAYER VI2 ;
  RECT 2687.800 312.820 2688.660 313.100 ;
  LAYER VI2 ;
  RECT 2688.260 312.820 2688.460 313.020 ;
  LAYER VI2 ;
  RECT 2687.860 312.820 2688.060 313.020 ;
  LAYER VI3 ;
  RECT 2687.800 309.140 2688.660 309.420 ;
  LAYER VI3 ;
  RECT 2688.260 309.140 2688.460 309.340 ;
  LAYER VI3 ;
  RECT 2687.860 309.140 2688.060 309.340 ;
  LAYER VI2 ;
  RECT 2687.800 309.140 2688.660 309.420 ;
  LAYER VI2 ;
  RECT 2688.260 309.140 2688.460 309.340 ;
  LAYER VI2 ;
  RECT 2687.860 309.140 2688.060 309.340 ;
  LAYER VI3 ;
  RECT 2687.800 305.460 2688.660 305.740 ;
  LAYER VI3 ;
  RECT 2688.260 305.460 2688.460 305.660 ;
  LAYER VI3 ;
  RECT 2687.860 305.460 2688.060 305.660 ;
  LAYER VI2 ;
  RECT 2687.800 305.460 2688.660 305.740 ;
  LAYER VI2 ;
  RECT 2688.260 305.460 2688.460 305.660 ;
  LAYER VI2 ;
  RECT 2687.860 305.460 2688.060 305.660 ;
  LAYER VI3 ;
  RECT 2687.800 301.780 2688.660 302.060 ;
  LAYER VI3 ;
  RECT 2688.260 301.780 2688.460 301.980 ;
  LAYER VI3 ;
  RECT 2687.860 301.780 2688.060 301.980 ;
  LAYER VI2 ;
  RECT 2687.800 301.780 2688.660 302.060 ;
  LAYER VI2 ;
  RECT 2688.260 301.780 2688.460 301.980 ;
  LAYER VI2 ;
  RECT 2687.860 301.780 2688.060 301.980 ;
  LAYER VI3 ;
  RECT 2687.800 298.100 2688.660 298.380 ;
  LAYER VI3 ;
  RECT 2688.260 298.100 2688.460 298.300 ;
  LAYER VI3 ;
  RECT 2687.860 298.100 2688.060 298.300 ;
  LAYER VI2 ;
  RECT 2687.800 298.100 2688.660 298.380 ;
  LAYER VI2 ;
  RECT 2688.260 298.100 2688.460 298.300 ;
  LAYER VI2 ;
  RECT 2687.860 298.100 2688.060 298.300 ;
  LAYER VI3 ;
  RECT 2687.800 294.420 2688.660 294.700 ;
  LAYER VI3 ;
  RECT 2688.260 294.420 2688.460 294.620 ;
  LAYER VI3 ;
  RECT 2687.860 294.420 2688.060 294.620 ;
  LAYER VI2 ;
  RECT 2687.800 294.420 2688.660 294.700 ;
  LAYER VI2 ;
  RECT 2688.260 294.420 2688.460 294.620 ;
  LAYER VI2 ;
  RECT 2687.860 294.420 2688.060 294.620 ;
  LAYER VI3 ;
  RECT 2687.800 290.740 2688.660 291.020 ;
  LAYER VI3 ;
  RECT 2688.260 290.740 2688.460 290.940 ;
  LAYER VI3 ;
  RECT 2687.860 290.740 2688.060 290.940 ;
  LAYER VI2 ;
  RECT 2687.800 290.740 2688.660 291.020 ;
  LAYER VI2 ;
  RECT 2688.260 290.740 2688.460 290.940 ;
  LAYER VI2 ;
  RECT 2687.860 290.740 2688.060 290.940 ;
  LAYER VI3 ;
  RECT 2687.800 287.060 2688.660 287.340 ;
  LAYER VI3 ;
  RECT 2688.260 287.060 2688.460 287.260 ;
  LAYER VI3 ;
  RECT 2687.860 287.060 2688.060 287.260 ;
  LAYER VI2 ;
  RECT 2687.800 287.060 2688.660 287.340 ;
  LAYER VI2 ;
  RECT 2688.260 287.060 2688.460 287.260 ;
  LAYER VI2 ;
  RECT 2687.860 287.060 2688.060 287.260 ;
  LAYER VI3 ;
  RECT 2687.800 283.380 2688.660 283.660 ;
  LAYER VI3 ;
  RECT 2688.260 283.380 2688.460 283.580 ;
  LAYER VI3 ;
  RECT 2687.860 283.380 2688.060 283.580 ;
  LAYER VI2 ;
  RECT 2687.800 283.380 2688.660 283.660 ;
  LAYER VI2 ;
  RECT 2688.260 283.380 2688.460 283.580 ;
  LAYER VI2 ;
  RECT 2687.860 283.380 2688.060 283.580 ;
  LAYER VI3 ;
  RECT 2687.800 279.700 2688.660 279.980 ;
  LAYER VI3 ;
  RECT 2688.260 279.700 2688.460 279.900 ;
  LAYER VI3 ;
  RECT 2687.860 279.700 2688.060 279.900 ;
  LAYER VI2 ;
  RECT 2687.800 279.700 2688.660 279.980 ;
  LAYER VI2 ;
  RECT 2688.260 279.700 2688.460 279.900 ;
  LAYER VI2 ;
  RECT 2687.860 279.700 2688.060 279.900 ;
  LAYER VI3 ;
  RECT 2687.800 276.020 2688.660 276.300 ;
  LAYER VI3 ;
  RECT 2688.260 276.020 2688.460 276.220 ;
  LAYER VI3 ;
  RECT 2687.860 276.020 2688.060 276.220 ;
  LAYER VI2 ;
  RECT 2687.800 276.020 2688.660 276.300 ;
  LAYER VI2 ;
  RECT 2688.260 276.020 2688.460 276.220 ;
  LAYER VI2 ;
  RECT 2687.860 276.020 2688.060 276.220 ;
  LAYER VI3 ;
  RECT 2687.800 272.340 2688.660 272.620 ;
  LAYER VI3 ;
  RECT 2688.260 272.340 2688.460 272.540 ;
  LAYER VI3 ;
  RECT 2687.860 272.340 2688.060 272.540 ;
  LAYER VI2 ;
  RECT 2687.800 272.340 2688.660 272.620 ;
  LAYER VI2 ;
  RECT 2688.260 272.340 2688.460 272.540 ;
  LAYER VI2 ;
  RECT 2687.860 272.340 2688.060 272.540 ;
  LAYER VI3 ;
  RECT 2687.800 268.660 2688.660 268.940 ;
  LAYER VI3 ;
  RECT 2688.260 268.660 2688.460 268.860 ;
  LAYER VI3 ;
  RECT 2687.860 268.660 2688.060 268.860 ;
  LAYER VI2 ;
  RECT 2687.800 268.660 2688.660 268.940 ;
  LAYER VI2 ;
  RECT 2688.260 268.660 2688.460 268.860 ;
  LAYER VI2 ;
  RECT 2687.860 268.660 2688.060 268.860 ;
  LAYER VI3 ;
  RECT 2687.800 264.980 2688.660 265.260 ;
  LAYER VI3 ;
  RECT 2688.260 264.980 2688.460 265.180 ;
  LAYER VI3 ;
  RECT 2687.860 264.980 2688.060 265.180 ;
  LAYER VI2 ;
  RECT 2687.800 264.980 2688.660 265.260 ;
  LAYER VI2 ;
  RECT 2688.260 264.980 2688.460 265.180 ;
  LAYER VI2 ;
  RECT 2687.860 264.980 2688.060 265.180 ;
  LAYER VI3 ;
  RECT 2687.800 261.300 2688.660 261.580 ;
  LAYER VI3 ;
  RECT 2688.260 261.300 2688.460 261.500 ;
  LAYER VI3 ;
  RECT 2687.860 261.300 2688.060 261.500 ;
  LAYER VI2 ;
  RECT 2687.800 261.300 2688.660 261.580 ;
  LAYER VI2 ;
  RECT 2688.260 261.300 2688.460 261.500 ;
  LAYER VI2 ;
  RECT 2687.860 261.300 2688.060 261.500 ;
  LAYER VI3 ;
  RECT 2687.800 257.620 2688.660 257.900 ;
  LAYER VI3 ;
  RECT 2688.260 257.620 2688.460 257.820 ;
  LAYER VI3 ;
  RECT 2687.860 257.620 2688.060 257.820 ;
  LAYER VI2 ;
  RECT 2687.800 257.620 2688.660 257.900 ;
  LAYER VI2 ;
  RECT 2688.260 257.620 2688.460 257.820 ;
  LAYER VI2 ;
  RECT 2687.860 257.620 2688.060 257.820 ;
  LAYER VI3 ;
  RECT 2687.800 253.940 2688.660 254.220 ;
  LAYER VI3 ;
  RECT 2688.260 253.940 2688.460 254.140 ;
  LAYER VI3 ;
  RECT 2687.860 253.940 2688.060 254.140 ;
  LAYER VI2 ;
  RECT 2687.800 253.940 2688.660 254.220 ;
  LAYER VI2 ;
  RECT 2688.260 253.940 2688.460 254.140 ;
  LAYER VI2 ;
  RECT 2687.860 253.940 2688.060 254.140 ;
  LAYER VI3 ;
  RECT 2687.800 250.260 2688.660 250.540 ;
  LAYER VI3 ;
  RECT 2688.260 250.260 2688.460 250.460 ;
  LAYER VI3 ;
  RECT 2687.860 250.260 2688.060 250.460 ;
  LAYER VI2 ;
  RECT 2687.800 250.260 2688.660 250.540 ;
  LAYER VI2 ;
  RECT 2688.260 250.260 2688.460 250.460 ;
  LAYER VI2 ;
  RECT 2687.860 250.260 2688.060 250.460 ;
  LAYER VI3 ;
  RECT 2687.800 246.580 2688.660 246.860 ;
  LAYER VI3 ;
  RECT 2688.260 246.580 2688.460 246.780 ;
  LAYER VI3 ;
  RECT 2687.860 246.580 2688.060 246.780 ;
  LAYER VI2 ;
  RECT 2687.800 246.580 2688.660 246.860 ;
  LAYER VI2 ;
  RECT 2688.260 246.580 2688.460 246.780 ;
  LAYER VI2 ;
  RECT 2687.860 246.580 2688.060 246.780 ;
  LAYER VI3 ;
  RECT 2687.800 242.900 2688.660 243.180 ;
  LAYER VI3 ;
  RECT 2688.260 242.900 2688.460 243.100 ;
  LAYER VI3 ;
  RECT 2687.860 242.900 2688.060 243.100 ;
  LAYER VI2 ;
  RECT 2687.800 242.900 2688.660 243.180 ;
  LAYER VI2 ;
  RECT 2688.260 242.900 2688.460 243.100 ;
  LAYER VI2 ;
  RECT 2687.860 242.900 2688.060 243.100 ;
  LAYER VI3 ;
  RECT 2687.800 239.220 2688.660 239.500 ;
  LAYER VI3 ;
  RECT 2688.260 239.220 2688.460 239.420 ;
  LAYER VI3 ;
  RECT 2687.860 239.220 2688.060 239.420 ;
  LAYER VI2 ;
  RECT 2687.800 239.220 2688.660 239.500 ;
  LAYER VI2 ;
  RECT 2688.260 239.220 2688.460 239.420 ;
  LAYER VI2 ;
  RECT 2687.860 239.220 2688.060 239.420 ;
  LAYER VI3 ;
  RECT 2687.800 235.540 2688.660 235.820 ;
  LAYER VI3 ;
  RECT 2688.260 235.540 2688.460 235.740 ;
  LAYER VI3 ;
  RECT 2687.860 235.540 2688.060 235.740 ;
  LAYER VI2 ;
  RECT 2687.800 235.540 2688.660 235.820 ;
  LAYER VI2 ;
  RECT 2688.260 235.540 2688.460 235.740 ;
  LAYER VI2 ;
  RECT 2687.860 235.540 2688.060 235.740 ;
  LAYER VI3 ;
  RECT 2687.800 231.860 2688.660 232.140 ;
  LAYER VI3 ;
  RECT 2688.260 231.860 2688.460 232.060 ;
  LAYER VI3 ;
  RECT 2687.860 231.860 2688.060 232.060 ;
  LAYER VI2 ;
  RECT 2687.800 231.860 2688.660 232.140 ;
  LAYER VI2 ;
  RECT 2688.260 231.860 2688.460 232.060 ;
  LAYER VI2 ;
  RECT 2687.860 231.860 2688.060 232.060 ;
  LAYER VI3 ;
  RECT 2687.800 228.180 2688.660 228.460 ;
  LAYER VI3 ;
  RECT 2688.260 228.180 2688.460 228.380 ;
  LAYER VI3 ;
  RECT 2687.860 228.180 2688.060 228.380 ;
  LAYER VI2 ;
  RECT 2687.800 228.180 2688.660 228.460 ;
  LAYER VI2 ;
  RECT 2688.260 228.180 2688.460 228.380 ;
  LAYER VI2 ;
  RECT 2687.860 228.180 2688.060 228.380 ;
  LAYER VI3 ;
  RECT 2687.800 224.500 2688.660 224.780 ;
  LAYER VI3 ;
  RECT 2688.260 224.500 2688.460 224.700 ;
  LAYER VI3 ;
  RECT 2687.860 224.500 2688.060 224.700 ;
  LAYER VI2 ;
  RECT 2687.800 224.500 2688.660 224.780 ;
  LAYER VI2 ;
  RECT 2688.260 224.500 2688.460 224.700 ;
  LAYER VI2 ;
  RECT 2687.860 224.500 2688.060 224.700 ;
  LAYER VI3 ;
  RECT 2687.800 220.820 2688.660 221.100 ;
  LAYER VI3 ;
  RECT 2688.260 220.820 2688.460 221.020 ;
  LAYER VI3 ;
  RECT 2687.860 220.820 2688.060 221.020 ;
  LAYER VI2 ;
  RECT 2687.800 220.820 2688.660 221.100 ;
  LAYER VI2 ;
  RECT 2688.260 220.820 2688.460 221.020 ;
  LAYER VI2 ;
  RECT 2687.860 220.820 2688.060 221.020 ;
  LAYER VI3 ;
  RECT 2687.800 217.140 2688.660 217.420 ;
  LAYER VI3 ;
  RECT 2688.260 217.140 2688.460 217.340 ;
  LAYER VI3 ;
  RECT 2687.860 217.140 2688.060 217.340 ;
  LAYER VI2 ;
  RECT 2687.800 217.140 2688.660 217.420 ;
  LAYER VI2 ;
  RECT 2688.260 217.140 2688.460 217.340 ;
  LAYER VI2 ;
  RECT 2687.860 217.140 2688.060 217.340 ;
  LAYER VI3 ;
  RECT 2687.800 213.460 2688.660 213.740 ;
  LAYER VI3 ;
  RECT 2688.260 213.460 2688.460 213.660 ;
  LAYER VI3 ;
  RECT 2687.860 213.460 2688.060 213.660 ;
  LAYER VI2 ;
  RECT 2687.800 213.460 2688.660 213.740 ;
  LAYER VI2 ;
  RECT 2688.260 213.460 2688.460 213.660 ;
  LAYER VI2 ;
  RECT 2687.860 213.460 2688.060 213.660 ;
  LAYER VI3 ;
  RECT 2687.800 209.780 2688.660 210.060 ;
  LAYER VI3 ;
  RECT 2688.260 209.780 2688.460 209.980 ;
  LAYER VI3 ;
  RECT 2687.860 209.780 2688.060 209.980 ;
  LAYER VI2 ;
  RECT 2687.800 209.780 2688.660 210.060 ;
  LAYER VI2 ;
  RECT 2688.260 209.780 2688.460 209.980 ;
  LAYER VI2 ;
  RECT 2687.860 209.780 2688.060 209.980 ;
  LAYER VI3 ;
  RECT 2687.800 206.100 2688.660 206.380 ;
  LAYER VI3 ;
  RECT 2688.260 206.100 2688.460 206.300 ;
  LAYER VI3 ;
  RECT 2687.860 206.100 2688.060 206.300 ;
  LAYER VI2 ;
  RECT 2687.800 206.100 2688.660 206.380 ;
  LAYER VI2 ;
  RECT 2688.260 206.100 2688.460 206.300 ;
  LAYER VI2 ;
  RECT 2687.860 206.100 2688.060 206.300 ;
  LAYER VI3 ;
  RECT 2687.800 202.420 2688.660 202.700 ;
  LAYER VI3 ;
  RECT 2688.260 202.420 2688.460 202.620 ;
  LAYER VI3 ;
  RECT 2687.860 202.420 2688.060 202.620 ;
  LAYER VI2 ;
  RECT 2687.800 202.420 2688.660 202.700 ;
  LAYER VI2 ;
  RECT 2688.260 202.420 2688.460 202.620 ;
  LAYER VI2 ;
  RECT 2687.860 202.420 2688.060 202.620 ;
  LAYER VI3 ;
  RECT 2687.800 198.740 2688.660 199.020 ;
  LAYER VI3 ;
  RECT 2688.260 198.740 2688.460 198.940 ;
  LAYER VI3 ;
  RECT 2687.860 198.740 2688.060 198.940 ;
  LAYER VI2 ;
  RECT 2687.800 198.740 2688.660 199.020 ;
  LAYER VI2 ;
  RECT 2688.260 198.740 2688.460 198.940 ;
  LAYER VI2 ;
  RECT 2687.860 198.740 2688.060 198.940 ;
  LAYER VI3 ;
  RECT 2687.800 195.060 2688.660 195.340 ;
  LAYER VI3 ;
  RECT 2688.260 195.060 2688.460 195.260 ;
  LAYER VI3 ;
  RECT 2687.860 195.060 2688.060 195.260 ;
  LAYER VI2 ;
  RECT 2687.800 195.060 2688.660 195.340 ;
  LAYER VI2 ;
  RECT 2688.260 195.060 2688.460 195.260 ;
  LAYER VI2 ;
  RECT 2687.860 195.060 2688.060 195.260 ;
  LAYER VI3 ;
  RECT 2687.800 191.380 2688.660 191.660 ;
  LAYER VI3 ;
  RECT 2688.260 191.380 2688.460 191.580 ;
  LAYER VI3 ;
  RECT 2687.860 191.380 2688.060 191.580 ;
  LAYER VI2 ;
  RECT 2687.800 191.380 2688.660 191.660 ;
  LAYER VI2 ;
  RECT 2688.260 191.380 2688.460 191.580 ;
  LAYER VI2 ;
  RECT 2687.860 191.380 2688.060 191.580 ;
  LAYER VI3 ;
  RECT 2687.800 187.700 2688.660 187.980 ;
  LAYER VI3 ;
  RECT 2688.260 187.700 2688.460 187.900 ;
  LAYER VI3 ;
  RECT 2687.860 187.700 2688.060 187.900 ;
  LAYER VI2 ;
  RECT 2687.800 187.700 2688.660 187.980 ;
  LAYER VI2 ;
  RECT 2688.260 187.700 2688.460 187.900 ;
  LAYER VI2 ;
  RECT 2687.860 187.700 2688.060 187.900 ;
  LAYER VI3 ;
  RECT 2687.800 184.020 2688.660 184.300 ;
  LAYER VI3 ;
  RECT 2688.260 184.020 2688.460 184.220 ;
  LAYER VI3 ;
  RECT 2687.860 184.020 2688.060 184.220 ;
  LAYER VI2 ;
  RECT 2687.800 184.020 2688.660 184.300 ;
  LAYER VI2 ;
  RECT 2688.260 184.020 2688.460 184.220 ;
  LAYER VI2 ;
  RECT 2687.860 184.020 2688.060 184.220 ;
  LAYER VI3 ;
  RECT 2687.800 180.340 2688.660 180.620 ;
  LAYER VI3 ;
  RECT 2688.260 180.340 2688.460 180.540 ;
  LAYER VI3 ;
  RECT 2687.860 180.340 2688.060 180.540 ;
  LAYER VI2 ;
  RECT 2687.800 180.340 2688.660 180.620 ;
  LAYER VI2 ;
  RECT 2688.260 180.340 2688.460 180.540 ;
  LAYER VI2 ;
  RECT 2687.860 180.340 2688.060 180.540 ;
  LAYER VI3 ;
  RECT 2687.800 176.660 2688.660 176.940 ;
  LAYER VI3 ;
  RECT 2688.260 176.660 2688.460 176.860 ;
  LAYER VI3 ;
  RECT 2687.860 176.660 2688.060 176.860 ;
  LAYER VI2 ;
  RECT 2687.800 176.660 2688.660 176.940 ;
  LAYER VI2 ;
  RECT 2688.260 176.660 2688.460 176.860 ;
  LAYER VI2 ;
  RECT 2687.860 176.660 2688.060 176.860 ;
  LAYER VI3 ;
  RECT 2687.800 172.980 2688.660 173.260 ;
  LAYER VI3 ;
  RECT 2688.260 172.980 2688.460 173.180 ;
  LAYER VI3 ;
  RECT 2687.860 172.980 2688.060 173.180 ;
  LAYER VI2 ;
  RECT 2687.800 172.980 2688.660 173.260 ;
  LAYER VI2 ;
  RECT 2688.260 172.980 2688.460 173.180 ;
  LAYER VI2 ;
  RECT 2687.860 172.980 2688.060 173.180 ;
  LAYER VI3 ;
  RECT 2687.800 169.300 2688.660 169.580 ;
  LAYER VI3 ;
  RECT 2688.260 169.300 2688.460 169.500 ;
  LAYER VI3 ;
  RECT 2687.860 169.300 2688.060 169.500 ;
  LAYER VI2 ;
  RECT 2687.800 169.300 2688.660 169.580 ;
  LAYER VI2 ;
  RECT 2688.260 169.300 2688.460 169.500 ;
  LAYER VI2 ;
  RECT 2687.860 169.300 2688.060 169.500 ;
  LAYER VI3 ;
  RECT 2687.800 165.620 2688.660 165.900 ;
  LAYER VI3 ;
  RECT 2688.260 165.620 2688.460 165.820 ;
  LAYER VI3 ;
  RECT 2687.860 165.620 2688.060 165.820 ;
  LAYER VI2 ;
  RECT 2687.800 165.620 2688.660 165.900 ;
  LAYER VI2 ;
  RECT 2688.260 165.620 2688.460 165.820 ;
  LAYER VI2 ;
  RECT 2687.860 165.620 2688.060 165.820 ;
  LAYER VI3 ;
  RECT 2687.800 161.940 2688.660 162.220 ;
  LAYER VI3 ;
  RECT 2688.260 161.940 2688.460 162.140 ;
  LAYER VI3 ;
  RECT 2687.860 161.940 2688.060 162.140 ;
  LAYER VI2 ;
  RECT 2687.800 161.940 2688.660 162.220 ;
  LAYER VI2 ;
  RECT 2688.260 161.940 2688.460 162.140 ;
  LAYER VI2 ;
  RECT 2687.860 161.940 2688.060 162.140 ;
  LAYER VI3 ;
  RECT 2687.800 158.260 2688.660 158.540 ;
  LAYER VI3 ;
  RECT 2688.260 158.260 2688.460 158.460 ;
  LAYER VI3 ;
  RECT 2687.860 158.260 2688.060 158.460 ;
  LAYER VI2 ;
  RECT 2687.800 158.260 2688.660 158.540 ;
  LAYER VI2 ;
  RECT 2688.260 158.260 2688.460 158.460 ;
  LAYER VI2 ;
  RECT 2687.860 158.260 2688.060 158.460 ;
  LAYER VI3 ;
  RECT 2687.800 154.580 2688.660 154.860 ;
  LAYER VI3 ;
  RECT 2688.260 154.580 2688.460 154.780 ;
  LAYER VI3 ;
  RECT 2687.860 154.580 2688.060 154.780 ;
  LAYER VI2 ;
  RECT 2687.800 154.580 2688.660 154.860 ;
  LAYER VI2 ;
  RECT 2688.260 154.580 2688.460 154.780 ;
  LAYER VI2 ;
  RECT 2687.860 154.580 2688.060 154.780 ;
  LAYER VI3 ;
  RECT 2687.800 150.900 2688.660 151.180 ;
  LAYER VI3 ;
  RECT 2688.260 150.900 2688.460 151.100 ;
  LAYER VI3 ;
  RECT 2687.860 150.900 2688.060 151.100 ;
  LAYER VI2 ;
  RECT 2687.800 150.900 2688.660 151.180 ;
  LAYER VI2 ;
  RECT 2688.260 150.900 2688.460 151.100 ;
  LAYER VI2 ;
  RECT 2687.860 150.900 2688.060 151.100 ;
  LAYER VI3 ;
  RECT 2687.800 147.220 2688.660 147.500 ;
  LAYER VI3 ;
  RECT 2688.260 147.220 2688.460 147.420 ;
  LAYER VI3 ;
  RECT 2687.860 147.220 2688.060 147.420 ;
  LAYER VI2 ;
  RECT 2687.800 147.220 2688.660 147.500 ;
  LAYER VI2 ;
  RECT 2688.260 147.220 2688.460 147.420 ;
  LAYER VI2 ;
  RECT 2687.860 147.220 2688.060 147.420 ;
  LAYER VI3 ;
  RECT 2687.800 143.540 2688.660 143.820 ;
  LAYER VI3 ;
  RECT 2688.260 143.540 2688.460 143.740 ;
  LAYER VI3 ;
  RECT 2687.860 143.540 2688.060 143.740 ;
  LAYER VI2 ;
  RECT 2687.800 143.540 2688.660 143.820 ;
  LAYER VI2 ;
  RECT 2688.260 143.540 2688.460 143.740 ;
  LAYER VI2 ;
  RECT 2687.860 143.540 2688.060 143.740 ;
  LAYER VI3 ;
  RECT 2687.800 139.860 2688.660 140.140 ;
  LAYER VI3 ;
  RECT 2688.260 139.860 2688.460 140.060 ;
  LAYER VI3 ;
  RECT 2687.860 139.860 2688.060 140.060 ;
  LAYER VI2 ;
  RECT 2687.800 139.860 2688.660 140.140 ;
  LAYER VI2 ;
  RECT 2688.260 139.860 2688.460 140.060 ;
  LAYER VI2 ;
  RECT 2687.860 139.860 2688.060 140.060 ;
  LAYER VI3 ;
  RECT 2687.800 136.180 2688.660 136.460 ;
  LAYER VI3 ;
  RECT 2688.260 136.180 2688.460 136.380 ;
  LAYER VI3 ;
  RECT 2687.860 136.180 2688.060 136.380 ;
  LAYER VI2 ;
  RECT 2687.800 136.180 2688.660 136.460 ;
  LAYER VI2 ;
  RECT 2688.260 136.180 2688.460 136.380 ;
  LAYER VI2 ;
  RECT 2687.860 136.180 2688.060 136.380 ;
  LAYER VI3 ;
  RECT 2687.800 132.500 2688.660 132.780 ;
  LAYER VI3 ;
  RECT 2688.260 132.500 2688.460 132.700 ;
  LAYER VI3 ;
  RECT 2687.860 132.500 2688.060 132.700 ;
  LAYER VI2 ;
  RECT 2687.800 132.500 2688.660 132.780 ;
  LAYER VI2 ;
  RECT 2688.260 132.500 2688.460 132.700 ;
  LAYER VI2 ;
  RECT 2687.860 132.500 2688.060 132.700 ;
  LAYER VI3 ;
  RECT 2687.800 128.820 2688.660 129.100 ;
  LAYER VI3 ;
  RECT 2688.260 128.820 2688.460 129.020 ;
  LAYER VI3 ;
  RECT 2687.860 128.820 2688.060 129.020 ;
  LAYER VI2 ;
  RECT 2687.800 128.820 2688.660 129.100 ;
  LAYER VI2 ;
  RECT 2688.260 128.820 2688.460 129.020 ;
  LAYER VI2 ;
  RECT 2687.860 128.820 2688.060 129.020 ;
  LAYER VI3 ;
  RECT 2687.800 125.140 2688.660 125.420 ;
  LAYER VI3 ;
  RECT 2688.260 125.140 2688.460 125.340 ;
  LAYER VI3 ;
  RECT 2687.860 125.140 2688.060 125.340 ;
  LAYER VI2 ;
  RECT 2687.800 125.140 2688.660 125.420 ;
  LAYER VI2 ;
  RECT 2688.260 125.140 2688.460 125.340 ;
  LAYER VI2 ;
  RECT 2687.860 125.140 2688.060 125.340 ;
  LAYER VI3 ;
  RECT 2687.800 121.460 2688.660 121.740 ;
  LAYER VI3 ;
  RECT 2688.260 121.460 2688.460 121.660 ;
  LAYER VI3 ;
  RECT 2687.860 121.460 2688.060 121.660 ;
  LAYER VI2 ;
  RECT 2687.800 121.460 2688.660 121.740 ;
  LAYER VI2 ;
  RECT 2688.260 121.460 2688.460 121.660 ;
  LAYER VI2 ;
  RECT 2687.860 121.460 2688.060 121.660 ;
  LAYER VI3 ;
  RECT 2687.800 117.780 2688.660 118.060 ;
  LAYER VI3 ;
  RECT 2688.260 117.780 2688.460 117.980 ;
  LAYER VI3 ;
  RECT 2687.860 117.780 2688.060 117.980 ;
  LAYER VI2 ;
  RECT 2687.800 117.780 2688.660 118.060 ;
  LAYER VI2 ;
  RECT 2688.260 117.780 2688.460 117.980 ;
  LAYER VI2 ;
  RECT 2687.860 117.780 2688.060 117.980 ;
  LAYER VI3 ;
  RECT 2687.800 114.100 2688.660 114.380 ;
  LAYER VI3 ;
  RECT 2688.260 114.100 2688.460 114.300 ;
  LAYER VI3 ;
  RECT 2687.860 114.100 2688.060 114.300 ;
  LAYER VI2 ;
  RECT 2687.800 114.100 2688.660 114.380 ;
  LAYER VI2 ;
  RECT 2688.260 114.100 2688.460 114.300 ;
  LAYER VI2 ;
  RECT 2687.860 114.100 2688.060 114.300 ;
  LAYER VI3 ;
  RECT 2687.800 110.420 2688.660 110.700 ;
  LAYER VI3 ;
  RECT 2688.260 110.420 2688.460 110.620 ;
  LAYER VI3 ;
  RECT 2687.860 110.420 2688.060 110.620 ;
  LAYER VI2 ;
  RECT 2687.800 110.420 2688.660 110.700 ;
  LAYER VI2 ;
  RECT 2688.260 110.420 2688.460 110.620 ;
  LAYER VI2 ;
  RECT 2687.860 110.420 2688.060 110.620 ;
  LAYER VI3 ;
  RECT 2687.800 106.740 2688.660 107.020 ;
  LAYER VI3 ;
  RECT 2688.260 106.740 2688.460 106.940 ;
  LAYER VI3 ;
  RECT 2687.860 106.740 2688.060 106.940 ;
  LAYER VI2 ;
  RECT 2687.800 106.740 2688.660 107.020 ;
  LAYER VI2 ;
  RECT 2688.260 106.740 2688.460 106.940 ;
  LAYER VI2 ;
  RECT 2687.860 106.740 2688.060 106.940 ;
  LAYER VI3 ;
  RECT 2687.800 103.060 2688.660 103.340 ;
  LAYER VI3 ;
  RECT 2688.260 103.060 2688.460 103.260 ;
  LAYER VI3 ;
  RECT 2687.860 103.060 2688.060 103.260 ;
  LAYER VI2 ;
  RECT 2687.800 103.060 2688.660 103.340 ;
  LAYER VI2 ;
  RECT 2688.260 103.060 2688.460 103.260 ;
  LAYER VI2 ;
  RECT 2687.860 103.060 2688.060 103.260 ;
  LAYER VI3 ;
  RECT 2687.800 99.380 2688.660 99.660 ;
  LAYER VI3 ;
  RECT 2688.260 99.380 2688.460 99.580 ;
  LAYER VI3 ;
  RECT 2687.860 99.380 2688.060 99.580 ;
  LAYER VI2 ;
  RECT 2687.800 99.380 2688.660 99.660 ;
  LAYER VI2 ;
  RECT 2688.260 99.380 2688.460 99.580 ;
  LAYER VI2 ;
  RECT 2687.860 99.380 2688.060 99.580 ;
  LAYER VI3 ;
  RECT 2687.800 95.700 2688.660 95.980 ;
  LAYER VI3 ;
  RECT 2688.260 95.700 2688.460 95.900 ;
  LAYER VI3 ;
  RECT 2687.860 95.700 2688.060 95.900 ;
  LAYER VI2 ;
  RECT 2687.800 95.700 2688.660 95.980 ;
  LAYER VI2 ;
  RECT 2688.260 95.700 2688.460 95.900 ;
  LAYER VI2 ;
  RECT 2687.860 95.700 2688.060 95.900 ;
  LAYER VI3 ;
  RECT 2687.800 92.020 2688.660 92.300 ;
  LAYER VI3 ;
  RECT 2688.260 92.020 2688.460 92.220 ;
  LAYER VI3 ;
  RECT 2687.860 92.020 2688.060 92.220 ;
  LAYER VI2 ;
  RECT 2687.800 92.020 2688.660 92.300 ;
  LAYER VI2 ;
  RECT 2688.260 92.020 2688.460 92.220 ;
  LAYER VI2 ;
  RECT 2687.860 92.020 2688.060 92.220 ;
  LAYER VI3 ;
  RECT 2687.800 88.340 2688.660 88.620 ;
  LAYER VI3 ;
  RECT 2688.260 88.340 2688.460 88.540 ;
  LAYER VI3 ;
  RECT 2687.860 88.340 2688.060 88.540 ;
  LAYER VI2 ;
  RECT 2687.800 88.340 2688.660 88.620 ;
  LAYER VI2 ;
  RECT 2688.260 88.340 2688.460 88.540 ;
  LAYER VI2 ;
  RECT 2687.860 88.340 2688.060 88.540 ;
  LAYER VI3 ;
  RECT 2687.800 84.660 2688.660 84.940 ;
  LAYER VI3 ;
  RECT 2688.260 84.660 2688.460 84.860 ;
  LAYER VI3 ;
  RECT 2687.860 84.660 2688.060 84.860 ;
  LAYER VI2 ;
  RECT 2687.800 84.660 2688.660 84.940 ;
  LAYER VI2 ;
  RECT 2688.260 84.660 2688.460 84.860 ;
  LAYER VI2 ;
  RECT 2687.860 84.660 2688.060 84.860 ;
  LAYER VI3 ;
  RECT 2687.800 80.980 2688.660 81.260 ;
  LAYER VI3 ;
  RECT 2688.260 80.980 2688.460 81.180 ;
  LAYER VI3 ;
  RECT 2687.860 80.980 2688.060 81.180 ;
  LAYER VI2 ;
  RECT 2687.800 80.980 2688.660 81.260 ;
  LAYER VI2 ;
  RECT 2688.260 80.980 2688.460 81.180 ;
  LAYER VI2 ;
  RECT 2687.860 80.980 2688.060 81.180 ;
  LAYER VI3 ;
  RECT 2687.800 77.300 2688.660 77.580 ;
  LAYER VI3 ;
  RECT 2688.260 77.300 2688.460 77.500 ;
  LAYER VI3 ;
  RECT 2687.860 77.300 2688.060 77.500 ;
  LAYER VI2 ;
  RECT 2687.800 77.300 2688.660 77.580 ;
  LAYER VI2 ;
  RECT 2688.260 77.300 2688.460 77.500 ;
  LAYER VI2 ;
  RECT 2687.860 77.300 2688.060 77.500 ;
  LAYER VI3 ;
  RECT 2687.800 73.620 2688.660 73.900 ;
  LAYER VI3 ;
  RECT 2688.260 73.620 2688.460 73.820 ;
  LAYER VI3 ;
  RECT 2687.860 73.620 2688.060 73.820 ;
  LAYER VI2 ;
  RECT 2687.800 73.620 2688.660 73.900 ;
  LAYER VI2 ;
  RECT 2688.260 73.620 2688.460 73.820 ;
  LAYER VI2 ;
  RECT 2687.860 73.620 2688.060 73.820 ;
  LAYER VI3 ;
  RECT 2687.800 69.940 2688.660 70.220 ;
  LAYER VI3 ;
  RECT 2688.260 69.940 2688.460 70.140 ;
  LAYER VI3 ;
  RECT 2687.860 69.940 2688.060 70.140 ;
  LAYER VI2 ;
  RECT 2687.800 69.940 2688.660 70.220 ;
  LAYER VI2 ;
  RECT 2688.260 69.940 2688.460 70.140 ;
  LAYER VI2 ;
  RECT 2687.860 69.940 2688.060 70.140 ;
  LAYER VI3 ;
  RECT 2687.800 65.600 2688.660 65.980 ;
  LAYER VI3 ;
  RECT 2688.200 65.660 2688.400 65.860 ;
  LAYER VI3 ;
  RECT 2687.800 65.660 2688.000 65.860 ;
  LAYER VI2 ;
  RECT 2687.800 65.600 2688.660 65.980 ;
  LAYER VI2 ;
  RECT 2688.200 65.660 2688.400 65.860 ;
  LAYER VI2 ;
  RECT 2687.800 65.660 2688.000 65.860 ;
  LAYER VI3 ;
  RECT 1376.820 560.790 1377.070 561.650 ;
  LAYER VI3 ;
  RECT 1376.820 561.250 1377.020 561.450 ;
  LAYER VI3 ;
  RECT 1376.820 560.850 1377.020 561.050 ;
  LAYER VI2 ;
  RECT 1376.820 560.790 1377.070 561.650 ;
  LAYER VI2 ;
  RECT 1376.820 561.250 1377.020 561.450 ;
  LAYER VI2 ;
  RECT 1376.820 560.850 1377.020 561.050 ;
  LAYER VI3 ;
  RECT 1417.740 560.790 1417.990 561.650 ;
  LAYER VI3 ;
  RECT 1417.740 561.250 1417.940 561.450 ;
  LAYER VI3 ;
  RECT 1417.740 560.850 1417.940 561.050 ;
  LAYER VI2 ;
  RECT 1417.740 560.790 1417.990 561.650 ;
  LAYER VI2 ;
  RECT 1417.740 561.250 1417.940 561.450 ;
  LAYER VI2 ;
  RECT 1417.740 560.850 1417.940 561.050 ;
  LAYER VI3 ;
  RECT 1458.660 560.790 1458.910 561.650 ;
  LAYER VI3 ;
  RECT 1458.660 561.250 1458.860 561.450 ;
  LAYER VI3 ;
  RECT 1458.660 560.850 1458.860 561.050 ;
  LAYER VI2 ;
  RECT 1458.660 560.790 1458.910 561.650 ;
  LAYER VI2 ;
  RECT 1458.660 561.250 1458.860 561.450 ;
  LAYER VI2 ;
  RECT 1458.660 560.850 1458.860 561.050 ;
  LAYER VI3 ;
  RECT 1499.580 560.790 1499.830 561.650 ;
  LAYER VI3 ;
  RECT 1499.580 561.250 1499.780 561.450 ;
  LAYER VI3 ;
  RECT 1499.580 560.850 1499.780 561.050 ;
  LAYER VI2 ;
  RECT 1499.580 560.790 1499.830 561.650 ;
  LAYER VI2 ;
  RECT 1499.580 561.250 1499.780 561.450 ;
  LAYER VI2 ;
  RECT 1499.580 560.850 1499.780 561.050 ;
  LAYER VI3 ;
  RECT 1540.500 560.790 1540.750 561.650 ;
  LAYER VI3 ;
  RECT 1540.500 561.250 1540.700 561.450 ;
  LAYER VI3 ;
  RECT 1540.500 560.850 1540.700 561.050 ;
  LAYER VI2 ;
  RECT 1540.500 560.790 1540.750 561.650 ;
  LAYER VI2 ;
  RECT 1540.500 561.250 1540.700 561.450 ;
  LAYER VI2 ;
  RECT 1540.500 560.850 1540.700 561.050 ;
  LAYER VI3 ;
  RECT 1581.420 560.790 1581.670 561.650 ;
  LAYER VI3 ;
  RECT 1581.420 561.250 1581.620 561.450 ;
  LAYER VI3 ;
  RECT 1581.420 560.850 1581.620 561.050 ;
  LAYER VI2 ;
  RECT 1581.420 560.790 1581.670 561.650 ;
  LAYER VI2 ;
  RECT 1581.420 561.250 1581.620 561.450 ;
  LAYER VI2 ;
  RECT 1581.420 560.850 1581.620 561.050 ;
  LAYER VI3 ;
  RECT 1622.340 560.790 1622.590 561.650 ;
  LAYER VI3 ;
  RECT 1622.340 561.250 1622.540 561.450 ;
  LAYER VI3 ;
  RECT 1622.340 560.850 1622.540 561.050 ;
  LAYER VI2 ;
  RECT 1622.340 560.790 1622.590 561.650 ;
  LAYER VI2 ;
  RECT 1622.340 561.250 1622.540 561.450 ;
  LAYER VI2 ;
  RECT 1622.340 560.850 1622.540 561.050 ;
  LAYER VI3 ;
  RECT 1663.260 560.790 1663.510 561.650 ;
  LAYER VI3 ;
  RECT 1663.260 561.250 1663.460 561.450 ;
  LAYER VI3 ;
  RECT 1663.260 560.850 1663.460 561.050 ;
  LAYER VI2 ;
  RECT 1663.260 560.790 1663.510 561.650 ;
  LAYER VI2 ;
  RECT 1663.260 561.250 1663.460 561.450 ;
  LAYER VI2 ;
  RECT 1663.260 560.850 1663.460 561.050 ;
  LAYER VI3 ;
  RECT 1704.180 560.790 1704.430 561.650 ;
  LAYER VI3 ;
  RECT 1704.180 561.250 1704.380 561.450 ;
  LAYER VI3 ;
  RECT 1704.180 560.850 1704.380 561.050 ;
  LAYER VI2 ;
  RECT 1704.180 560.790 1704.430 561.650 ;
  LAYER VI2 ;
  RECT 1704.180 561.250 1704.380 561.450 ;
  LAYER VI2 ;
  RECT 1704.180 560.850 1704.380 561.050 ;
  LAYER VI3 ;
  RECT 1745.100 560.790 1745.350 561.650 ;
  LAYER VI3 ;
  RECT 1745.100 561.250 1745.300 561.450 ;
  LAYER VI3 ;
  RECT 1745.100 560.850 1745.300 561.050 ;
  LAYER VI2 ;
  RECT 1745.100 560.790 1745.350 561.650 ;
  LAYER VI2 ;
  RECT 1745.100 561.250 1745.300 561.450 ;
  LAYER VI2 ;
  RECT 1745.100 560.850 1745.300 561.050 ;
  LAYER VI3 ;
  RECT 1786.020 560.790 1786.270 561.650 ;
  LAYER VI3 ;
  RECT 1786.020 561.250 1786.220 561.450 ;
  LAYER VI3 ;
  RECT 1786.020 560.850 1786.220 561.050 ;
  LAYER VI2 ;
  RECT 1786.020 560.790 1786.270 561.650 ;
  LAYER VI2 ;
  RECT 1786.020 561.250 1786.220 561.450 ;
  LAYER VI2 ;
  RECT 1786.020 560.850 1786.220 561.050 ;
  LAYER VI3 ;
  RECT 1826.940 560.790 1827.190 561.650 ;
  LAYER VI3 ;
  RECT 1826.940 561.250 1827.140 561.450 ;
  LAYER VI3 ;
  RECT 1826.940 560.850 1827.140 561.050 ;
  LAYER VI2 ;
  RECT 1826.940 560.790 1827.190 561.650 ;
  LAYER VI2 ;
  RECT 1826.940 561.250 1827.140 561.450 ;
  LAYER VI2 ;
  RECT 1826.940 560.850 1827.140 561.050 ;
  LAYER VI3 ;
  RECT 1867.860 560.790 1868.110 561.650 ;
  LAYER VI3 ;
  RECT 1867.860 561.250 1868.060 561.450 ;
  LAYER VI3 ;
  RECT 1867.860 560.850 1868.060 561.050 ;
  LAYER VI2 ;
  RECT 1867.860 560.790 1868.110 561.650 ;
  LAYER VI2 ;
  RECT 1867.860 561.250 1868.060 561.450 ;
  LAYER VI2 ;
  RECT 1867.860 560.850 1868.060 561.050 ;
  LAYER VI3 ;
  RECT 1908.780 560.790 1909.030 561.650 ;
  LAYER VI3 ;
  RECT 1908.780 561.250 1908.980 561.450 ;
  LAYER VI3 ;
  RECT 1908.780 560.850 1908.980 561.050 ;
  LAYER VI2 ;
  RECT 1908.780 560.790 1909.030 561.650 ;
  LAYER VI2 ;
  RECT 1908.780 561.250 1908.980 561.450 ;
  LAYER VI2 ;
  RECT 1908.780 560.850 1908.980 561.050 ;
  LAYER VI3 ;
  RECT 1949.700 560.790 1949.950 561.650 ;
  LAYER VI3 ;
  RECT 1949.700 561.250 1949.900 561.450 ;
  LAYER VI3 ;
  RECT 1949.700 560.850 1949.900 561.050 ;
  LAYER VI2 ;
  RECT 1949.700 560.790 1949.950 561.650 ;
  LAYER VI2 ;
  RECT 1949.700 561.250 1949.900 561.450 ;
  LAYER VI2 ;
  RECT 1949.700 560.850 1949.900 561.050 ;
  LAYER VI3 ;
  RECT 1990.620 560.790 1990.870 561.650 ;
  LAYER VI3 ;
  RECT 1990.620 561.250 1990.820 561.450 ;
  LAYER VI3 ;
  RECT 1990.620 560.850 1990.820 561.050 ;
  LAYER VI2 ;
  RECT 1990.620 560.790 1990.870 561.650 ;
  LAYER VI2 ;
  RECT 1990.620 561.250 1990.820 561.450 ;
  LAYER VI2 ;
  RECT 1990.620 560.850 1990.820 561.050 ;
  LAYER VI3 ;
  RECT 2031.540 560.790 2031.790 561.650 ;
  LAYER VI3 ;
  RECT 2031.540 561.250 2031.740 561.450 ;
  LAYER VI3 ;
  RECT 2031.540 560.850 2031.740 561.050 ;
  LAYER VI2 ;
  RECT 2031.540 560.790 2031.790 561.650 ;
  LAYER VI2 ;
  RECT 2031.540 561.250 2031.740 561.450 ;
  LAYER VI2 ;
  RECT 2031.540 560.850 2031.740 561.050 ;
  LAYER VI3 ;
  RECT 2072.460 560.790 2072.710 561.650 ;
  LAYER VI3 ;
  RECT 2072.460 561.250 2072.660 561.450 ;
  LAYER VI3 ;
  RECT 2072.460 560.850 2072.660 561.050 ;
  LAYER VI2 ;
  RECT 2072.460 560.790 2072.710 561.650 ;
  LAYER VI2 ;
  RECT 2072.460 561.250 2072.660 561.450 ;
  LAYER VI2 ;
  RECT 2072.460 560.850 2072.660 561.050 ;
  LAYER VI3 ;
  RECT 2113.380 560.790 2113.630 561.650 ;
  LAYER VI3 ;
  RECT 2113.380 561.250 2113.580 561.450 ;
  LAYER VI3 ;
  RECT 2113.380 560.850 2113.580 561.050 ;
  LAYER VI2 ;
  RECT 2113.380 560.790 2113.630 561.650 ;
  LAYER VI2 ;
  RECT 2113.380 561.250 2113.580 561.450 ;
  LAYER VI2 ;
  RECT 2113.380 560.850 2113.580 561.050 ;
  LAYER VI3 ;
  RECT 2154.300 560.790 2154.550 561.650 ;
  LAYER VI3 ;
  RECT 2154.300 561.250 2154.500 561.450 ;
  LAYER VI3 ;
  RECT 2154.300 560.850 2154.500 561.050 ;
  LAYER VI2 ;
  RECT 2154.300 560.790 2154.550 561.650 ;
  LAYER VI2 ;
  RECT 2154.300 561.250 2154.500 561.450 ;
  LAYER VI2 ;
  RECT 2154.300 560.850 2154.500 561.050 ;
  LAYER VI3 ;
  RECT 2195.220 560.790 2195.470 561.650 ;
  LAYER VI3 ;
  RECT 2195.220 561.250 2195.420 561.450 ;
  LAYER VI3 ;
  RECT 2195.220 560.850 2195.420 561.050 ;
  LAYER VI2 ;
  RECT 2195.220 560.790 2195.470 561.650 ;
  LAYER VI2 ;
  RECT 2195.220 561.250 2195.420 561.450 ;
  LAYER VI2 ;
  RECT 2195.220 560.850 2195.420 561.050 ;
  LAYER VI3 ;
  RECT 2236.140 560.790 2236.390 561.650 ;
  LAYER VI3 ;
  RECT 2236.140 561.250 2236.340 561.450 ;
  LAYER VI3 ;
  RECT 2236.140 560.850 2236.340 561.050 ;
  LAYER VI2 ;
  RECT 2236.140 560.790 2236.390 561.650 ;
  LAYER VI2 ;
  RECT 2236.140 561.250 2236.340 561.450 ;
  LAYER VI2 ;
  RECT 2236.140 560.850 2236.340 561.050 ;
  LAYER VI3 ;
  RECT 2277.060 560.790 2277.310 561.650 ;
  LAYER VI3 ;
  RECT 2277.060 561.250 2277.260 561.450 ;
  LAYER VI3 ;
  RECT 2277.060 560.850 2277.260 561.050 ;
  LAYER VI2 ;
  RECT 2277.060 560.790 2277.310 561.650 ;
  LAYER VI2 ;
  RECT 2277.060 561.250 2277.260 561.450 ;
  LAYER VI2 ;
  RECT 2277.060 560.850 2277.260 561.050 ;
  LAYER VI3 ;
  RECT 2317.980 560.790 2318.230 561.650 ;
  LAYER VI3 ;
  RECT 2317.980 561.250 2318.180 561.450 ;
  LAYER VI3 ;
  RECT 2317.980 560.850 2318.180 561.050 ;
  LAYER VI2 ;
  RECT 2317.980 560.790 2318.230 561.650 ;
  LAYER VI2 ;
  RECT 2317.980 561.250 2318.180 561.450 ;
  LAYER VI2 ;
  RECT 2317.980 560.850 2318.180 561.050 ;
  LAYER VI3 ;
  RECT 2358.900 560.790 2359.150 561.650 ;
  LAYER VI3 ;
  RECT 2358.900 561.250 2359.100 561.450 ;
  LAYER VI3 ;
  RECT 2358.900 560.850 2359.100 561.050 ;
  LAYER VI2 ;
  RECT 2358.900 560.790 2359.150 561.650 ;
  LAYER VI2 ;
  RECT 2358.900 561.250 2359.100 561.450 ;
  LAYER VI2 ;
  RECT 2358.900 560.850 2359.100 561.050 ;
  LAYER VI3 ;
  RECT 2399.820 560.790 2400.070 561.650 ;
  LAYER VI3 ;
  RECT 2399.820 561.250 2400.020 561.450 ;
  LAYER VI3 ;
  RECT 2399.820 560.850 2400.020 561.050 ;
  LAYER VI2 ;
  RECT 2399.820 560.790 2400.070 561.650 ;
  LAYER VI2 ;
  RECT 2399.820 561.250 2400.020 561.450 ;
  LAYER VI2 ;
  RECT 2399.820 560.850 2400.020 561.050 ;
  LAYER VI3 ;
  RECT 2440.740 560.790 2440.990 561.650 ;
  LAYER VI3 ;
  RECT 2440.740 561.250 2440.940 561.450 ;
  LAYER VI3 ;
  RECT 2440.740 560.850 2440.940 561.050 ;
  LAYER VI2 ;
  RECT 2440.740 560.790 2440.990 561.650 ;
  LAYER VI2 ;
  RECT 2440.740 561.250 2440.940 561.450 ;
  LAYER VI2 ;
  RECT 2440.740 560.850 2440.940 561.050 ;
  LAYER VI3 ;
  RECT 2481.660 560.790 2481.910 561.650 ;
  LAYER VI3 ;
  RECT 2481.660 561.250 2481.860 561.450 ;
  LAYER VI3 ;
  RECT 2481.660 560.850 2481.860 561.050 ;
  LAYER VI2 ;
  RECT 2481.660 560.790 2481.910 561.650 ;
  LAYER VI2 ;
  RECT 2481.660 561.250 2481.860 561.450 ;
  LAYER VI2 ;
  RECT 2481.660 560.850 2481.860 561.050 ;
  LAYER VI3 ;
  RECT 2522.580 560.790 2522.830 561.650 ;
  LAYER VI3 ;
  RECT 2522.580 561.250 2522.780 561.450 ;
  LAYER VI3 ;
  RECT 2522.580 560.850 2522.780 561.050 ;
  LAYER VI2 ;
  RECT 2522.580 560.790 2522.830 561.650 ;
  LAYER VI2 ;
  RECT 2522.580 561.250 2522.780 561.450 ;
  LAYER VI2 ;
  RECT 2522.580 560.850 2522.780 561.050 ;
  LAYER VI3 ;
  RECT 2563.500 560.790 2563.750 561.650 ;
  LAYER VI3 ;
  RECT 2563.500 561.250 2563.700 561.450 ;
  LAYER VI3 ;
  RECT 2563.500 560.850 2563.700 561.050 ;
  LAYER VI2 ;
  RECT 2563.500 560.790 2563.750 561.650 ;
  LAYER VI2 ;
  RECT 2563.500 561.250 2563.700 561.450 ;
  LAYER VI2 ;
  RECT 2563.500 560.850 2563.700 561.050 ;
  LAYER VI3 ;
  RECT 2604.420 560.790 2604.670 561.650 ;
  LAYER VI3 ;
  RECT 2604.420 561.250 2604.620 561.450 ;
  LAYER VI3 ;
  RECT 2604.420 560.850 2604.620 561.050 ;
  LAYER VI2 ;
  RECT 2604.420 560.790 2604.670 561.650 ;
  LAYER VI2 ;
  RECT 2604.420 561.250 2604.620 561.450 ;
  LAYER VI2 ;
  RECT 2604.420 560.850 2604.620 561.050 ;
  LAYER VI3 ;
  RECT 2645.340 560.790 2645.590 561.650 ;
  LAYER VI3 ;
  RECT 2645.340 561.250 2645.540 561.450 ;
  LAYER VI3 ;
  RECT 2645.340 560.850 2645.540 561.050 ;
  LAYER VI2 ;
  RECT 2645.340 560.790 2645.590 561.650 ;
  LAYER VI2 ;
  RECT 2645.340 561.250 2645.540 561.450 ;
  LAYER VI2 ;
  RECT 2645.340 560.850 2645.540 561.050 ;
  LAYER VI3 ;
  RECT 1359.810 560.790 1362.320 561.650 ;
  LAYER VI3 ;
  RECT 1361.810 561.250 1362.010 561.450 ;
  LAYER VI3 ;
  RECT 1361.810 560.850 1362.010 561.050 ;
  LAYER VI3 ;
  RECT 1361.410 561.250 1361.610 561.450 ;
  LAYER VI3 ;
  RECT 1361.410 560.850 1361.610 561.050 ;
  LAYER VI3 ;
  RECT 1361.010 561.250 1361.210 561.450 ;
  LAYER VI3 ;
  RECT 1361.010 560.850 1361.210 561.050 ;
  LAYER VI3 ;
  RECT 1360.610 561.250 1360.810 561.450 ;
  LAYER VI3 ;
  RECT 1360.610 560.850 1360.810 561.050 ;
  LAYER VI3 ;
  RECT 1360.210 561.250 1360.410 561.450 ;
  LAYER VI3 ;
  RECT 1360.210 560.850 1360.410 561.050 ;
  LAYER VI3 ;
  RECT 1359.810 561.250 1360.010 561.450 ;
  LAYER VI3 ;
  RECT 1359.810 560.850 1360.010 561.050 ;
  LAYER VI2 ;
  RECT 1359.810 560.790 1362.320 561.650 ;
  LAYER VI2 ;
  RECT 1361.810 561.250 1362.010 561.450 ;
  LAYER VI2 ;
  RECT 1361.810 560.850 1362.010 561.050 ;
  LAYER VI2 ;
  RECT 1361.410 561.250 1361.610 561.450 ;
  LAYER VI2 ;
  RECT 1361.410 560.850 1361.610 561.050 ;
  LAYER VI2 ;
  RECT 1361.010 561.250 1361.210 561.450 ;
  LAYER VI2 ;
  RECT 1361.010 560.850 1361.210 561.050 ;
  LAYER VI2 ;
  RECT 1360.610 561.250 1360.810 561.450 ;
  LAYER VI2 ;
  RECT 1360.610 560.850 1360.810 561.050 ;
  LAYER VI2 ;
  RECT 1360.210 561.250 1360.410 561.450 ;
  LAYER VI2 ;
  RECT 1360.210 560.850 1360.410 561.050 ;
  LAYER VI2 ;
  RECT 1359.810 561.250 1360.010 561.450 ;
  LAYER VI2 ;
  RECT 1359.810 560.850 1360.010 561.050 ;
  LAYER VI3 ;
  RECT 1347.390 560.790 1349.780 561.650 ;
  LAYER VI3 ;
  RECT 1349.390 561.250 1349.590 561.450 ;
  LAYER VI3 ;
  RECT 1349.390 560.850 1349.590 561.050 ;
  LAYER VI3 ;
  RECT 1348.990 561.250 1349.190 561.450 ;
  LAYER VI3 ;
  RECT 1348.990 560.850 1349.190 561.050 ;
  LAYER VI3 ;
  RECT 1348.590 561.250 1348.790 561.450 ;
  LAYER VI3 ;
  RECT 1348.590 560.850 1348.790 561.050 ;
  LAYER VI3 ;
  RECT 1348.190 561.250 1348.390 561.450 ;
  LAYER VI3 ;
  RECT 1348.190 560.850 1348.390 561.050 ;
  LAYER VI3 ;
  RECT 1347.790 561.250 1347.990 561.450 ;
  LAYER VI3 ;
  RECT 1347.790 560.850 1347.990 561.050 ;
  LAYER VI3 ;
  RECT 1347.390 561.250 1347.590 561.450 ;
  LAYER VI3 ;
  RECT 1347.390 560.850 1347.590 561.050 ;
  LAYER VI2 ;
  RECT 1347.390 560.790 1349.780 561.650 ;
  LAYER VI2 ;
  RECT 1349.390 561.250 1349.590 561.450 ;
  LAYER VI2 ;
  RECT 1349.390 560.850 1349.590 561.050 ;
  LAYER VI2 ;
  RECT 1348.990 561.250 1349.190 561.450 ;
  LAYER VI2 ;
  RECT 1348.990 560.850 1349.190 561.050 ;
  LAYER VI2 ;
  RECT 1348.590 561.250 1348.790 561.450 ;
  LAYER VI2 ;
  RECT 1348.590 560.850 1348.790 561.050 ;
  LAYER VI2 ;
  RECT 1348.190 561.250 1348.390 561.450 ;
  LAYER VI2 ;
  RECT 1348.190 560.850 1348.390 561.050 ;
  LAYER VI2 ;
  RECT 1347.790 561.250 1347.990 561.450 ;
  LAYER VI2 ;
  RECT 1347.790 560.850 1347.990 561.050 ;
  LAYER VI2 ;
  RECT 1347.390 561.250 1347.590 561.450 ;
  LAYER VI2 ;
  RECT 1347.390 560.850 1347.590 561.050 ;
  LAYER VI3 ;
  RECT 1339.880 560.790 1342.940 561.650 ;
  LAYER VI3 ;
  RECT 1342.680 561.250 1342.880 561.450 ;
  LAYER VI3 ;
  RECT 1342.680 560.850 1342.880 561.050 ;
  LAYER VI3 ;
  RECT 1342.280 561.250 1342.480 561.450 ;
  LAYER VI3 ;
  RECT 1342.280 560.850 1342.480 561.050 ;
  LAYER VI3 ;
  RECT 1341.880 561.250 1342.080 561.450 ;
  LAYER VI3 ;
  RECT 1341.880 560.850 1342.080 561.050 ;
  LAYER VI3 ;
  RECT 1341.480 561.250 1341.680 561.450 ;
  LAYER VI3 ;
  RECT 1341.480 560.850 1341.680 561.050 ;
  LAYER VI3 ;
  RECT 1341.080 561.250 1341.280 561.450 ;
  LAYER VI3 ;
  RECT 1341.080 560.850 1341.280 561.050 ;
  LAYER VI3 ;
  RECT 1340.680 561.250 1340.880 561.450 ;
  LAYER VI3 ;
  RECT 1340.680 560.850 1340.880 561.050 ;
  LAYER VI3 ;
  RECT 1340.280 561.250 1340.480 561.450 ;
  LAYER VI3 ;
  RECT 1340.280 560.850 1340.480 561.050 ;
  LAYER VI3 ;
  RECT 1339.880 561.250 1340.080 561.450 ;
  LAYER VI3 ;
  RECT 1339.880 560.850 1340.080 561.050 ;
  LAYER VI2 ;
  RECT 1339.880 560.790 1342.940 561.650 ;
  LAYER VI2 ;
  RECT 1342.680 561.250 1342.880 561.450 ;
  LAYER VI2 ;
  RECT 1342.680 560.850 1342.880 561.050 ;
  LAYER VI2 ;
  RECT 1342.280 561.250 1342.480 561.450 ;
  LAYER VI2 ;
  RECT 1342.280 560.850 1342.480 561.050 ;
  LAYER VI2 ;
  RECT 1341.880 561.250 1342.080 561.450 ;
  LAYER VI2 ;
  RECT 1341.880 560.850 1342.080 561.050 ;
  LAYER VI2 ;
  RECT 1341.480 561.250 1341.680 561.450 ;
  LAYER VI2 ;
  RECT 1341.480 560.850 1341.680 561.050 ;
  LAYER VI2 ;
  RECT 1341.080 561.250 1341.280 561.450 ;
  LAYER VI2 ;
  RECT 1341.080 560.850 1341.280 561.050 ;
  LAYER VI2 ;
  RECT 1340.680 561.250 1340.880 561.450 ;
  LAYER VI2 ;
  RECT 1340.680 560.850 1340.880 561.050 ;
  LAYER VI2 ;
  RECT 1340.280 561.250 1340.480 561.450 ;
  LAYER VI2 ;
  RECT 1340.280 560.850 1340.480 561.050 ;
  LAYER VI2 ;
  RECT 1339.880 561.250 1340.080 561.450 ;
  LAYER VI2 ;
  RECT 1339.880 560.850 1340.080 561.050 ;
  LAYER VI3 ;
  RECT 1364.060 560.790 1366.910 561.650 ;
  LAYER VI3 ;
  RECT 1366.460 561.250 1366.660 561.450 ;
  LAYER VI3 ;
  RECT 1366.460 560.850 1366.660 561.050 ;
  LAYER VI3 ;
  RECT 1366.060 561.250 1366.260 561.450 ;
  LAYER VI3 ;
  RECT 1366.060 560.850 1366.260 561.050 ;
  LAYER VI3 ;
  RECT 1365.660 561.250 1365.860 561.450 ;
  LAYER VI3 ;
  RECT 1365.660 560.850 1365.860 561.050 ;
  LAYER VI3 ;
  RECT 1365.260 561.250 1365.460 561.450 ;
  LAYER VI3 ;
  RECT 1365.260 560.850 1365.460 561.050 ;
  LAYER VI3 ;
  RECT 1364.860 561.250 1365.060 561.450 ;
  LAYER VI3 ;
  RECT 1364.860 560.850 1365.060 561.050 ;
  LAYER VI3 ;
  RECT 1364.460 561.250 1364.660 561.450 ;
  LAYER VI3 ;
  RECT 1364.460 560.850 1364.660 561.050 ;
  LAYER VI3 ;
  RECT 1364.060 561.250 1364.260 561.450 ;
  LAYER VI3 ;
  RECT 1364.060 560.850 1364.260 561.050 ;
  LAYER VI2 ;
  RECT 1364.060 560.790 1366.910 561.650 ;
  LAYER VI2 ;
  RECT 1366.460 561.250 1366.660 561.450 ;
  LAYER VI2 ;
  RECT 1366.460 560.850 1366.660 561.050 ;
  LAYER VI2 ;
  RECT 1366.060 561.250 1366.260 561.450 ;
  LAYER VI2 ;
  RECT 1366.060 560.850 1366.260 561.050 ;
  LAYER VI2 ;
  RECT 1365.660 561.250 1365.860 561.450 ;
  LAYER VI2 ;
  RECT 1365.660 560.850 1365.860 561.050 ;
  LAYER VI2 ;
  RECT 1365.260 561.250 1365.460 561.450 ;
  LAYER VI2 ;
  RECT 1365.260 560.850 1365.460 561.050 ;
  LAYER VI2 ;
  RECT 1364.860 561.250 1365.060 561.450 ;
  LAYER VI2 ;
  RECT 1364.860 560.850 1365.060 561.050 ;
  LAYER VI2 ;
  RECT 1364.460 561.250 1364.660 561.450 ;
  LAYER VI2 ;
  RECT 1364.460 560.850 1364.660 561.050 ;
  LAYER VI2 ;
  RECT 1364.060 561.250 1364.260 561.450 ;
  LAYER VI2 ;
  RECT 1364.060 560.850 1364.260 561.050 ;
  LAYER VI3 ;
  RECT 1368.360 560.790 1371.610 561.650 ;
  LAYER VI3 ;
  RECT 1371.160 561.250 1371.360 561.450 ;
  LAYER VI3 ;
  RECT 1371.160 560.850 1371.360 561.050 ;
  LAYER VI3 ;
  RECT 1370.760 561.250 1370.960 561.450 ;
  LAYER VI3 ;
  RECT 1370.760 560.850 1370.960 561.050 ;
  LAYER VI3 ;
  RECT 1370.360 561.250 1370.560 561.450 ;
  LAYER VI3 ;
  RECT 1370.360 560.850 1370.560 561.050 ;
  LAYER VI3 ;
  RECT 1369.960 561.250 1370.160 561.450 ;
  LAYER VI3 ;
  RECT 1369.960 560.850 1370.160 561.050 ;
  LAYER VI3 ;
  RECT 1369.560 561.250 1369.760 561.450 ;
  LAYER VI3 ;
  RECT 1369.560 560.850 1369.760 561.050 ;
  LAYER VI3 ;
  RECT 1369.160 561.250 1369.360 561.450 ;
  LAYER VI3 ;
  RECT 1369.160 560.850 1369.360 561.050 ;
  LAYER VI3 ;
  RECT 1368.760 561.250 1368.960 561.450 ;
  LAYER VI3 ;
  RECT 1368.760 560.850 1368.960 561.050 ;
  LAYER VI3 ;
  RECT 1368.360 561.250 1368.560 561.450 ;
  LAYER VI3 ;
  RECT 1368.360 560.850 1368.560 561.050 ;
  LAYER VI2 ;
  RECT 1368.360 560.790 1371.610 561.650 ;
  LAYER VI2 ;
  RECT 1371.160 561.250 1371.360 561.450 ;
  LAYER VI2 ;
  RECT 1371.160 560.850 1371.360 561.050 ;
  LAYER VI2 ;
  RECT 1370.760 561.250 1370.960 561.450 ;
  LAYER VI2 ;
  RECT 1370.760 560.850 1370.960 561.050 ;
  LAYER VI2 ;
  RECT 1370.360 561.250 1370.560 561.450 ;
  LAYER VI2 ;
  RECT 1370.360 560.850 1370.560 561.050 ;
  LAYER VI2 ;
  RECT 1369.960 561.250 1370.160 561.450 ;
  LAYER VI2 ;
  RECT 1369.960 560.850 1370.160 561.050 ;
  LAYER VI2 ;
  RECT 1369.560 561.250 1369.760 561.450 ;
  LAYER VI2 ;
  RECT 1369.560 560.850 1369.760 561.050 ;
  LAYER VI2 ;
  RECT 1369.160 561.250 1369.360 561.450 ;
  LAYER VI2 ;
  RECT 1369.160 560.850 1369.360 561.050 ;
  LAYER VI2 ;
  RECT 1368.760 561.250 1368.960 561.450 ;
  LAYER VI2 ;
  RECT 1368.760 560.850 1368.960 561.050 ;
  LAYER VI2 ;
  RECT 1368.360 561.250 1368.560 561.450 ;
  LAYER VI2 ;
  RECT 1368.360 560.850 1368.560 561.050 ;
  LAYER VI3 ;
  RECT 1337.160 560.790 1338.920 561.650 ;
  LAYER VI3 ;
  RECT 1338.360 561.250 1338.560 561.450 ;
  LAYER VI3 ;
  RECT 1338.360 560.850 1338.560 561.050 ;
  LAYER VI3 ;
  RECT 1337.960 561.250 1338.160 561.450 ;
  LAYER VI3 ;
  RECT 1337.960 560.850 1338.160 561.050 ;
  LAYER VI3 ;
  RECT 1337.560 561.250 1337.760 561.450 ;
  LAYER VI3 ;
  RECT 1337.560 560.850 1337.760 561.050 ;
  LAYER VI3 ;
  RECT 1337.160 561.250 1337.360 561.450 ;
  LAYER VI3 ;
  RECT 1337.160 560.850 1337.360 561.050 ;
  LAYER VI2 ;
  RECT 1337.160 560.790 1338.920 561.650 ;
  LAYER VI2 ;
  RECT 1338.360 561.250 1338.560 561.450 ;
  LAYER VI2 ;
  RECT 1338.360 560.850 1338.560 561.050 ;
  LAYER VI2 ;
  RECT 1337.960 561.250 1338.160 561.450 ;
  LAYER VI2 ;
  RECT 1337.960 560.850 1338.160 561.050 ;
  LAYER VI2 ;
  RECT 1337.560 561.250 1337.760 561.450 ;
  LAYER VI2 ;
  RECT 1337.560 560.850 1337.760 561.050 ;
  LAYER VI2 ;
  RECT 1337.160 561.250 1337.360 561.450 ;
  LAYER VI2 ;
  RECT 1337.160 560.850 1337.360 561.050 ;
  LAYER VI3 ;
  RECT 1319.820 560.790 1321.580 561.650 ;
  LAYER VI3 ;
  RECT 1321.020 561.250 1321.220 561.450 ;
  LAYER VI3 ;
  RECT 1321.020 560.850 1321.220 561.050 ;
  LAYER VI3 ;
  RECT 1320.620 561.250 1320.820 561.450 ;
  LAYER VI3 ;
  RECT 1320.620 560.850 1320.820 561.050 ;
  LAYER VI3 ;
  RECT 1320.220 561.250 1320.420 561.450 ;
  LAYER VI3 ;
  RECT 1320.220 560.850 1320.420 561.050 ;
  LAYER VI3 ;
  RECT 1319.820 561.250 1320.020 561.450 ;
  LAYER VI3 ;
  RECT 1319.820 560.850 1320.020 561.050 ;
  LAYER VI2 ;
  RECT 1319.820 560.790 1321.580 561.650 ;
  LAYER VI2 ;
  RECT 1321.020 561.250 1321.220 561.450 ;
  LAYER VI2 ;
  RECT 1321.020 560.850 1321.220 561.050 ;
  LAYER VI2 ;
  RECT 1320.620 561.250 1320.820 561.450 ;
  LAYER VI2 ;
  RECT 1320.620 560.850 1320.820 561.050 ;
  LAYER VI2 ;
  RECT 1320.220 561.250 1320.420 561.450 ;
  LAYER VI2 ;
  RECT 1320.220 560.850 1320.420 561.050 ;
  LAYER VI2 ;
  RECT 1319.820 561.250 1320.020 561.450 ;
  LAYER VI2 ;
  RECT 1319.820 560.850 1320.020 561.050 ;
  LAYER VI3 ;
  RECT 1323.820 560.790 1325.580 561.650 ;
  LAYER VI3 ;
  RECT 1325.020 561.250 1325.220 561.450 ;
  LAYER VI3 ;
  RECT 1325.020 560.850 1325.220 561.050 ;
  LAYER VI3 ;
  RECT 1324.620 561.250 1324.820 561.450 ;
  LAYER VI3 ;
  RECT 1324.620 560.850 1324.820 561.050 ;
  LAYER VI3 ;
  RECT 1324.220 561.250 1324.420 561.450 ;
  LAYER VI3 ;
  RECT 1324.220 560.850 1324.420 561.050 ;
  LAYER VI3 ;
  RECT 1323.820 561.250 1324.020 561.450 ;
  LAYER VI3 ;
  RECT 1323.820 560.850 1324.020 561.050 ;
  LAYER VI2 ;
  RECT 1323.820 560.790 1325.580 561.650 ;
  LAYER VI2 ;
  RECT 1325.020 561.250 1325.220 561.450 ;
  LAYER VI2 ;
  RECT 1325.020 560.850 1325.220 561.050 ;
  LAYER VI2 ;
  RECT 1324.620 561.250 1324.820 561.450 ;
  LAYER VI2 ;
  RECT 1324.620 560.850 1324.820 561.050 ;
  LAYER VI2 ;
  RECT 1324.220 561.250 1324.420 561.450 ;
  LAYER VI2 ;
  RECT 1324.220 560.850 1324.420 561.050 ;
  LAYER VI2 ;
  RECT 1323.820 561.250 1324.020 561.450 ;
  LAYER VI2 ;
  RECT 1323.820 560.850 1324.020 561.050 ;
  LAYER VI3 ;
  RECT 1327.820 560.790 1329.580 561.650 ;
  LAYER VI3 ;
  RECT 1329.020 561.250 1329.220 561.450 ;
  LAYER VI3 ;
  RECT 1329.020 560.850 1329.220 561.050 ;
  LAYER VI3 ;
  RECT 1328.620 561.250 1328.820 561.450 ;
  LAYER VI3 ;
  RECT 1328.620 560.850 1328.820 561.050 ;
  LAYER VI3 ;
  RECT 1328.220 561.250 1328.420 561.450 ;
  LAYER VI3 ;
  RECT 1328.220 560.850 1328.420 561.050 ;
  LAYER VI3 ;
  RECT 1327.820 561.250 1328.020 561.450 ;
  LAYER VI3 ;
  RECT 1327.820 560.850 1328.020 561.050 ;
  LAYER VI2 ;
  RECT 1327.820 560.790 1329.580 561.650 ;
  LAYER VI2 ;
  RECT 1329.020 561.250 1329.220 561.450 ;
  LAYER VI2 ;
  RECT 1329.020 560.850 1329.220 561.050 ;
  LAYER VI2 ;
  RECT 1328.620 561.250 1328.820 561.450 ;
  LAYER VI2 ;
  RECT 1328.620 560.850 1328.820 561.050 ;
  LAYER VI2 ;
  RECT 1328.220 561.250 1328.420 561.450 ;
  LAYER VI2 ;
  RECT 1328.220 560.850 1328.420 561.050 ;
  LAYER VI2 ;
  RECT 1327.820 561.250 1328.020 561.450 ;
  LAYER VI2 ;
  RECT 1327.820 560.850 1328.020 561.050 ;
  LAYER VI3 ;
  RECT 1331.820 560.790 1333.580 561.650 ;
  LAYER VI3 ;
  RECT 1333.020 561.250 1333.220 561.450 ;
  LAYER VI3 ;
  RECT 1333.020 560.850 1333.220 561.050 ;
  LAYER VI3 ;
  RECT 1332.620 561.250 1332.820 561.450 ;
  LAYER VI3 ;
  RECT 1332.620 560.850 1332.820 561.050 ;
  LAYER VI3 ;
  RECT 1332.220 561.250 1332.420 561.450 ;
  LAYER VI3 ;
  RECT 1332.220 560.850 1332.420 561.050 ;
  LAYER VI3 ;
  RECT 1331.820 561.250 1332.020 561.450 ;
  LAYER VI3 ;
  RECT 1331.820 560.850 1332.020 561.050 ;
  LAYER VI2 ;
  RECT 1331.820 560.790 1333.580 561.650 ;
  LAYER VI2 ;
  RECT 1333.020 561.250 1333.220 561.450 ;
  LAYER VI2 ;
  RECT 1333.020 560.850 1333.220 561.050 ;
  LAYER VI2 ;
  RECT 1332.620 561.250 1332.820 561.450 ;
  LAYER VI2 ;
  RECT 1332.620 560.850 1332.820 561.050 ;
  LAYER VI2 ;
  RECT 1332.220 561.250 1332.420 561.450 ;
  LAYER VI2 ;
  RECT 1332.220 560.850 1332.420 561.050 ;
  LAYER VI2 ;
  RECT 1331.820 561.250 1332.020 561.450 ;
  LAYER VI2 ;
  RECT 1331.820 560.850 1332.020 561.050 ;
  LAYER VI3 ;
  RECT 4.280 65.600 5.140 65.980 ;
  LAYER VI3 ;
  RECT 4.680 65.660 4.880 65.860 ;
  LAYER VI3 ;
  RECT 4.280 65.660 4.480 65.860 ;
  LAYER VI2 ;
  RECT 4.280 65.600 5.140 65.980 ;
  LAYER VI2 ;
  RECT 4.680 65.660 4.880 65.860 ;
  LAYER VI2 ;
  RECT 4.280 65.660 4.480 65.860 ;
  LAYER VI3 ;
  RECT 4.280 69.940 5.140 70.220 ;
  LAYER VI3 ;
  RECT 4.740 69.940 4.940 70.140 ;
  LAYER VI3 ;
  RECT 4.340 69.940 4.540 70.140 ;
  LAYER VI2 ;
  RECT 4.280 69.940 5.140 70.220 ;
  LAYER VI2 ;
  RECT 4.740 69.940 4.940 70.140 ;
  LAYER VI2 ;
  RECT 4.340 69.940 4.540 70.140 ;
  LAYER VI3 ;
  RECT 4.280 73.620 5.140 73.900 ;
  LAYER VI3 ;
  RECT 4.740 73.620 4.940 73.820 ;
  LAYER VI3 ;
  RECT 4.340 73.620 4.540 73.820 ;
  LAYER VI2 ;
  RECT 4.280 73.620 5.140 73.900 ;
  LAYER VI2 ;
  RECT 4.740 73.620 4.940 73.820 ;
  LAYER VI2 ;
  RECT 4.340 73.620 4.540 73.820 ;
  LAYER VI3 ;
  RECT 4.280 77.300 5.140 77.580 ;
  LAYER VI3 ;
  RECT 4.740 77.300 4.940 77.500 ;
  LAYER VI3 ;
  RECT 4.340 77.300 4.540 77.500 ;
  LAYER VI2 ;
  RECT 4.280 77.300 5.140 77.580 ;
  LAYER VI2 ;
  RECT 4.740 77.300 4.940 77.500 ;
  LAYER VI2 ;
  RECT 4.340 77.300 4.540 77.500 ;
  LAYER VI3 ;
  RECT 4.280 80.980 5.140 81.260 ;
  LAYER VI3 ;
  RECT 4.740 80.980 4.940 81.180 ;
  LAYER VI3 ;
  RECT 4.340 80.980 4.540 81.180 ;
  LAYER VI2 ;
  RECT 4.280 80.980 5.140 81.260 ;
  LAYER VI2 ;
  RECT 4.740 80.980 4.940 81.180 ;
  LAYER VI2 ;
  RECT 4.340 80.980 4.540 81.180 ;
  LAYER VI3 ;
  RECT 4.280 84.660 5.140 84.940 ;
  LAYER VI3 ;
  RECT 4.740 84.660 4.940 84.860 ;
  LAYER VI3 ;
  RECT 4.340 84.660 4.540 84.860 ;
  LAYER VI2 ;
  RECT 4.280 84.660 5.140 84.940 ;
  LAYER VI2 ;
  RECT 4.740 84.660 4.940 84.860 ;
  LAYER VI2 ;
  RECT 4.340 84.660 4.540 84.860 ;
  LAYER VI3 ;
  RECT 4.280 88.340 5.140 88.620 ;
  LAYER VI3 ;
  RECT 4.740 88.340 4.940 88.540 ;
  LAYER VI3 ;
  RECT 4.340 88.340 4.540 88.540 ;
  LAYER VI2 ;
  RECT 4.280 88.340 5.140 88.620 ;
  LAYER VI2 ;
  RECT 4.740 88.340 4.940 88.540 ;
  LAYER VI2 ;
  RECT 4.340 88.340 4.540 88.540 ;
  LAYER VI3 ;
  RECT 4.280 92.020 5.140 92.300 ;
  LAYER VI3 ;
  RECT 4.740 92.020 4.940 92.220 ;
  LAYER VI3 ;
  RECT 4.340 92.020 4.540 92.220 ;
  LAYER VI2 ;
  RECT 4.280 92.020 5.140 92.300 ;
  LAYER VI2 ;
  RECT 4.740 92.020 4.940 92.220 ;
  LAYER VI2 ;
  RECT 4.340 92.020 4.540 92.220 ;
  LAYER VI3 ;
  RECT 4.280 95.700 5.140 95.980 ;
  LAYER VI3 ;
  RECT 4.740 95.700 4.940 95.900 ;
  LAYER VI3 ;
  RECT 4.340 95.700 4.540 95.900 ;
  LAYER VI2 ;
  RECT 4.280 95.700 5.140 95.980 ;
  LAYER VI2 ;
  RECT 4.740 95.700 4.940 95.900 ;
  LAYER VI2 ;
  RECT 4.340 95.700 4.540 95.900 ;
  LAYER VI3 ;
  RECT 4.280 99.380 5.140 99.660 ;
  LAYER VI3 ;
  RECT 4.740 99.380 4.940 99.580 ;
  LAYER VI3 ;
  RECT 4.340 99.380 4.540 99.580 ;
  LAYER VI2 ;
  RECT 4.280 99.380 5.140 99.660 ;
  LAYER VI2 ;
  RECT 4.740 99.380 4.940 99.580 ;
  LAYER VI2 ;
  RECT 4.340 99.380 4.540 99.580 ;
  LAYER VI3 ;
  RECT 4.280 103.060 5.140 103.340 ;
  LAYER VI3 ;
  RECT 4.740 103.060 4.940 103.260 ;
  LAYER VI3 ;
  RECT 4.340 103.060 4.540 103.260 ;
  LAYER VI2 ;
  RECT 4.280 103.060 5.140 103.340 ;
  LAYER VI2 ;
  RECT 4.740 103.060 4.940 103.260 ;
  LAYER VI2 ;
  RECT 4.340 103.060 4.540 103.260 ;
  LAYER VI3 ;
  RECT 4.280 106.740 5.140 107.020 ;
  LAYER VI3 ;
  RECT 4.740 106.740 4.940 106.940 ;
  LAYER VI3 ;
  RECT 4.340 106.740 4.540 106.940 ;
  LAYER VI2 ;
  RECT 4.280 106.740 5.140 107.020 ;
  LAYER VI2 ;
  RECT 4.740 106.740 4.940 106.940 ;
  LAYER VI2 ;
  RECT 4.340 106.740 4.540 106.940 ;
  LAYER VI3 ;
  RECT 4.280 110.420 5.140 110.700 ;
  LAYER VI3 ;
  RECT 4.740 110.420 4.940 110.620 ;
  LAYER VI3 ;
  RECT 4.340 110.420 4.540 110.620 ;
  LAYER VI2 ;
  RECT 4.280 110.420 5.140 110.700 ;
  LAYER VI2 ;
  RECT 4.740 110.420 4.940 110.620 ;
  LAYER VI2 ;
  RECT 4.340 110.420 4.540 110.620 ;
  LAYER VI3 ;
  RECT 4.280 114.100 5.140 114.380 ;
  LAYER VI3 ;
  RECT 4.740 114.100 4.940 114.300 ;
  LAYER VI3 ;
  RECT 4.340 114.100 4.540 114.300 ;
  LAYER VI2 ;
  RECT 4.280 114.100 5.140 114.380 ;
  LAYER VI2 ;
  RECT 4.740 114.100 4.940 114.300 ;
  LAYER VI2 ;
  RECT 4.340 114.100 4.540 114.300 ;
  LAYER VI3 ;
  RECT 4.280 117.780 5.140 118.060 ;
  LAYER VI3 ;
  RECT 4.740 117.780 4.940 117.980 ;
  LAYER VI3 ;
  RECT 4.340 117.780 4.540 117.980 ;
  LAYER VI2 ;
  RECT 4.280 117.780 5.140 118.060 ;
  LAYER VI2 ;
  RECT 4.740 117.780 4.940 117.980 ;
  LAYER VI2 ;
  RECT 4.340 117.780 4.540 117.980 ;
  LAYER VI3 ;
  RECT 4.280 121.460 5.140 121.740 ;
  LAYER VI3 ;
  RECT 4.740 121.460 4.940 121.660 ;
  LAYER VI3 ;
  RECT 4.340 121.460 4.540 121.660 ;
  LAYER VI2 ;
  RECT 4.280 121.460 5.140 121.740 ;
  LAYER VI2 ;
  RECT 4.740 121.460 4.940 121.660 ;
  LAYER VI2 ;
  RECT 4.340 121.460 4.540 121.660 ;
  LAYER VI3 ;
  RECT 4.280 125.140 5.140 125.420 ;
  LAYER VI3 ;
  RECT 4.740 125.140 4.940 125.340 ;
  LAYER VI3 ;
  RECT 4.340 125.140 4.540 125.340 ;
  LAYER VI2 ;
  RECT 4.280 125.140 5.140 125.420 ;
  LAYER VI2 ;
  RECT 4.740 125.140 4.940 125.340 ;
  LAYER VI2 ;
  RECT 4.340 125.140 4.540 125.340 ;
  LAYER VI3 ;
  RECT 4.280 128.820 5.140 129.100 ;
  LAYER VI3 ;
  RECT 4.740 128.820 4.940 129.020 ;
  LAYER VI3 ;
  RECT 4.340 128.820 4.540 129.020 ;
  LAYER VI2 ;
  RECT 4.280 128.820 5.140 129.100 ;
  LAYER VI2 ;
  RECT 4.740 128.820 4.940 129.020 ;
  LAYER VI2 ;
  RECT 4.340 128.820 4.540 129.020 ;
  LAYER VI3 ;
  RECT 4.280 132.500 5.140 132.780 ;
  LAYER VI3 ;
  RECT 4.740 132.500 4.940 132.700 ;
  LAYER VI3 ;
  RECT 4.340 132.500 4.540 132.700 ;
  LAYER VI2 ;
  RECT 4.280 132.500 5.140 132.780 ;
  LAYER VI2 ;
  RECT 4.740 132.500 4.940 132.700 ;
  LAYER VI2 ;
  RECT 4.340 132.500 4.540 132.700 ;
  LAYER VI3 ;
  RECT 4.280 136.180 5.140 136.460 ;
  LAYER VI3 ;
  RECT 4.740 136.180 4.940 136.380 ;
  LAYER VI3 ;
  RECT 4.340 136.180 4.540 136.380 ;
  LAYER VI2 ;
  RECT 4.280 136.180 5.140 136.460 ;
  LAYER VI2 ;
  RECT 4.740 136.180 4.940 136.380 ;
  LAYER VI2 ;
  RECT 4.340 136.180 4.540 136.380 ;
  LAYER VI3 ;
  RECT 4.280 139.860 5.140 140.140 ;
  LAYER VI3 ;
  RECT 4.740 139.860 4.940 140.060 ;
  LAYER VI3 ;
  RECT 4.340 139.860 4.540 140.060 ;
  LAYER VI2 ;
  RECT 4.280 139.860 5.140 140.140 ;
  LAYER VI2 ;
  RECT 4.740 139.860 4.940 140.060 ;
  LAYER VI2 ;
  RECT 4.340 139.860 4.540 140.060 ;
  LAYER VI3 ;
  RECT 4.280 143.540 5.140 143.820 ;
  LAYER VI3 ;
  RECT 4.740 143.540 4.940 143.740 ;
  LAYER VI3 ;
  RECT 4.340 143.540 4.540 143.740 ;
  LAYER VI2 ;
  RECT 4.280 143.540 5.140 143.820 ;
  LAYER VI2 ;
  RECT 4.740 143.540 4.940 143.740 ;
  LAYER VI2 ;
  RECT 4.340 143.540 4.540 143.740 ;
  LAYER VI3 ;
  RECT 4.280 147.220 5.140 147.500 ;
  LAYER VI3 ;
  RECT 4.740 147.220 4.940 147.420 ;
  LAYER VI3 ;
  RECT 4.340 147.220 4.540 147.420 ;
  LAYER VI2 ;
  RECT 4.280 147.220 5.140 147.500 ;
  LAYER VI2 ;
  RECT 4.740 147.220 4.940 147.420 ;
  LAYER VI2 ;
  RECT 4.340 147.220 4.540 147.420 ;
  LAYER VI3 ;
  RECT 4.280 150.900 5.140 151.180 ;
  LAYER VI3 ;
  RECT 4.740 150.900 4.940 151.100 ;
  LAYER VI3 ;
  RECT 4.340 150.900 4.540 151.100 ;
  LAYER VI2 ;
  RECT 4.280 150.900 5.140 151.180 ;
  LAYER VI2 ;
  RECT 4.740 150.900 4.940 151.100 ;
  LAYER VI2 ;
  RECT 4.340 150.900 4.540 151.100 ;
  LAYER VI3 ;
  RECT 4.280 154.580 5.140 154.860 ;
  LAYER VI3 ;
  RECT 4.740 154.580 4.940 154.780 ;
  LAYER VI3 ;
  RECT 4.340 154.580 4.540 154.780 ;
  LAYER VI2 ;
  RECT 4.280 154.580 5.140 154.860 ;
  LAYER VI2 ;
  RECT 4.740 154.580 4.940 154.780 ;
  LAYER VI2 ;
  RECT 4.340 154.580 4.540 154.780 ;
  LAYER VI3 ;
  RECT 4.280 158.260 5.140 158.540 ;
  LAYER VI3 ;
  RECT 4.740 158.260 4.940 158.460 ;
  LAYER VI3 ;
  RECT 4.340 158.260 4.540 158.460 ;
  LAYER VI2 ;
  RECT 4.280 158.260 5.140 158.540 ;
  LAYER VI2 ;
  RECT 4.740 158.260 4.940 158.460 ;
  LAYER VI2 ;
  RECT 4.340 158.260 4.540 158.460 ;
  LAYER VI3 ;
  RECT 4.280 161.940 5.140 162.220 ;
  LAYER VI3 ;
  RECT 4.740 161.940 4.940 162.140 ;
  LAYER VI3 ;
  RECT 4.340 161.940 4.540 162.140 ;
  LAYER VI2 ;
  RECT 4.280 161.940 5.140 162.220 ;
  LAYER VI2 ;
  RECT 4.740 161.940 4.940 162.140 ;
  LAYER VI2 ;
  RECT 4.340 161.940 4.540 162.140 ;
  LAYER VI3 ;
  RECT 4.280 165.620 5.140 165.900 ;
  LAYER VI3 ;
  RECT 4.740 165.620 4.940 165.820 ;
  LAYER VI3 ;
  RECT 4.340 165.620 4.540 165.820 ;
  LAYER VI2 ;
  RECT 4.280 165.620 5.140 165.900 ;
  LAYER VI2 ;
  RECT 4.740 165.620 4.940 165.820 ;
  LAYER VI2 ;
  RECT 4.340 165.620 4.540 165.820 ;
  LAYER VI3 ;
  RECT 4.280 169.300 5.140 169.580 ;
  LAYER VI3 ;
  RECT 4.740 169.300 4.940 169.500 ;
  LAYER VI3 ;
  RECT 4.340 169.300 4.540 169.500 ;
  LAYER VI2 ;
  RECT 4.280 169.300 5.140 169.580 ;
  LAYER VI2 ;
  RECT 4.740 169.300 4.940 169.500 ;
  LAYER VI2 ;
  RECT 4.340 169.300 4.540 169.500 ;
  LAYER VI3 ;
  RECT 4.280 172.980 5.140 173.260 ;
  LAYER VI3 ;
  RECT 4.740 172.980 4.940 173.180 ;
  LAYER VI3 ;
  RECT 4.340 172.980 4.540 173.180 ;
  LAYER VI2 ;
  RECT 4.280 172.980 5.140 173.260 ;
  LAYER VI2 ;
  RECT 4.740 172.980 4.940 173.180 ;
  LAYER VI2 ;
  RECT 4.340 172.980 4.540 173.180 ;
  LAYER VI3 ;
  RECT 4.280 176.660 5.140 176.940 ;
  LAYER VI3 ;
  RECT 4.740 176.660 4.940 176.860 ;
  LAYER VI3 ;
  RECT 4.340 176.660 4.540 176.860 ;
  LAYER VI2 ;
  RECT 4.280 176.660 5.140 176.940 ;
  LAYER VI2 ;
  RECT 4.740 176.660 4.940 176.860 ;
  LAYER VI2 ;
  RECT 4.340 176.660 4.540 176.860 ;
  LAYER VI3 ;
  RECT 4.280 180.340 5.140 180.620 ;
  LAYER VI3 ;
  RECT 4.740 180.340 4.940 180.540 ;
  LAYER VI3 ;
  RECT 4.340 180.340 4.540 180.540 ;
  LAYER VI2 ;
  RECT 4.280 180.340 5.140 180.620 ;
  LAYER VI2 ;
  RECT 4.740 180.340 4.940 180.540 ;
  LAYER VI2 ;
  RECT 4.340 180.340 4.540 180.540 ;
  LAYER VI3 ;
  RECT 4.280 184.020 5.140 184.300 ;
  LAYER VI3 ;
  RECT 4.740 184.020 4.940 184.220 ;
  LAYER VI3 ;
  RECT 4.340 184.020 4.540 184.220 ;
  LAYER VI2 ;
  RECT 4.280 184.020 5.140 184.300 ;
  LAYER VI2 ;
  RECT 4.740 184.020 4.940 184.220 ;
  LAYER VI2 ;
  RECT 4.340 184.020 4.540 184.220 ;
  LAYER VI3 ;
  RECT 4.280 187.700 5.140 187.980 ;
  LAYER VI3 ;
  RECT 4.740 187.700 4.940 187.900 ;
  LAYER VI3 ;
  RECT 4.340 187.700 4.540 187.900 ;
  LAYER VI2 ;
  RECT 4.280 187.700 5.140 187.980 ;
  LAYER VI2 ;
  RECT 4.740 187.700 4.940 187.900 ;
  LAYER VI2 ;
  RECT 4.340 187.700 4.540 187.900 ;
  LAYER VI3 ;
  RECT 4.280 191.380 5.140 191.660 ;
  LAYER VI3 ;
  RECT 4.740 191.380 4.940 191.580 ;
  LAYER VI3 ;
  RECT 4.340 191.380 4.540 191.580 ;
  LAYER VI2 ;
  RECT 4.280 191.380 5.140 191.660 ;
  LAYER VI2 ;
  RECT 4.740 191.380 4.940 191.580 ;
  LAYER VI2 ;
  RECT 4.340 191.380 4.540 191.580 ;
  LAYER VI3 ;
  RECT 4.280 195.060 5.140 195.340 ;
  LAYER VI3 ;
  RECT 4.740 195.060 4.940 195.260 ;
  LAYER VI3 ;
  RECT 4.340 195.060 4.540 195.260 ;
  LAYER VI2 ;
  RECT 4.280 195.060 5.140 195.340 ;
  LAYER VI2 ;
  RECT 4.740 195.060 4.940 195.260 ;
  LAYER VI2 ;
  RECT 4.340 195.060 4.540 195.260 ;
  LAYER VI3 ;
  RECT 4.280 198.740 5.140 199.020 ;
  LAYER VI3 ;
  RECT 4.740 198.740 4.940 198.940 ;
  LAYER VI3 ;
  RECT 4.340 198.740 4.540 198.940 ;
  LAYER VI2 ;
  RECT 4.280 198.740 5.140 199.020 ;
  LAYER VI2 ;
  RECT 4.740 198.740 4.940 198.940 ;
  LAYER VI2 ;
  RECT 4.340 198.740 4.540 198.940 ;
  LAYER VI3 ;
  RECT 4.280 202.420 5.140 202.700 ;
  LAYER VI3 ;
  RECT 4.740 202.420 4.940 202.620 ;
  LAYER VI3 ;
  RECT 4.340 202.420 4.540 202.620 ;
  LAYER VI2 ;
  RECT 4.280 202.420 5.140 202.700 ;
  LAYER VI2 ;
  RECT 4.740 202.420 4.940 202.620 ;
  LAYER VI2 ;
  RECT 4.340 202.420 4.540 202.620 ;
  LAYER VI3 ;
  RECT 4.280 206.100 5.140 206.380 ;
  LAYER VI3 ;
  RECT 4.740 206.100 4.940 206.300 ;
  LAYER VI3 ;
  RECT 4.340 206.100 4.540 206.300 ;
  LAYER VI2 ;
  RECT 4.280 206.100 5.140 206.380 ;
  LAYER VI2 ;
  RECT 4.740 206.100 4.940 206.300 ;
  LAYER VI2 ;
  RECT 4.340 206.100 4.540 206.300 ;
  LAYER VI3 ;
  RECT 4.280 209.780 5.140 210.060 ;
  LAYER VI3 ;
  RECT 4.740 209.780 4.940 209.980 ;
  LAYER VI3 ;
  RECT 4.340 209.780 4.540 209.980 ;
  LAYER VI2 ;
  RECT 4.280 209.780 5.140 210.060 ;
  LAYER VI2 ;
  RECT 4.740 209.780 4.940 209.980 ;
  LAYER VI2 ;
  RECT 4.340 209.780 4.540 209.980 ;
  LAYER VI3 ;
  RECT 4.280 213.460 5.140 213.740 ;
  LAYER VI3 ;
  RECT 4.740 213.460 4.940 213.660 ;
  LAYER VI3 ;
  RECT 4.340 213.460 4.540 213.660 ;
  LAYER VI2 ;
  RECT 4.280 213.460 5.140 213.740 ;
  LAYER VI2 ;
  RECT 4.740 213.460 4.940 213.660 ;
  LAYER VI2 ;
  RECT 4.340 213.460 4.540 213.660 ;
  LAYER VI3 ;
  RECT 4.280 217.140 5.140 217.420 ;
  LAYER VI3 ;
  RECT 4.740 217.140 4.940 217.340 ;
  LAYER VI3 ;
  RECT 4.340 217.140 4.540 217.340 ;
  LAYER VI2 ;
  RECT 4.280 217.140 5.140 217.420 ;
  LAYER VI2 ;
  RECT 4.740 217.140 4.940 217.340 ;
  LAYER VI2 ;
  RECT 4.340 217.140 4.540 217.340 ;
  LAYER VI3 ;
  RECT 4.280 220.820 5.140 221.100 ;
  LAYER VI3 ;
  RECT 4.740 220.820 4.940 221.020 ;
  LAYER VI3 ;
  RECT 4.340 220.820 4.540 221.020 ;
  LAYER VI2 ;
  RECT 4.280 220.820 5.140 221.100 ;
  LAYER VI2 ;
  RECT 4.740 220.820 4.940 221.020 ;
  LAYER VI2 ;
  RECT 4.340 220.820 4.540 221.020 ;
  LAYER VI3 ;
  RECT 4.280 224.500 5.140 224.780 ;
  LAYER VI3 ;
  RECT 4.740 224.500 4.940 224.700 ;
  LAYER VI3 ;
  RECT 4.340 224.500 4.540 224.700 ;
  LAYER VI2 ;
  RECT 4.280 224.500 5.140 224.780 ;
  LAYER VI2 ;
  RECT 4.740 224.500 4.940 224.700 ;
  LAYER VI2 ;
  RECT 4.340 224.500 4.540 224.700 ;
  LAYER VI3 ;
  RECT 4.280 228.180 5.140 228.460 ;
  LAYER VI3 ;
  RECT 4.740 228.180 4.940 228.380 ;
  LAYER VI3 ;
  RECT 4.340 228.180 4.540 228.380 ;
  LAYER VI2 ;
  RECT 4.280 228.180 5.140 228.460 ;
  LAYER VI2 ;
  RECT 4.740 228.180 4.940 228.380 ;
  LAYER VI2 ;
  RECT 4.340 228.180 4.540 228.380 ;
  LAYER VI3 ;
  RECT 4.280 231.860 5.140 232.140 ;
  LAYER VI3 ;
  RECT 4.740 231.860 4.940 232.060 ;
  LAYER VI3 ;
  RECT 4.340 231.860 4.540 232.060 ;
  LAYER VI2 ;
  RECT 4.280 231.860 5.140 232.140 ;
  LAYER VI2 ;
  RECT 4.740 231.860 4.940 232.060 ;
  LAYER VI2 ;
  RECT 4.340 231.860 4.540 232.060 ;
  LAYER VI3 ;
  RECT 4.280 235.540 5.140 235.820 ;
  LAYER VI3 ;
  RECT 4.740 235.540 4.940 235.740 ;
  LAYER VI3 ;
  RECT 4.340 235.540 4.540 235.740 ;
  LAYER VI2 ;
  RECT 4.280 235.540 5.140 235.820 ;
  LAYER VI2 ;
  RECT 4.740 235.540 4.940 235.740 ;
  LAYER VI2 ;
  RECT 4.340 235.540 4.540 235.740 ;
  LAYER VI3 ;
  RECT 4.280 239.220 5.140 239.500 ;
  LAYER VI3 ;
  RECT 4.740 239.220 4.940 239.420 ;
  LAYER VI3 ;
  RECT 4.340 239.220 4.540 239.420 ;
  LAYER VI2 ;
  RECT 4.280 239.220 5.140 239.500 ;
  LAYER VI2 ;
  RECT 4.740 239.220 4.940 239.420 ;
  LAYER VI2 ;
  RECT 4.340 239.220 4.540 239.420 ;
  LAYER VI3 ;
  RECT 4.280 242.900 5.140 243.180 ;
  LAYER VI3 ;
  RECT 4.740 242.900 4.940 243.100 ;
  LAYER VI3 ;
  RECT 4.340 242.900 4.540 243.100 ;
  LAYER VI2 ;
  RECT 4.280 242.900 5.140 243.180 ;
  LAYER VI2 ;
  RECT 4.740 242.900 4.940 243.100 ;
  LAYER VI2 ;
  RECT 4.340 242.900 4.540 243.100 ;
  LAYER VI3 ;
  RECT 4.280 246.580 5.140 246.860 ;
  LAYER VI3 ;
  RECT 4.740 246.580 4.940 246.780 ;
  LAYER VI3 ;
  RECT 4.340 246.580 4.540 246.780 ;
  LAYER VI2 ;
  RECT 4.280 246.580 5.140 246.860 ;
  LAYER VI2 ;
  RECT 4.740 246.580 4.940 246.780 ;
  LAYER VI2 ;
  RECT 4.340 246.580 4.540 246.780 ;
  LAYER VI3 ;
  RECT 4.280 250.260 5.140 250.540 ;
  LAYER VI3 ;
  RECT 4.740 250.260 4.940 250.460 ;
  LAYER VI3 ;
  RECT 4.340 250.260 4.540 250.460 ;
  LAYER VI2 ;
  RECT 4.280 250.260 5.140 250.540 ;
  LAYER VI2 ;
  RECT 4.740 250.260 4.940 250.460 ;
  LAYER VI2 ;
  RECT 4.340 250.260 4.540 250.460 ;
  LAYER VI3 ;
  RECT 4.280 253.940 5.140 254.220 ;
  LAYER VI3 ;
  RECT 4.740 253.940 4.940 254.140 ;
  LAYER VI3 ;
  RECT 4.340 253.940 4.540 254.140 ;
  LAYER VI2 ;
  RECT 4.280 253.940 5.140 254.220 ;
  LAYER VI2 ;
  RECT 4.740 253.940 4.940 254.140 ;
  LAYER VI2 ;
  RECT 4.340 253.940 4.540 254.140 ;
  LAYER VI3 ;
  RECT 4.280 257.620 5.140 257.900 ;
  LAYER VI3 ;
  RECT 4.740 257.620 4.940 257.820 ;
  LAYER VI3 ;
  RECT 4.340 257.620 4.540 257.820 ;
  LAYER VI2 ;
  RECT 4.280 257.620 5.140 257.900 ;
  LAYER VI2 ;
  RECT 4.740 257.620 4.940 257.820 ;
  LAYER VI2 ;
  RECT 4.340 257.620 4.540 257.820 ;
  LAYER VI3 ;
  RECT 4.280 261.300 5.140 261.580 ;
  LAYER VI3 ;
  RECT 4.740 261.300 4.940 261.500 ;
  LAYER VI3 ;
  RECT 4.340 261.300 4.540 261.500 ;
  LAYER VI2 ;
  RECT 4.280 261.300 5.140 261.580 ;
  LAYER VI2 ;
  RECT 4.740 261.300 4.940 261.500 ;
  LAYER VI2 ;
  RECT 4.340 261.300 4.540 261.500 ;
  LAYER VI3 ;
  RECT 4.280 264.980 5.140 265.260 ;
  LAYER VI3 ;
  RECT 4.740 264.980 4.940 265.180 ;
  LAYER VI3 ;
  RECT 4.340 264.980 4.540 265.180 ;
  LAYER VI2 ;
  RECT 4.280 264.980 5.140 265.260 ;
  LAYER VI2 ;
  RECT 4.740 264.980 4.940 265.180 ;
  LAYER VI2 ;
  RECT 4.340 264.980 4.540 265.180 ;
  LAYER VI3 ;
  RECT 4.280 268.660 5.140 268.940 ;
  LAYER VI3 ;
  RECT 4.740 268.660 4.940 268.860 ;
  LAYER VI3 ;
  RECT 4.340 268.660 4.540 268.860 ;
  LAYER VI2 ;
  RECT 4.280 268.660 5.140 268.940 ;
  LAYER VI2 ;
  RECT 4.740 268.660 4.940 268.860 ;
  LAYER VI2 ;
  RECT 4.340 268.660 4.540 268.860 ;
  LAYER VI3 ;
  RECT 4.280 272.340 5.140 272.620 ;
  LAYER VI3 ;
  RECT 4.740 272.340 4.940 272.540 ;
  LAYER VI3 ;
  RECT 4.340 272.340 4.540 272.540 ;
  LAYER VI2 ;
  RECT 4.280 272.340 5.140 272.620 ;
  LAYER VI2 ;
  RECT 4.740 272.340 4.940 272.540 ;
  LAYER VI2 ;
  RECT 4.340 272.340 4.540 272.540 ;
  LAYER VI3 ;
  RECT 4.280 276.020 5.140 276.300 ;
  LAYER VI3 ;
  RECT 4.740 276.020 4.940 276.220 ;
  LAYER VI3 ;
  RECT 4.340 276.020 4.540 276.220 ;
  LAYER VI2 ;
  RECT 4.280 276.020 5.140 276.300 ;
  LAYER VI2 ;
  RECT 4.740 276.020 4.940 276.220 ;
  LAYER VI2 ;
  RECT 4.340 276.020 4.540 276.220 ;
  LAYER VI3 ;
  RECT 4.280 279.700 5.140 279.980 ;
  LAYER VI3 ;
  RECT 4.740 279.700 4.940 279.900 ;
  LAYER VI3 ;
  RECT 4.340 279.700 4.540 279.900 ;
  LAYER VI2 ;
  RECT 4.280 279.700 5.140 279.980 ;
  LAYER VI2 ;
  RECT 4.740 279.700 4.940 279.900 ;
  LAYER VI2 ;
  RECT 4.340 279.700 4.540 279.900 ;
  LAYER VI3 ;
  RECT 4.280 283.380 5.140 283.660 ;
  LAYER VI3 ;
  RECT 4.740 283.380 4.940 283.580 ;
  LAYER VI3 ;
  RECT 4.340 283.380 4.540 283.580 ;
  LAYER VI2 ;
  RECT 4.280 283.380 5.140 283.660 ;
  LAYER VI2 ;
  RECT 4.740 283.380 4.940 283.580 ;
  LAYER VI2 ;
  RECT 4.340 283.380 4.540 283.580 ;
  LAYER VI3 ;
  RECT 4.280 287.060 5.140 287.340 ;
  LAYER VI3 ;
  RECT 4.740 287.060 4.940 287.260 ;
  LAYER VI3 ;
  RECT 4.340 287.060 4.540 287.260 ;
  LAYER VI2 ;
  RECT 4.280 287.060 5.140 287.340 ;
  LAYER VI2 ;
  RECT 4.740 287.060 4.940 287.260 ;
  LAYER VI2 ;
  RECT 4.340 287.060 4.540 287.260 ;
  LAYER VI3 ;
  RECT 4.280 290.740 5.140 291.020 ;
  LAYER VI3 ;
  RECT 4.740 290.740 4.940 290.940 ;
  LAYER VI3 ;
  RECT 4.340 290.740 4.540 290.940 ;
  LAYER VI2 ;
  RECT 4.280 290.740 5.140 291.020 ;
  LAYER VI2 ;
  RECT 4.740 290.740 4.940 290.940 ;
  LAYER VI2 ;
  RECT 4.340 290.740 4.540 290.940 ;
  LAYER VI3 ;
  RECT 4.280 294.420 5.140 294.700 ;
  LAYER VI3 ;
  RECT 4.740 294.420 4.940 294.620 ;
  LAYER VI3 ;
  RECT 4.340 294.420 4.540 294.620 ;
  LAYER VI2 ;
  RECT 4.280 294.420 5.140 294.700 ;
  LAYER VI2 ;
  RECT 4.740 294.420 4.940 294.620 ;
  LAYER VI2 ;
  RECT 4.340 294.420 4.540 294.620 ;
  LAYER VI3 ;
  RECT 4.280 298.100 5.140 298.380 ;
  LAYER VI3 ;
  RECT 4.740 298.100 4.940 298.300 ;
  LAYER VI3 ;
  RECT 4.340 298.100 4.540 298.300 ;
  LAYER VI2 ;
  RECT 4.280 298.100 5.140 298.380 ;
  LAYER VI2 ;
  RECT 4.740 298.100 4.940 298.300 ;
  LAYER VI2 ;
  RECT 4.340 298.100 4.540 298.300 ;
  LAYER VI3 ;
  RECT 4.280 301.780 5.140 302.060 ;
  LAYER VI3 ;
  RECT 4.740 301.780 4.940 301.980 ;
  LAYER VI3 ;
  RECT 4.340 301.780 4.540 301.980 ;
  LAYER VI2 ;
  RECT 4.280 301.780 5.140 302.060 ;
  LAYER VI2 ;
  RECT 4.740 301.780 4.940 301.980 ;
  LAYER VI2 ;
  RECT 4.340 301.780 4.540 301.980 ;
  LAYER VI3 ;
  RECT 4.280 305.460 5.140 305.740 ;
  LAYER VI3 ;
  RECT 4.740 305.460 4.940 305.660 ;
  LAYER VI3 ;
  RECT 4.340 305.460 4.540 305.660 ;
  LAYER VI2 ;
  RECT 4.280 305.460 5.140 305.740 ;
  LAYER VI2 ;
  RECT 4.740 305.460 4.940 305.660 ;
  LAYER VI2 ;
  RECT 4.340 305.460 4.540 305.660 ;
  LAYER VI3 ;
  RECT 4.280 309.140 5.140 309.420 ;
  LAYER VI3 ;
  RECT 4.740 309.140 4.940 309.340 ;
  LAYER VI3 ;
  RECT 4.340 309.140 4.540 309.340 ;
  LAYER VI2 ;
  RECT 4.280 309.140 5.140 309.420 ;
  LAYER VI2 ;
  RECT 4.740 309.140 4.940 309.340 ;
  LAYER VI2 ;
  RECT 4.340 309.140 4.540 309.340 ;
  LAYER VI3 ;
  RECT 4.280 312.820 5.140 313.100 ;
  LAYER VI3 ;
  RECT 4.740 312.820 4.940 313.020 ;
  LAYER VI3 ;
  RECT 4.340 312.820 4.540 313.020 ;
  LAYER VI2 ;
  RECT 4.280 312.820 5.140 313.100 ;
  LAYER VI2 ;
  RECT 4.740 312.820 4.940 313.020 ;
  LAYER VI2 ;
  RECT 4.340 312.820 4.540 313.020 ;
  LAYER VI3 ;
  RECT 4.280 316.500 5.140 316.780 ;
  LAYER VI3 ;
  RECT 4.740 316.500 4.940 316.700 ;
  LAYER VI3 ;
  RECT 4.340 316.500 4.540 316.700 ;
  LAYER VI2 ;
  RECT 4.280 316.500 5.140 316.780 ;
  LAYER VI2 ;
  RECT 4.740 316.500 4.940 316.700 ;
  LAYER VI2 ;
  RECT 4.340 316.500 4.540 316.700 ;
  LAYER VI3 ;
  RECT 4.280 320.180 5.140 320.460 ;
  LAYER VI3 ;
  RECT 4.740 320.180 4.940 320.380 ;
  LAYER VI3 ;
  RECT 4.340 320.180 4.540 320.380 ;
  LAYER VI2 ;
  RECT 4.280 320.180 5.140 320.460 ;
  LAYER VI2 ;
  RECT 4.740 320.180 4.940 320.380 ;
  LAYER VI2 ;
  RECT 4.340 320.180 4.540 320.380 ;
  LAYER VI3 ;
  RECT 4.280 323.860 5.140 324.140 ;
  LAYER VI3 ;
  RECT 4.740 323.860 4.940 324.060 ;
  LAYER VI3 ;
  RECT 4.340 323.860 4.540 324.060 ;
  LAYER VI2 ;
  RECT 4.280 323.860 5.140 324.140 ;
  LAYER VI2 ;
  RECT 4.740 323.860 4.940 324.060 ;
  LAYER VI2 ;
  RECT 4.340 323.860 4.540 324.060 ;
  LAYER VI3 ;
  RECT 4.280 327.540 5.140 327.820 ;
  LAYER VI3 ;
  RECT 4.740 327.540 4.940 327.740 ;
  LAYER VI3 ;
  RECT 4.340 327.540 4.540 327.740 ;
  LAYER VI2 ;
  RECT 4.280 327.540 5.140 327.820 ;
  LAYER VI2 ;
  RECT 4.740 327.540 4.940 327.740 ;
  LAYER VI2 ;
  RECT 4.340 327.540 4.540 327.740 ;
  LAYER VI3 ;
  RECT 4.280 331.220 5.140 331.500 ;
  LAYER VI3 ;
  RECT 4.740 331.220 4.940 331.420 ;
  LAYER VI3 ;
  RECT 4.340 331.220 4.540 331.420 ;
  LAYER VI2 ;
  RECT 4.280 331.220 5.140 331.500 ;
  LAYER VI2 ;
  RECT 4.740 331.220 4.940 331.420 ;
  LAYER VI2 ;
  RECT 4.340 331.220 4.540 331.420 ;
  LAYER VI3 ;
  RECT 4.280 334.900 5.140 335.180 ;
  LAYER VI3 ;
  RECT 4.740 334.900 4.940 335.100 ;
  LAYER VI3 ;
  RECT 4.340 334.900 4.540 335.100 ;
  LAYER VI2 ;
  RECT 4.280 334.900 5.140 335.180 ;
  LAYER VI2 ;
  RECT 4.740 334.900 4.940 335.100 ;
  LAYER VI2 ;
  RECT 4.340 334.900 4.540 335.100 ;
  LAYER VI3 ;
  RECT 4.280 338.580 5.140 338.860 ;
  LAYER VI3 ;
  RECT 4.740 338.580 4.940 338.780 ;
  LAYER VI3 ;
  RECT 4.340 338.580 4.540 338.780 ;
  LAYER VI2 ;
  RECT 4.280 338.580 5.140 338.860 ;
  LAYER VI2 ;
  RECT 4.740 338.580 4.940 338.780 ;
  LAYER VI2 ;
  RECT 4.340 338.580 4.540 338.780 ;
  LAYER VI3 ;
  RECT 4.280 342.260 5.140 342.540 ;
  LAYER VI3 ;
  RECT 4.740 342.260 4.940 342.460 ;
  LAYER VI3 ;
  RECT 4.340 342.260 4.540 342.460 ;
  LAYER VI2 ;
  RECT 4.280 342.260 5.140 342.540 ;
  LAYER VI2 ;
  RECT 4.740 342.260 4.940 342.460 ;
  LAYER VI2 ;
  RECT 4.340 342.260 4.540 342.460 ;
  LAYER VI3 ;
  RECT 4.280 345.940 5.140 346.220 ;
  LAYER VI3 ;
  RECT 4.740 345.940 4.940 346.140 ;
  LAYER VI3 ;
  RECT 4.340 345.940 4.540 346.140 ;
  LAYER VI2 ;
  RECT 4.280 345.940 5.140 346.220 ;
  LAYER VI2 ;
  RECT 4.740 345.940 4.940 346.140 ;
  LAYER VI2 ;
  RECT 4.340 345.940 4.540 346.140 ;
  LAYER VI3 ;
  RECT 4.280 349.620 5.140 349.900 ;
  LAYER VI3 ;
  RECT 4.740 349.620 4.940 349.820 ;
  LAYER VI3 ;
  RECT 4.340 349.620 4.540 349.820 ;
  LAYER VI2 ;
  RECT 4.280 349.620 5.140 349.900 ;
  LAYER VI2 ;
  RECT 4.740 349.620 4.940 349.820 ;
  LAYER VI2 ;
  RECT 4.340 349.620 4.540 349.820 ;
  LAYER VI3 ;
  RECT 4.280 353.300 5.140 353.580 ;
  LAYER VI3 ;
  RECT 4.740 353.300 4.940 353.500 ;
  LAYER VI3 ;
  RECT 4.340 353.300 4.540 353.500 ;
  LAYER VI2 ;
  RECT 4.280 353.300 5.140 353.580 ;
  LAYER VI2 ;
  RECT 4.740 353.300 4.940 353.500 ;
  LAYER VI2 ;
  RECT 4.340 353.300 4.540 353.500 ;
  LAYER VI3 ;
  RECT 4.280 356.980 5.140 357.260 ;
  LAYER VI3 ;
  RECT 4.740 356.980 4.940 357.180 ;
  LAYER VI3 ;
  RECT 4.340 356.980 4.540 357.180 ;
  LAYER VI2 ;
  RECT 4.280 356.980 5.140 357.260 ;
  LAYER VI2 ;
  RECT 4.740 356.980 4.940 357.180 ;
  LAYER VI2 ;
  RECT 4.340 356.980 4.540 357.180 ;
  LAYER VI3 ;
  RECT 4.280 360.660 5.140 360.940 ;
  LAYER VI3 ;
  RECT 4.740 360.660 4.940 360.860 ;
  LAYER VI3 ;
  RECT 4.340 360.660 4.540 360.860 ;
  LAYER VI2 ;
  RECT 4.280 360.660 5.140 360.940 ;
  LAYER VI2 ;
  RECT 4.740 360.660 4.940 360.860 ;
  LAYER VI2 ;
  RECT 4.340 360.660 4.540 360.860 ;
  LAYER VI3 ;
  RECT 4.280 364.340 5.140 364.620 ;
  LAYER VI3 ;
  RECT 4.740 364.340 4.940 364.540 ;
  LAYER VI3 ;
  RECT 4.340 364.340 4.540 364.540 ;
  LAYER VI2 ;
  RECT 4.280 364.340 5.140 364.620 ;
  LAYER VI2 ;
  RECT 4.740 364.340 4.940 364.540 ;
  LAYER VI2 ;
  RECT 4.340 364.340 4.540 364.540 ;
  LAYER VI3 ;
  RECT 4.280 368.020 5.140 368.300 ;
  LAYER VI3 ;
  RECT 4.740 368.020 4.940 368.220 ;
  LAYER VI3 ;
  RECT 4.340 368.020 4.540 368.220 ;
  LAYER VI2 ;
  RECT 4.280 368.020 5.140 368.300 ;
  LAYER VI2 ;
  RECT 4.740 368.020 4.940 368.220 ;
  LAYER VI2 ;
  RECT 4.340 368.020 4.540 368.220 ;
  LAYER VI3 ;
  RECT 4.280 371.700 5.140 371.980 ;
  LAYER VI3 ;
  RECT 4.740 371.700 4.940 371.900 ;
  LAYER VI3 ;
  RECT 4.340 371.700 4.540 371.900 ;
  LAYER VI2 ;
  RECT 4.280 371.700 5.140 371.980 ;
  LAYER VI2 ;
  RECT 4.740 371.700 4.940 371.900 ;
  LAYER VI2 ;
  RECT 4.340 371.700 4.540 371.900 ;
  LAYER VI3 ;
  RECT 4.280 375.380 5.140 375.660 ;
  LAYER VI3 ;
  RECT 4.740 375.380 4.940 375.580 ;
  LAYER VI3 ;
  RECT 4.340 375.380 4.540 375.580 ;
  LAYER VI2 ;
  RECT 4.280 375.380 5.140 375.660 ;
  LAYER VI2 ;
  RECT 4.740 375.380 4.940 375.580 ;
  LAYER VI2 ;
  RECT 4.340 375.380 4.540 375.580 ;
  LAYER VI3 ;
  RECT 4.280 379.060 5.140 379.340 ;
  LAYER VI3 ;
  RECT 4.740 379.060 4.940 379.260 ;
  LAYER VI3 ;
  RECT 4.340 379.060 4.540 379.260 ;
  LAYER VI2 ;
  RECT 4.280 379.060 5.140 379.340 ;
  LAYER VI2 ;
  RECT 4.740 379.060 4.940 379.260 ;
  LAYER VI2 ;
  RECT 4.340 379.060 4.540 379.260 ;
  LAYER VI3 ;
  RECT 4.280 382.740 5.140 383.020 ;
  LAYER VI3 ;
  RECT 4.740 382.740 4.940 382.940 ;
  LAYER VI3 ;
  RECT 4.340 382.740 4.540 382.940 ;
  LAYER VI2 ;
  RECT 4.280 382.740 5.140 383.020 ;
  LAYER VI2 ;
  RECT 4.740 382.740 4.940 382.940 ;
  LAYER VI2 ;
  RECT 4.340 382.740 4.540 382.940 ;
  LAYER VI3 ;
  RECT 4.280 386.420 5.140 386.700 ;
  LAYER VI3 ;
  RECT 4.740 386.420 4.940 386.620 ;
  LAYER VI3 ;
  RECT 4.340 386.420 4.540 386.620 ;
  LAYER VI2 ;
  RECT 4.280 386.420 5.140 386.700 ;
  LAYER VI2 ;
  RECT 4.740 386.420 4.940 386.620 ;
  LAYER VI2 ;
  RECT 4.340 386.420 4.540 386.620 ;
  LAYER VI3 ;
  RECT 4.280 390.100 5.140 390.380 ;
  LAYER VI3 ;
  RECT 4.740 390.100 4.940 390.300 ;
  LAYER VI3 ;
  RECT 4.340 390.100 4.540 390.300 ;
  LAYER VI2 ;
  RECT 4.280 390.100 5.140 390.380 ;
  LAYER VI2 ;
  RECT 4.740 390.100 4.940 390.300 ;
  LAYER VI2 ;
  RECT 4.340 390.100 4.540 390.300 ;
  LAYER VI3 ;
  RECT 4.280 393.780 5.140 394.060 ;
  LAYER VI3 ;
  RECT 4.740 393.780 4.940 393.980 ;
  LAYER VI3 ;
  RECT 4.340 393.780 4.540 393.980 ;
  LAYER VI2 ;
  RECT 4.280 393.780 5.140 394.060 ;
  LAYER VI2 ;
  RECT 4.740 393.780 4.940 393.980 ;
  LAYER VI2 ;
  RECT 4.340 393.780 4.540 393.980 ;
  LAYER VI3 ;
  RECT 4.280 397.460 5.140 397.740 ;
  LAYER VI3 ;
  RECT 4.740 397.460 4.940 397.660 ;
  LAYER VI3 ;
  RECT 4.340 397.460 4.540 397.660 ;
  LAYER VI2 ;
  RECT 4.280 397.460 5.140 397.740 ;
  LAYER VI2 ;
  RECT 4.740 397.460 4.940 397.660 ;
  LAYER VI2 ;
  RECT 4.340 397.460 4.540 397.660 ;
  LAYER VI3 ;
  RECT 4.280 401.140 5.140 401.420 ;
  LAYER VI3 ;
  RECT 4.740 401.140 4.940 401.340 ;
  LAYER VI3 ;
  RECT 4.340 401.140 4.540 401.340 ;
  LAYER VI2 ;
  RECT 4.280 401.140 5.140 401.420 ;
  LAYER VI2 ;
  RECT 4.740 401.140 4.940 401.340 ;
  LAYER VI2 ;
  RECT 4.340 401.140 4.540 401.340 ;
  LAYER VI3 ;
  RECT 4.280 404.820 5.140 405.100 ;
  LAYER VI3 ;
  RECT 4.740 404.820 4.940 405.020 ;
  LAYER VI3 ;
  RECT 4.340 404.820 4.540 405.020 ;
  LAYER VI2 ;
  RECT 4.280 404.820 5.140 405.100 ;
  LAYER VI2 ;
  RECT 4.740 404.820 4.940 405.020 ;
  LAYER VI2 ;
  RECT 4.340 404.820 4.540 405.020 ;
  LAYER VI3 ;
  RECT 4.280 408.500 5.140 408.780 ;
  LAYER VI3 ;
  RECT 4.740 408.500 4.940 408.700 ;
  LAYER VI3 ;
  RECT 4.340 408.500 4.540 408.700 ;
  LAYER VI2 ;
  RECT 4.280 408.500 5.140 408.780 ;
  LAYER VI2 ;
  RECT 4.740 408.500 4.940 408.700 ;
  LAYER VI2 ;
  RECT 4.340 408.500 4.540 408.700 ;
  LAYER VI3 ;
  RECT 4.280 412.180 5.140 412.460 ;
  LAYER VI3 ;
  RECT 4.740 412.180 4.940 412.380 ;
  LAYER VI3 ;
  RECT 4.340 412.180 4.540 412.380 ;
  LAYER VI2 ;
  RECT 4.280 412.180 5.140 412.460 ;
  LAYER VI2 ;
  RECT 4.740 412.180 4.940 412.380 ;
  LAYER VI2 ;
  RECT 4.340 412.180 4.540 412.380 ;
  LAYER VI3 ;
  RECT 4.280 415.860 5.140 416.140 ;
  LAYER VI3 ;
  RECT 4.740 415.860 4.940 416.060 ;
  LAYER VI3 ;
  RECT 4.340 415.860 4.540 416.060 ;
  LAYER VI2 ;
  RECT 4.280 415.860 5.140 416.140 ;
  LAYER VI2 ;
  RECT 4.740 415.860 4.940 416.060 ;
  LAYER VI2 ;
  RECT 4.340 415.860 4.540 416.060 ;
  LAYER VI3 ;
  RECT 4.280 419.540 5.140 419.820 ;
  LAYER VI3 ;
  RECT 4.740 419.540 4.940 419.740 ;
  LAYER VI3 ;
  RECT 4.340 419.540 4.540 419.740 ;
  LAYER VI2 ;
  RECT 4.280 419.540 5.140 419.820 ;
  LAYER VI2 ;
  RECT 4.740 419.540 4.940 419.740 ;
  LAYER VI2 ;
  RECT 4.340 419.540 4.540 419.740 ;
  LAYER VI3 ;
  RECT 4.280 423.220 5.140 423.500 ;
  LAYER VI3 ;
  RECT 4.740 423.220 4.940 423.420 ;
  LAYER VI3 ;
  RECT 4.340 423.220 4.540 423.420 ;
  LAYER VI2 ;
  RECT 4.280 423.220 5.140 423.500 ;
  LAYER VI2 ;
  RECT 4.740 423.220 4.940 423.420 ;
  LAYER VI2 ;
  RECT 4.340 423.220 4.540 423.420 ;
  LAYER VI3 ;
  RECT 4.280 426.900 5.140 427.180 ;
  LAYER VI3 ;
  RECT 4.740 426.900 4.940 427.100 ;
  LAYER VI3 ;
  RECT 4.340 426.900 4.540 427.100 ;
  LAYER VI2 ;
  RECT 4.280 426.900 5.140 427.180 ;
  LAYER VI2 ;
  RECT 4.740 426.900 4.940 427.100 ;
  LAYER VI2 ;
  RECT 4.340 426.900 4.540 427.100 ;
  LAYER VI3 ;
  RECT 4.280 430.580 5.140 430.860 ;
  LAYER VI3 ;
  RECT 4.740 430.580 4.940 430.780 ;
  LAYER VI3 ;
  RECT 4.340 430.580 4.540 430.780 ;
  LAYER VI2 ;
  RECT 4.280 430.580 5.140 430.860 ;
  LAYER VI2 ;
  RECT 4.740 430.580 4.940 430.780 ;
  LAYER VI2 ;
  RECT 4.340 430.580 4.540 430.780 ;
  LAYER VI3 ;
  RECT 4.280 434.260 5.140 434.540 ;
  LAYER VI3 ;
  RECT 4.740 434.260 4.940 434.460 ;
  LAYER VI3 ;
  RECT 4.340 434.260 4.540 434.460 ;
  LAYER VI2 ;
  RECT 4.280 434.260 5.140 434.540 ;
  LAYER VI2 ;
  RECT 4.740 434.260 4.940 434.460 ;
  LAYER VI2 ;
  RECT 4.340 434.260 4.540 434.460 ;
  LAYER VI3 ;
  RECT 4.280 437.940 5.140 438.220 ;
  LAYER VI3 ;
  RECT 4.740 437.940 4.940 438.140 ;
  LAYER VI3 ;
  RECT 4.340 437.940 4.540 438.140 ;
  LAYER VI2 ;
  RECT 4.280 437.940 5.140 438.220 ;
  LAYER VI2 ;
  RECT 4.740 437.940 4.940 438.140 ;
  LAYER VI2 ;
  RECT 4.340 437.940 4.540 438.140 ;
  LAYER VI3 ;
  RECT 4.280 441.620 5.140 441.900 ;
  LAYER VI3 ;
  RECT 4.740 441.620 4.940 441.820 ;
  LAYER VI3 ;
  RECT 4.340 441.620 4.540 441.820 ;
  LAYER VI2 ;
  RECT 4.280 441.620 5.140 441.900 ;
  LAYER VI2 ;
  RECT 4.740 441.620 4.940 441.820 ;
  LAYER VI2 ;
  RECT 4.340 441.620 4.540 441.820 ;
  LAYER VI3 ;
  RECT 4.280 445.300 5.140 445.580 ;
  LAYER VI3 ;
  RECT 4.740 445.300 4.940 445.500 ;
  LAYER VI3 ;
  RECT 4.340 445.300 4.540 445.500 ;
  LAYER VI2 ;
  RECT 4.280 445.300 5.140 445.580 ;
  LAYER VI2 ;
  RECT 4.740 445.300 4.940 445.500 ;
  LAYER VI2 ;
  RECT 4.340 445.300 4.540 445.500 ;
  LAYER VI3 ;
  RECT 4.280 448.980 5.140 449.260 ;
  LAYER VI3 ;
  RECT 4.740 448.980 4.940 449.180 ;
  LAYER VI3 ;
  RECT 4.340 448.980 4.540 449.180 ;
  LAYER VI2 ;
  RECT 4.280 448.980 5.140 449.260 ;
  LAYER VI2 ;
  RECT 4.740 448.980 4.940 449.180 ;
  LAYER VI2 ;
  RECT 4.340 448.980 4.540 449.180 ;
  LAYER VI3 ;
  RECT 4.280 452.660 5.140 452.940 ;
  LAYER VI3 ;
  RECT 4.740 452.660 4.940 452.860 ;
  LAYER VI3 ;
  RECT 4.340 452.660 4.540 452.860 ;
  LAYER VI2 ;
  RECT 4.280 452.660 5.140 452.940 ;
  LAYER VI2 ;
  RECT 4.740 452.660 4.940 452.860 ;
  LAYER VI2 ;
  RECT 4.340 452.660 4.540 452.860 ;
  LAYER VI3 ;
  RECT 4.280 456.340 5.140 456.620 ;
  LAYER VI3 ;
  RECT 4.740 456.340 4.940 456.540 ;
  LAYER VI3 ;
  RECT 4.340 456.340 4.540 456.540 ;
  LAYER VI2 ;
  RECT 4.280 456.340 5.140 456.620 ;
  LAYER VI2 ;
  RECT 4.740 456.340 4.940 456.540 ;
  LAYER VI2 ;
  RECT 4.340 456.340 4.540 456.540 ;
  LAYER VI3 ;
  RECT 4.280 460.020 5.140 460.300 ;
  LAYER VI3 ;
  RECT 4.740 460.020 4.940 460.220 ;
  LAYER VI3 ;
  RECT 4.340 460.020 4.540 460.220 ;
  LAYER VI2 ;
  RECT 4.280 460.020 5.140 460.300 ;
  LAYER VI2 ;
  RECT 4.740 460.020 4.940 460.220 ;
  LAYER VI2 ;
  RECT 4.340 460.020 4.540 460.220 ;
  LAYER VI3 ;
  RECT 4.280 463.700 5.140 463.980 ;
  LAYER VI3 ;
  RECT 4.740 463.700 4.940 463.900 ;
  LAYER VI3 ;
  RECT 4.340 463.700 4.540 463.900 ;
  LAYER VI2 ;
  RECT 4.280 463.700 5.140 463.980 ;
  LAYER VI2 ;
  RECT 4.740 463.700 4.940 463.900 ;
  LAYER VI2 ;
  RECT 4.340 463.700 4.540 463.900 ;
  LAYER VI3 ;
  RECT 4.280 467.380 5.140 467.660 ;
  LAYER VI3 ;
  RECT 4.740 467.380 4.940 467.580 ;
  LAYER VI3 ;
  RECT 4.340 467.380 4.540 467.580 ;
  LAYER VI2 ;
  RECT 4.280 467.380 5.140 467.660 ;
  LAYER VI2 ;
  RECT 4.740 467.380 4.940 467.580 ;
  LAYER VI2 ;
  RECT 4.340 467.380 4.540 467.580 ;
  LAYER VI3 ;
  RECT 4.280 471.060 5.140 471.340 ;
  LAYER VI3 ;
  RECT 4.740 471.060 4.940 471.260 ;
  LAYER VI3 ;
  RECT 4.340 471.060 4.540 471.260 ;
  LAYER VI2 ;
  RECT 4.280 471.060 5.140 471.340 ;
  LAYER VI2 ;
  RECT 4.740 471.060 4.940 471.260 ;
  LAYER VI2 ;
  RECT 4.340 471.060 4.540 471.260 ;
  LAYER VI3 ;
  RECT 4.280 474.740 5.140 475.020 ;
  LAYER VI3 ;
  RECT 4.740 474.740 4.940 474.940 ;
  LAYER VI3 ;
  RECT 4.340 474.740 4.540 474.940 ;
  LAYER VI2 ;
  RECT 4.280 474.740 5.140 475.020 ;
  LAYER VI2 ;
  RECT 4.740 474.740 4.940 474.940 ;
  LAYER VI2 ;
  RECT 4.340 474.740 4.540 474.940 ;
  LAYER VI3 ;
  RECT 4.280 478.420 5.140 478.700 ;
  LAYER VI3 ;
  RECT 4.740 478.420 4.940 478.620 ;
  LAYER VI3 ;
  RECT 4.340 478.420 4.540 478.620 ;
  LAYER VI2 ;
  RECT 4.280 478.420 5.140 478.700 ;
  LAYER VI2 ;
  RECT 4.740 478.420 4.940 478.620 ;
  LAYER VI2 ;
  RECT 4.340 478.420 4.540 478.620 ;
  LAYER VI3 ;
  RECT 4.280 482.100 5.140 482.380 ;
  LAYER VI3 ;
  RECT 4.740 482.100 4.940 482.300 ;
  LAYER VI3 ;
  RECT 4.340 482.100 4.540 482.300 ;
  LAYER VI2 ;
  RECT 4.280 482.100 5.140 482.380 ;
  LAYER VI2 ;
  RECT 4.740 482.100 4.940 482.300 ;
  LAYER VI2 ;
  RECT 4.340 482.100 4.540 482.300 ;
  LAYER VI3 ;
  RECT 4.280 485.780 5.140 486.060 ;
  LAYER VI3 ;
  RECT 4.740 485.780 4.940 485.980 ;
  LAYER VI3 ;
  RECT 4.340 485.780 4.540 485.980 ;
  LAYER VI2 ;
  RECT 4.280 485.780 5.140 486.060 ;
  LAYER VI2 ;
  RECT 4.740 485.780 4.940 485.980 ;
  LAYER VI2 ;
  RECT 4.340 485.780 4.540 485.980 ;
  LAYER VI3 ;
  RECT 4.280 489.460 5.140 489.740 ;
  LAYER VI3 ;
  RECT 4.740 489.460 4.940 489.660 ;
  LAYER VI3 ;
  RECT 4.340 489.460 4.540 489.660 ;
  LAYER VI2 ;
  RECT 4.280 489.460 5.140 489.740 ;
  LAYER VI2 ;
  RECT 4.740 489.460 4.940 489.660 ;
  LAYER VI2 ;
  RECT 4.340 489.460 4.540 489.660 ;
  LAYER VI3 ;
  RECT 4.280 493.140 5.140 493.420 ;
  LAYER VI3 ;
  RECT 4.740 493.140 4.940 493.340 ;
  LAYER VI3 ;
  RECT 4.340 493.140 4.540 493.340 ;
  LAYER VI2 ;
  RECT 4.280 493.140 5.140 493.420 ;
  LAYER VI2 ;
  RECT 4.740 493.140 4.940 493.340 ;
  LAYER VI2 ;
  RECT 4.340 493.140 4.540 493.340 ;
  LAYER VI3 ;
  RECT 4.280 496.820 5.140 497.100 ;
  LAYER VI3 ;
  RECT 4.740 496.820 4.940 497.020 ;
  LAYER VI3 ;
  RECT 4.340 496.820 4.540 497.020 ;
  LAYER VI2 ;
  RECT 4.280 496.820 5.140 497.100 ;
  LAYER VI2 ;
  RECT 4.740 496.820 4.940 497.020 ;
  LAYER VI2 ;
  RECT 4.340 496.820 4.540 497.020 ;
  LAYER VI3 ;
  RECT 4.280 500.500 5.140 500.780 ;
  LAYER VI3 ;
  RECT 4.740 500.500 4.940 500.700 ;
  LAYER VI3 ;
  RECT 4.340 500.500 4.540 500.700 ;
  LAYER VI2 ;
  RECT 4.280 500.500 5.140 500.780 ;
  LAYER VI2 ;
  RECT 4.740 500.500 4.940 500.700 ;
  LAYER VI2 ;
  RECT 4.340 500.500 4.540 500.700 ;
  LAYER VI3 ;
  RECT 4.280 504.180 5.140 504.460 ;
  LAYER VI3 ;
  RECT 4.740 504.180 4.940 504.380 ;
  LAYER VI3 ;
  RECT 4.340 504.180 4.540 504.380 ;
  LAYER VI2 ;
  RECT 4.280 504.180 5.140 504.460 ;
  LAYER VI2 ;
  RECT 4.740 504.180 4.940 504.380 ;
  LAYER VI2 ;
  RECT 4.340 504.180 4.540 504.380 ;
  LAYER VI3 ;
  RECT 4.280 507.860 5.140 508.140 ;
  LAYER VI3 ;
  RECT 4.740 507.860 4.940 508.060 ;
  LAYER VI3 ;
  RECT 4.340 507.860 4.540 508.060 ;
  LAYER VI2 ;
  RECT 4.280 507.860 5.140 508.140 ;
  LAYER VI2 ;
  RECT 4.740 507.860 4.940 508.060 ;
  LAYER VI2 ;
  RECT 4.340 507.860 4.540 508.060 ;
  LAYER VI3 ;
  RECT 4.280 511.540 5.140 511.820 ;
  LAYER VI3 ;
  RECT 4.740 511.540 4.940 511.740 ;
  LAYER VI3 ;
  RECT 4.340 511.540 4.540 511.740 ;
  LAYER VI2 ;
  RECT 4.280 511.540 5.140 511.820 ;
  LAYER VI2 ;
  RECT 4.740 511.540 4.940 511.740 ;
  LAYER VI2 ;
  RECT 4.340 511.540 4.540 511.740 ;
  LAYER VI3 ;
  RECT 4.280 515.220 5.140 515.500 ;
  LAYER VI3 ;
  RECT 4.740 515.220 4.940 515.420 ;
  LAYER VI3 ;
  RECT 4.340 515.220 4.540 515.420 ;
  LAYER VI2 ;
  RECT 4.280 515.220 5.140 515.500 ;
  LAYER VI2 ;
  RECT 4.740 515.220 4.940 515.420 ;
  LAYER VI2 ;
  RECT 4.340 515.220 4.540 515.420 ;
  LAYER VI3 ;
  RECT 4.280 518.900 5.140 519.180 ;
  LAYER VI3 ;
  RECT 4.740 518.900 4.940 519.100 ;
  LAYER VI3 ;
  RECT 4.340 518.900 4.540 519.100 ;
  LAYER VI2 ;
  RECT 4.280 518.900 5.140 519.180 ;
  LAYER VI2 ;
  RECT 4.740 518.900 4.940 519.100 ;
  LAYER VI2 ;
  RECT 4.340 518.900 4.540 519.100 ;
  LAYER VI3 ;
  RECT 4.280 522.580 5.140 522.860 ;
  LAYER VI3 ;
  RECT 4.740 522.580 4.940 522.780 ;
  LAYER VI3 ;
  RECT 4.340 522.580 4.540 522.780 ;
  LAYER VI2 ;
  RECT 4.280 522.580 5.140 522.860 ;
  LAYER VI2 ;
  RECT 4.740 522.580 4.940 522.780 ;
  LAYER VI2 ;
  RECT 4.340 522.580 4.540 522.780 ;
  LAYER VI3 ;
  RECT 4.280 526.260 5.140 526.540 ;
  LAYER VI3 ;
  RECT 4.740 526.260 4.940 526.460 ;
  LAYER VI3 ;
  RECT 4.340 526.260 4.540 526.460 ;
  LAYER VI2 ;
  RECT 4.280 526.260 5.140 526.540 ;
  LAYER VI2 ;
  RECT 4.740 526.260 4.940 526.460 ;
  LAYER VI2 ;
  RECT 4.340 526.260 4.540 526.460 ;
  LAYER VI3 ;
  RECT 4.280 529.940 5.140 530.220 ;
  LAYER VI3 ;
  RECT 4.740 529.940 4.940 530.140 ;
  LAYER VI3 ;
  RECT 4.340 529.940 4.540 530.140 ;
  LAYER VI2 ;
  RECT 4.280 529.940 5.140 530.220 ;
  LAYER VI2 ;
  RECT 4.740 529.940 4.940 530.140 ;
  LAYER VI2 ;
  RECT 4.340 529.940 4.540 530.140 ;
  LAYER VI3 ;
  RECT 4.280 533.620 5.140 533.900 ;
  LAYER VI3 ;
  RECT 4.740 533.620 4.940 533.820 ;
  LAYER VI3 ;
  RECT 4.340 533.620 4.540 533.820 ;
  LAYER VI2 ;
  RECT 4.280 533.620 5.140 533.900 ;
  LAYER VI2 ;
  RECT 4.740 533.620 4.940 533.820 ;
  LAYER VI2 ;
  RECT 4.340 533.620 4.540 533.820 ;
  LAYER VI3 ;
  RECT 4.280 537.300 5.140 537.580 ;
  LAYER VI3 ;
  RECT 4.740 537.300 4.940 537.500 ;
  LAYER VI3 ;
  RECT 4.340 537.300 4.540 537.500 ;
  LAYER VI2 ;
  RECT 4.280 537.300 5.140 537.580 ;
  LAYER VI2 ;
  RECT 4.740 537.300 4.940 537.500 ;
  LAYER VI2 ;
  RECT 4.340 537.300 4.540 537.500 ;
  LAYER VI3 ;
  RECT 4.280 540.980 5.140 541.260 ;
  LAYER VI3 ;
  RECT 4.740 540.980 4.940 541.180 ;
  LAYER VI3 ;
  RECT 4.340 540.980 4.540 541.180 ;
  LAYER VI2 ;
  RECT 4.280 540.980 5.140 541.260 ;
  LAYER VI2 ;
  RECT 4.740 540.980 4.940 541.180 ;
  LAYER VI2 ;
  RECT 4.340 540.980 4.540 541.180 ;
  LAYER VI3 ;
  RECT 4.280 544.660 5.140 544.940 ;
  LAYER VI3 ;
  RECT 4.740 544.660 4.940 544.860 ;
  LAYER VI3 ;
  RECT 4.340 544.660 4.540 544.860 ;
  LAYER VI2 ;
  RECT 4.280 544.660 5.140 544.940 ;
  LAYER VI2 ;
  RECT 4.740 544.660 4.940 544.860 ;
  LAYER VI2 ;
  RECT 4.340 544.660 4.540 544.860 ;
  LAYER VI3 ;
  RECT 4.280 548.340 5.140 548.620 ;
  LAYER VI3 ;
  RECT 4.740 548.340 4.940 548.540 ;
  LAYER VI3 ;
  RECT 4.340 548.340 4.540 548.540 ;
  LAYER VI2 ;
  RECT 4.280 548.340 5.140 548.620 ;
  LAYER VI2 ;
  RECT 4.740 548.340 4.940 548.540 ;
  LAYER VI2 ;
  RECT 4.340 548.340 4.540 548.540 ;
  LAYER VI3 ;
  RECT 4.280 552.020 5.140 552.300 ;
  LAYER VI3 ;
  RECT 4.740 552.020 4.940 552.220 ;
  LAYER VI3 ;
  RECT 4.340 552.020 4.540 552.220 ;
  LAYER VI2 ;
  RECT 4.280 552.020 5.140 552.300 ;
  LAYER VI2 ;
  RECT 4.740 552.020 4.940 552.220 ;
  LAYER VI2 ;
  RECT 4.340 552.020 4.540 552.220 ;
  LAYER VI3 ;
  RECT 4.280 559.940 5.140 560.320 ;
  LAYER VI3 ;
  RECT 4.680 560.000 4.880 560.200 ;
  LAYER VI3 ;
  RECT 4.280 560.000 4.480 560.200 ;
  LAYER VI2 ;
  RECT 4.280 559.940 5.140 560.320 ;
  LAYER VI2 ;
  RECT 4.680 560.000 4.880 560.200 ;
  LAYER VI2 ;
  RECT 4.280 560.000 4.480 560.200 ;
  LAYER VI3 ;
  RECT 47.350 560.790 47.600 561.650 ;
  LAYER VI3 ;
  RECT 47.350 561.250 47.550 561.450 ;
  LAYER VI3 ;
  RECT 47.350 560.850 47.550 561.050 ;
  LAYER VI2 ;
  RECT 47.350 560.790 47.600 561.650 ;
  LAYER VI2 ;
  RECT 47.350 561.250 47.550 561.450 ;
  LAYER VI2 ;
  RECT 47.350 560.850 47.550 561.050 ;
  LAYER VI3 ;
  RECT 88.270 560.790 88.520 561.650 ;
  LAYER VI3 ;
  RECT 88.270 561.250 88.470 561.450 ;
  LAYER VI3 ;
  RECT 88.270 560.850 88.470 561.050 ;
  LAYER VI2 ;
  RECT 88.270 560.790 88.520 561.650 ;
  LAYER VI2 ;
  RECT 88.270 561.250 88.470 561.450 ;
  LAYER VI2 ;
  RECT 88.270 560.850 88.470 561.050 ;
  LAYER VI3 ;
  RECT 129.190 560.790 129.440 561.650 ;
  LAYER VI3 ;
  RECT 129.190 561.250 129.390 561.450 ;
  LAYER VI3 ;
  RECT 129.190 560.850 129.390 561.050 ;
  LAYER VI2 ;
  RECT 129.190 560.790 129.440 561.650 ;
  LAYER VI2 ;
  RECT 129.190 561.250 129.390 561.450 ;
  LAYER VI2 ;
  RECT 129.190 560.850 129.390 561.050 ;
  LAYER VI3 ;
  RECT 170.110 560.790 170.360 561.650 ;
  LAYER VI3 ;
  RECT 170.110 561.250 170.310 561.450 ;
  LAYER VI3 ;
  RECT 170.110 560.850 170.310 561.050 ;
  LAYER VI2 ;
  RECT 170.110 560.790 170.360 561.650 ;
  LAYER VI2 ;
  RECT 170.110 561.250 170.310 561.450 ;
  LAYER VI2 ;
  RECT 170.110 560.850 170.310 561.050 ;
  LAYER VI3 ;
  RECT 211.030 560.790 211.280 561.650 ;
  LAYER VI3 ;
  RECT 211.030 561.250 211.230 561.450 ;
  LAYER VI3 ;
  RECT 211.030 560.850 211.230 561.050 ;
  LAYER VI2 ;
  RECT 211.030 560.790 211.280 561.650 ;
  LAYER VI2 ;
  RECT 211.030 561.250 211.230 561.450 ;
  LAYER VI2 ;
  RECT 211.030 560.850 211.230 561.050 ;
  LAYER VI3 ;
  RECT 251.950 560.790 252.200 561.650 ;
  LAYER VI3 ;
  RECT 251.950 561.250 252.150 561.450 ;
  LAYER VI3 ;
  RECT 251.950 560.850 252.150 561.050 ;
  LAYER VI2 ;
  RECT 251.950 560.790 252.200 561.650 ;
  LAYER VI2 ;
  RECT 251.950 561.250 252.150 561.450 ;
  LAYER VI2 ;
  RECT 251.950 560.850 252.150 561.050 ;
  LAYER VI3 ;
  RECT 292.870 560.790 293.120 561.650 ;
  LAYER VI3 ;
  RECT 292.870 561.250 293.070 561.450 ;
  LAYER VI3 ;
  RECT 292.870 560.850 293.070 561.050 ;
  LAYER VI2 ;
  RECT 292.870 560.790 293.120 561.650 ;
  LAYER VI2 ;
  RECT 292.870 561.250 293.070 561.450 ;
  LAYER VI2 ;
  RECT 292.870 560.850 293.070 561.050 ;
  LAYER VI3 ;
  RECT 333.790 560.790 334.040 561.650 ;
  LAYER VI3 ;
  RECT 333.790 561.250 333.990 561.450 ;
  LAYER VI3 ;
  RECT 333.790 560.850 333.990 561.050 ;
  LAYER VI2 ;
  RECT 333.790 560.790 334.040 561.650 ;
  LAYER VI2 ;
  RECT 333.790 561.250 333.990 561.450 ;
  LAYER VI2 ;
  RECT 333.790 560.850 333.990 561.050 ;
  LAYER VI3 ;
  RECT 374.710 560.790 374.960 561.650 ;
  LAYER VI3 ;
  RECT 374.710 561.250 374.910 561.450 ;
  LAYER VI3 ;
  RECT 374.710 560.850 374.910 561.050 ;
  LAYER VI2 ;
  RECT 374.710 560.790 374.960 561.650 ;
  LAYER VI2 ;
  RECT 374.710 561.250 374.910 561.450 ;
  LAYER VI2 ;
  RECT 374.710 560.850 374.910 561.050 ;
  LAYER VI3 ;
  RECT 415.630 560.790 415.880 561.650 ;
  LAYER VI3 ;
  RECT 415.630 561.250 415.830 561.450 ;
  LAYER VI3 ;
  RECT 415.630 560.850 415.830 561.050 ;
  LAYER VI2 ;
  RECT 415.630 560.790 415.880 561.650 ;
  LAYER VI2 ;
  RECT 415.630 561.250 415.830 561.450 ;
  LAYER VI2 ;
  RECT 415.630 560.850 415.830 561.050 ;
  LAYER VI3 ;
  RECT 456.550 560.790 456.800 561.650 ;
  LAYER VI3 ;
  RECT 456.550 561.250 456.750 561.450 ;
  LAYER VI3 ;
  RECT 456.550 560.850 456.750 561.050 ;
  LAYER VI2 ;
  RECT 456.550 560.790 456.800 561.650 ;
  LAYER VI2 ;
  RECT 456.550 561.250 456.750 561.450 ;
  LAYER VI2 ;
  RECT 456.550 560.850 456.750 561.050 ;
  LAYER VI3 ;
  RECT 497.470 560.790 497.720 561.650 ;
  LAYER VI3 ;
  RECT 497.470 561.250 497.670 561.450 ;
  LAYER VI3 ;
  RECT 497.470 560.850 497.670 561.050 ;
  LAYER VI2 ;
  RECT 497.470 560.790 497.720 561.650 ;
  LAYER VI2 ;
  RECT 497.470 561.250 497.670 561.450 ;
  LAYER VI2 ;
  RECT 497.470 560.850 497.670 561.050 ;
  LAYER VI3 ;
  RECT 538.390 560.790 538.640 561.650 ;
  LAYER VI3 ;
  RECT 538.390 561.250 538.590 561.450 ;
  LAYER VI3 ;
  RECT 538.390 560.850 538.590 561.050 ;
  LAYER VI2 ;
  RECT 538.390 560.790 538.640 561.650 ;
  LAYER VI2 ;
  RECT 538.390 561.250 538.590 561.450 ;
  LAYER VI2 ;
  RECT 538.390 560.850 538.590 561.050 ;
  LAYER VI3 ;
  RECT 579.310 560.790 579.560 561.650 ;
  LAYER VI3 ;
  RECT 579.310 561.250 579.510 561.450 ;
  LAYER VI3 ;
  RECT 579.310 560.850 579.510 561.050 ;
  LAYER VI2 ;
  RECT 579.310 560.790 579.560 561.650 ;
  LAYER VI2 ;
  RECT 579.310 561.250 579.510 561.450 ;
  LAYER VI2 ;
  RECT 579.310 560.850 579.510 561.050 ;
  LAYER VI3 ;
  RECT 620.230 560.790 620.480 561.650 ;
  LAYER VI3 ;
  RECT 620.230 561.250 620.430 561.450 ;
  LAYER VI3 ;
  RECT 620.230 560.850 620.430 561.050 ;
  LAYER VI2 ;
  RECT 620.230 560.790 620.480 561.650 ;
  LAYER VI2 ;
  RECT 620.230 561.250 620.430 561.450 ;
  LAYER VI2 ;
  RECT 620.230 560.850 620.430 561.050 ;
  LAYER VI3 ;
  RECT 661.150 560.790 661.400 561.650 ;
  LAYER VI3 ;
  RECT 661.150 561.250 661.350 561.450 ;
  LAYER VI3 ;
  RECT 661.150 560.850 661.350 561.050 ;
  LAYER VI2 ;
  RECT 661.150 560.790 661.400 561.650 ;
  LAYER VI2 ;
  RECT 661.150 561.250 661.350 561.450 ;
  LAYER VI2 ;
  RECT 661.150 560.850 661.350 561.050 ;
  LAYER VI3 ;
  RECT 702.070 560.790 702.320 561.650 ;
  LAYER VI3 ;
  RECT 702.070 561.250 702.270 561.450 ;
  LAYER VI3 ;
  RECT 702.070 560.850 702.270 561.050 ;
  LAYER VI2 ;
  RECT 702.070 560.790 702.320 561.650 ;
  LAYER VI2 ;
  RECT 702.070 561.250 702.270 561.450 ;
  LAYER VI2 ;
  RECT 702.070 560.850 702.270 561.050 ;
  LAYER VI3 ;
  RECT 742.990 560.790 743.240 561.650 ;
  LAYER VI3 ;
  RECT 742.990 561.250 743.190 561.450 ;
  LAYER VI3 ;
  RECT 742.990 560.850 743.190 561.050 ;
  LAYER VI2 ;
  RECT 742.990 560.790 743.240 561.650 ;
  LAYER VI2 ;
  RECT 742.990 561.250 743.190 561.450 ;
  LAYER VI2 ;
  RECT 742.990 560.850 743.190 561.050 ;
  LAYER VI3 ;
  RECT 783.910 560.790 784.160 561.650 ;
  LAYER VI3 ;
  RECT 783.910 561.250 784.110 561.450 ;
  LAYER VI3 ;
  RECT 783.910 560.850 784.110 561.050 ;
  LAYER VI2 ;
  RECT 783.910 560.790 784.160 561.650 ;
  LAYER VI2 ;
  RECT 783.910 561.250 784.110 561.450 ;
  LAYER VI2 ;
  RECT 783.910 560.850 784.110 561.050 ;
  LAYER VI3 ;
  RECT 824.830 560.790 825.080 561.650 ;
  LAYER VI3 ;
  RECT 824.830 561.250 825.030 561.450 ;
  LAYER VI3 ;
  RECT 824.830 560.850 825.030 561.050 ;
  LAYER VI2 ;
  RECT 824.830 560.790 825.080 561.650 ;
  LAYER VI2 ;
  RECT 824.830 561.250 825.030 561.450 ;
  LAYER VI2 ;
  RECT 824.830 560.850 825.030 561.050 ;
  LAYER VI3 ;
  RECT 865.750 560.790 866.000 561.650 ;
  LAYER VI3 ;
  RECT 865.750 561.250 865.950 561.450 ;
  LAYER VI3 ;
  RECT 865.750 560.850 865.950 561.050 ;
  LAYER VI2 ;
  RECT 865.750 560.790 866.000 561.650 ;
  LAYER VI2 ;
  RECT 865.750 561.250 865.950 561.450 ;
  LAYER VI2 ;
  RECT 865.750 560.850 865.950 561.050 ;
  LAYER VI3 ;
  RECT 906.670 560.790 906.920 561.650 ;
  LAYER VI3 ;
  RECT 906.670 561.250 906.870 561.450 ;
  LAYER VI3 ;
  RECT 906.670 560.850 906.870 561.050 ;
  LAYER VI2 ;
  RECT 906.670 560.790 906.920 561.650 ;
  LAYER VI2 ;
  RECT 906.670 561.250 906.870 561.450 ;
  LAYER VI2 ;
  RECT 906.670 560.850 906.870 561.050 ;
  LAYER VI3 ;
  RECT 947.590 560.790 947.840 561.650 ;
  LAYER VI3 ;
  RECT 947.590 561.250 947.790 561.450 ;
  LAYER VI3 ;
  RECT 947.590 560.850 947.790 561.050 ;
  LAYER VI2 ;
  RECT 947.590 560.790 947.840 561.650 ;
  LAYER VI2 ;
  RECT 947.590 561.250 947.790 561.450 ;
  LAYER VI2 ;
  RECT 947.590 560.850 947.790 561.050 ;
  LAYER VI3 ;
  RECT 988.510 560.790 988.760 561.650 ;
  LAYER VI3 ;
  RECT 988.510 561.250 988.710 561.450 ;
  LAYER VI3 ;
  RECT 988.510 560.850 988.710 561.050 ;
  LAYER VI2 ;
  RECT 988.510 560.790 988.760 561.650 ;
  LAYER VI2 ;
  RECT 988.510 561.250 988.710 561.450 ;
  LAYER VI2 ;
  RECT 988.510 560.850 988.710 561.050 ;
  LAYER VI3 ;
  RECT 1029.430 560.790 1029.680 561.650 ;
  LAYER VI3 ;
  RECT 1029.430 561.250 1029.630 561.450 ;
  LAYER VI3 ;
  RECT 1029.430 560.850 1029.630 561.050 ;
  LAYER VI2 ;
  RECT 1029.430 560.790 1029.680 561.650 ;
  LAYER VI2 ;
  RECT 1029.430 561.250 1029.630 561.450 ;
  LAYER VI2 ;
  RECT 1029.430 560.850 1029.630 561.050 ;
  LAYER VI3 ;
  RECT 1070.350 560.790 1070.600 561.650 ;
  LAYER VI3 ;
  RECT 1070.350 561.250 1070.550 561.450 ;
  LAYER VI3 ;
  RECT 1070.350 560.850 1070.550 561.050 ;
  LAYER VI2 ;
  RECT 1070.350 560.790 1070.600 561.650 ;
  LAYER VI2 ;
  RECT 1070.350 561.250 1070.550 561.450 ;
  LAYER VI2 ;
  RECT 1070.350 560.850 1070.550 561.050 ;
  LAYER VI3 ;
  RECT 1111.270 560.790 1111.520 561.650 ;
  LAYER VI3 ;
  RECT 1111.270 561.250 1111.470 561.450 ;
  LAYER VI3 ;
  RECT 1111.270 560.850 1111.470 561.050 ;
  LAYER VI2 ;
  RECT 1111.270 560.790 1111.520 561.650 ;
  LAYER VI2 ;
  RECT 1111.270 561.250 1111.470 561.450 ;
  LAYER VI2 ;
  RECT 1111.270 560.850 1111.470 561.050 ;
  LAYER VI3 ;
  RECT 1152.190 560.790 1152.440 561.650 ;
  LAYER VI3 ;
  RECT 1152.190 561.250 1152.390 561.450 ;
  LAYER VI3 ;
  RECT 1152.190 560.850 1152.390 561.050 ;
  LAYER VI2 ;
  RECT 1152.190 560.790 1152.440 561.650 ;
  LAYER VI2 ;
  RECT 1152.190 561.250 1152.390 561.450 ;
  LAYER VI2 ;
  RECT 1152.190 560.850 1152.390 561.050 ;
  LAYER VI3 ;
  RECT 1193.110 560.790 1193.360 561.650 ;
  LAYER VI3 ;
  RECT 1193.110 561.250 1193.310 561.450 ;
  LAYER VI3 ;
  RECT 1193.110 560.850 1193.310 561.050 ;
  LAYER VI2 ;
  RECT 1193.110 560.790 1193.360 561.650 ;
  LAYER VI2 ;
  RECT 1193.110 561.250 1193.310 561.450 ;
  LAYER VI2 ;
  RECT 1193.110 560.850 1193.310 561.050 ;
  LAYER VI3 ;
  RECT 1234.030 560.790 1234.280 561.650 ;
  LAYER VI3 ;
  RECT 1234.030 561.250 1234.230 561.450 ;
  LAYER VI3 ;
  RECT 1234.030 560.850 1234.230 561.050 ;
  LAYER VI2 ;
  RECT 1234.030 560.790 1234.280 561.650 ;
  LAYER VI2 ;
  RECT 1234.030 561.250 1234.230 561.450 ;
  LAYER VI2 ;
  RECT 1234.030 560.850 1234.230 561.050 ;
  LAYER VI3 ;
  RECT 1274.950 560.790 1275.200 561.650 ;
  LAYER VI3 ;
  RECT 1274.950 561.250 1275.150 561.450 ;
  LAYER VI3 ;
  RECT 1274.950 560.850 1275.150 561.050 ;
  LAYER VI2 ;
  RECT 1274.950 560.790 1275.200 561.650 ;
  LAYER VI2 ;
  RECT 1274.950 561.250 1275.150 561.450 ;
  LAYER VI2 ;
  RECT 1274.950 560.850 1275.150 561.050 ;
END
END SHKD110_4224X8X16BM1
END LIBRARY





