# ________________________________________________________________________________________________
# 
# 
#             Synchronous One-Port Register File Compiler
# 
#                 UMC 0.11um LL AE Logic Process
# 
# ________________________________________________________________________________________________
# 
#               
#         Copyright (C) 2024 Faraday Technology Corporation. All Rights Reserved.       
#                
#         This source code is an unpublished work belongs to Faraday Technology Corporation       
#         It is considered a trade secret and is not to be divulged or       
#         used by parties who have not received written authorization from       
#         Faraday Technology Corporation       
#                
#         Faraday's home page can be found at: http://www.faraday-tech.com/       
#                
# ________________________________________________________________________________________________
# 
#        IP Name            :  FSR0K_B_SY                
#        IP Version         :  1.4.0                     
#        IP Release Status  :  Active                    
#        Word               :  128                       
#        Bit                :  7                         
#        Byte               :  1                         
#        Mux                :  4                         
#        Output Loading     :  0.01                      
#        Clock Input Slew   :  0.016                     
#        Data Input Slew    :  0.016                     
#        Ring Type          :  Ringless Model            
#        Ring Width         :  0                         
#        Bus Format         :  0                         
#        Memaker Path       :  /home/mem/Desktop/memlib  
#        GUI Version        :  m20230904                 
#        Date               :  2024/09/06 21:04:36       
# ________________________________________________________________________________________________
# 

VERSION 5.5 ;
NAMESCASESENSITIVE ON ;
MACRO SYKB110_128X7X1CM4
CLASS BLOCK ;
FOREIGN SYKB110_128X7X1CM4 0.000 0.000 ;
ORIGIN 0.000 0.000 ;
SIZE 99.555 BY 68.179 ;
SYMMETRY x y r90 ;
SITE core ;
PIN VCC
  DIRECTION INOUT ;
  USE POWER ;
 PORT
  LAYER ME4 ;
  RECT 69.257 0.000 69.977 33.870 ;
 END
 PORT
  LAYER ME4 ;
  RECT 65.253 0.000 65.973 33.870 ;
 END
 PORT
  LAYER ME4 ;
  RECT 77.265 0.000 77.985 33.870 ;
 END
 PORT
  LAYER ME4 ;
  RECT 73.261 0.000 73.981 33.870 ;
 END
 PORT
  LAYER ME4 ;
  RECT 85.273 0.000 85.993 33.870 ;
 END
 PORT
  LAYER ME4 ;
  RECT 81.269 0.000 81.989 33.870 ;
 END
 PORT
  LAYER ME4 ;
  RECT 93.281 0.000 94.001 33.870 ;
 END
 PORT
  LAYER ME4 ;
  RECT 89.277 0.000 89.997 33.870 ;
 END
 PORT
  LAYER ME4 ;
  RECT 98.255 0.000 98.635 68.179 ;
 END
 PORT
  LAYER ME4 ;
  RECT 62.621 0.921 63.001 68.179 ;
 END
 PORT
  LAYER ME4 ;
  RECT 48.365 0.000 48.965 68.179 ;
 END
 PORT
  LAYER ME4 ;
  RECT 52.545 0.000 53.265 68.179 ;
 END
 PORT
  LAYER ME4 ;
  RECT 54.655 0.000 55.775 68.179 ;
 END
 PORT
  LAYER ME4 ;
  RECT 60.685 0.000 61.405 68.179 ;
 END
 PORT
  LAYER ME4 ;
  RECT 41.420 0.000 42.540 68.179 ;
 END
 PORT
  LAYER ME4 ;
  RECT 44.135 0.000 44.855 68.179 ;
 END
 PORT
  LAYER ME4 ;
  RECT 39.046 0.000 39.766 67.420 ;
 END
 PORT
  LAYER ME4 ;
  RECT 37.006 0.921 37.726 68.179 ;
 END
 PORT
  LAYER ME4 ;
  RECT 34.886 0.000 35.606 68.179 ;
 END
 PORT
  LAYER ME4 ;
  RECT 32.846 0.921 33.566 68.179 ;
 END
 PORT
  LAYER ME4 ;
  RECT 0.920 0.000 1.300 68.179 ;
 END
 PORT
  LAYER ME4 ;
  RECT 7.556 0.000 8.276 33.870 ;
 END
 PORT
  LAYER ME4 ;
  RECT 3.552 0.000 4.272 33.870 ;
 END
 PORT
  LAYER ME4 ;
  RECT 15.564 0.000 16.284 33.870 ;
 END
 PORT
  LAYER ME4 ;
  RECT 11.560 0.000 12.280 33.870 ;
 END
 PORT
  LAYER ME4 ;
  RECT 23.572 0.000 24.292 33.870 ;
 END
 PORT
  LAYER ME4 ;
  RECT 19.568 0.000 20.288 33.870 ;
 END
 PORT
  LAYER ME4 ;
  RECT 30.726 0.000 31.446 68.179 ;
 END
 PORT
  LAYER ME4 ;
  RECT 28.546 0.000 28.926 68.179 ;
 END
 PORT
  LAYER ME4 ;
  RECT 71.449 35.220 71.789 68.179 ;
 END
 PORT
  LAYER ME4 ;
  RECT 69.447 35.220 69.787 68.179 ;
 END
 PORT
  LAYER ME4 ;
  RECT 67.445 35.220 67.785 68.179 ;
 END
 PORT
  LAYER ME4 ;
  RECT 65.443 35.220 65.783 68.179 ;
 END
 PORT
  LAYER ME4 ;
  RECT 79.457 35.220 79.797 68.179 ;
 END
 PORT
  LAYER ME4 ;
  RECT 77.455 35.220 77.795 68.179 ;
 END
 PORT
  LAYER ME4 ;
  RECT 75.453 35.220 75.793 68.179 ;
 END
 PORT
  LAYER ME4 ;
  RECT 73.451 35.220 73.791 68.179 ;
 END
 PORT
  LAYER ME4 ;
  RECT 87.465 35.220 87.805 68.179 ;
 END
 PORT
  LAYER ME4 ;
  RECT 85.463 35.220 85.803 68.179 ;
 END
 PORT
  LAYER ME4 ;
  RECT 83.461 35.220 83.801 68.179 ;
 END
 PORT
  LAYER ME4 ;
  RECT 81.459 35.220 81.799 68.179 ;
 END
 PORT
  LAYER ME4 ;
  RECT 95.473 35.220 95.813 68.179 ;
 END
 PORT
  LAYER ME4 ;
  RECT 93.471 35.220 93.811 68.179 ;
 END
 PORT
  LAYER ME4 ;
  RECT 91.469 35.220 91.809 68.179 ;
 END
 PORT
  LAYER ME4 ;
  RECT 89.467 35.220 89.807 68.179 ;
 END
 PORT
  LAYER ME4 ;
  RECT 9.748 35.220 10.088 68.179 ;
 END
 PORT
  LAYER ME4 ;
  RECT 7.746 35.220 8.086 68.179 ;
 END
 PORT
  LAYER ME4 ;
  RECT 5.744 35.220 6.084 68.179 ;
 END
 PORT
  LAYER ME4 ;
  RECT 3.742 35.220 4.082 68.179 ;
 END
 PORT
  LAYER ME4 ;
  RECT 17.756 35.220 18.096 68.179 ;
 END
 PORT
  LAYER ME4 ;
  RECT 15.754 35.220 16.094 68.179 ;
 END
 PORT
  LAYER ME4 ;
  RECT 13.752 35.220 14.092 68.179 ;
 END
 PORT
  LAYER ME4 ;
  RECT 11.750 35.220 12.090 68.179 ;
 END
 PORT
  LAYER ME4 ;
  RECT 25.764 35.220 26.104 68.179 ;
 END
 PORT
  LAYER ME4 ;
  RECT 23.762 35.220 24.102 68.179 ;
 END
 PORT
  LAYER ME4 ;
  RECT 21.760 35.220 22.100 68.179 ;
 END
 PORT
  LAYER ME4 ;
  RECT 19.758 35.220 20.098 68.179 ;
 END
END VCC
PIN GND
  DIRECTION INOUT ;
  USE GROUND ;
 PORT
  LAYER ME4 ;
  RECT 64.442 0.921 64.782 68.179 ;
 END
 PORT
  LAYER ME4 ;
  RECT 71.259 0.000 71.979 31.570 ;
 END
 PORT
  LAYER ME4 ;
  RECT 72.450 0.000 72.790 68.179 ;
 END
 PORT
  LAYER ME4 ;
  RECT 66.444 0.000 66.784 68.179 ;
 END
 PORT
  LAYER ME4 ;
  RECT 67.255 0.000 67.975 31.570 ;
 END
 PORT
  LAYER ME4 ;
  RECT 68.446 0.921 68.786 68.179 ;
 END
 PORT
  LAYER ME4 ;
  RECT 70.448 0.921 70.788 68.179 ;
 END
 PORT
  LAYER ME4 ;
  RECT 79.267 0.000 79.987 31.570 ;
 END
 PORT
  LAYER ME4 ;
  RECT 80.458 0.000 80.798 68.179 ;
 END
 PORT
  LAYER ME4 ;
  RECT 74.452 0.000 74.792 68.179 ;
 END
 PORT
  LAYER ME4 ;
  RECT 75.263 0.000 75.983 31.570 ;
 END
 PORT
  LAYER ME4 ;
  RECT 76.454 0.921 76.794 68.179 ;
 END
 PORT
  LAYER ME4 ;
  RECT 78.456 0.921 78.796 68.179 ;
 END
 PORT
  LAYER ME4 ;
  RECT 87.275 0.000 87.995 31.570 ;
 END
 PORT
  LAYER ME4 ;
  RECT 88.466 0.000 88.806 68.179 ;
 END
 PORT
  LAYER ME4 ;
  RECT 82.460 0.000 82.800 68.179 ;
 END
 PORT
  LAYER ME4 ;
  RECT 83.271 0.000 83.991 31.570 ;
 END
 PORT
  LAYER ME4 ;
  RECT 84.462 0.921 84.802 68.179 ;
 END
 PORT
  LAYER ME4 ;
  RECT 86.464 0.921 86.804 68.179 ;
 END
 PORT
  LAYER ME4 ;
  RECT 95.283 0.000 96.003 31.570 ;
 END
 PORT
  LAYER ME4 ;
  RECT 96.474 0.000 96.814 68.179 ;
 END
 PORT
  LAYER ME4 ;
  RECT 90.468 0.000 90.808 68.179 ;
 END
 PORT
  LAYER ME4 ;
  RECT 91.279 0.000 91.999 31.570 ;
 END
 PORT
  LAYER ME4 ;
  RECT 92.470 0.921 92.810 68.179 ;
 END
 PORT
  LAYER ME4 ;
  RECT 94.472 0.921 94.812 68.179 ;
 END
 PORT
  LAYER ME4 ;
  RECT 97.475 0.000 97.815 68.179 ;
 END
 PORT
  LAYER ME4 ;
  RECT 63.441 0.921 63.781 68.179 ;
 END
 PORT
  LAYER ME4 ;
  RECT 45.585 0.000 46.305 68.179 ;
 END
 PORT
  LAYER ME4 ;
  RECT 51.579 0.000 52.299 68.179 ;
 END
 PORT
  LAYER ME4 ;
  RECT 57.050 0.000 57.770 68.179 ;
 END
 PORT
  LAYER ME4 ;
  RECT 58.765 0.000 59.485 68.179 ;
 END
 PORT
  LAYER ME4 ;
  RECT 61.761 0.000 62.361 68.179 ;
 END
 PORT
  LAYER ME4 ;
  RECT 38.026 0.000 38.746 68.179 ;
 END
 PORT
  LAYER ME4 ;
  RECT 35.986 0.921 36.706 67.420 ;
 END
 PORT
  LAYER ME4 ;
  RECT 33.866 0.000 34.586 68.179 ;
 END
 PORT
  LAYER ME4 ;
  RECT 31.826 0.921 32.546 68.179 ;
 END
 PORT
  LAYER ME4 ;
  RECT 1.740 0.000 2.080 68.179 ;
 END
 PORT
  LAYER ME4 ;
  RECT 2.741 0.921 3.081 68.179 ;
 END
 PORT
  LAYER ME4 ;
  RECT 9.558 0.000 10.278 31.570 ;
 END
 PORT
  LAYER ME4 ;
  RECT 10.749 0.000 11.089 68.179 ;
 END
 PORT
  LAYER ME4 ;
  RECT 4.743 0.000 5.083 68.179 ;
 END
 PORT
  LAYER ME4 ;
  RECT 5.554 0.000 6.274 31.570 ;
 END
 PORT
  LAYER ME4 ;
  RECT 6.745 0.921 7.085 68.179 ;
 END
 PORT
  LAYER ME4 ;
  RECT 8.747 0.921 9.087 68.179 ;
 END
 PORT
  LAYER ME4 ;
  RECT 17.566 0.000 18.286 31.570 ;
 END
 PORT
  LAYER ME4 ;
  RECT 18.757 0.000 19.097 68.179 ;
 END
 PORT
  LAYER ME4 ;
  RECT 12.751 0.000 13.091 68.179 ;
 END
 PORT
  LAYER ME4 ;
  RECT 13.562 0.000 14.282 31.570 ;
 END
 PORT
  LAYER ME4 ;
  RECT 14.753 0.921 15.093 68.179 ;
 END
 PORT
  LAYER ME4 ;
  RECT 16.755 0.921 17.095 68.179 ;
 END
 PORT
  LAYER ME4 ;
  RECT 25.574 0.000 26.294 31.570 ;
 END
 PORT
  LAYER ME4 ;
  RECT 26.765 0.000 27.105 68.179 ;
 END
 PORT
  LAYER ME4 ;
  RECT 20.759 0.000 21.099 68.179 ;
 END
 PORT
  LAYER ME4 ;
  RECT 21.570 0.000 22.290 31.570 ;
 END
 PORT
  LAYER ME4 ;
  RECT 22.761 0.921 23.101 68.179 ;
 END
 PORT
  LAYER ME4 ;
  RECT 24.763 0.921 25.103 68.179 ;
 END
 PORT
  LAYER ME4 ;
  RECT 29.706 0.000 30.426 68.179 ;
 END
 PORT
  LAYER ME4 ;
  RECT 27.766 0.000 28.106 68.179 ;
 END
END GND
PIN DI2
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 24.622 0.000 24.902 0.720 ;
  LAYER ME3 ;
  RECT 24.622 0.000 24.902 0.720 ;
  LAYER ME2 ;
  RECT 24.622 0.000 24.902 0.720 ;
  LAYER ME1 ;
  RECT 24.622 0.000 24.902 0.720 ;
 END
 ANTENNAPARTIALMETALAREA                  0.522 LAYER ME1 ;
 ANTENNAGATEAREA                          0.072 LAYER ME1 ;
 ANTENNAGATEAREA                          0.072 LAYER ME2 ;
 ANTENNAGATEAREA                          0.072 LAYER ME3 ;
 ANTENNAGATEAREA                          0.072 LAYER ME4 ;
 ANTENNADIFFAREA                          0.218 LAYER ME1 ;
 ANTENNADIFFAREA                          0.218 LAYER ME2 ;
 ANTENNADIFFAREA                          0.218 LAYER ME3 ;
 ANTENNADIFFAREA                          0.218 LAYER ME4 ;
 ANTENNAMAXAREACAR                       10.048 LAYER ME1 ;
 ANTENNAMAXAREACAR                       12.848 LAYER ME2 ;
 ANTENNAMAXAREACAR                       15.648 LAYER ME3 ;
 ANTENNAMAXAREACAR                       18.448 LAYER ME4 ;
END DI2
PIN DO2
  DIRECTION OUTPUT ;
 PORT
  LAYER ME4 ;
  RECT 22.564 0.000 22.844 0.720 ;
  LAYER ME3 ;
  RECT 22.564 0.000 22.844 0.720 ;
  LAYER ME2 ;
  RECT 22.564 0.000 22.844 0.720 ;
  LAYER ME1 ;
  RECT 22.564 0.000 22.844 0.720 ;
 END
 ANTENNAPARTIALMETALAREA                  2.030 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME3 ;
 ANTENNADIFFAREA                          1.293 LAYER ME4 ;
END DO2
PIN DI1
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 16.614 0.000 16.894 0.720 ;
  LAYER ME3 ;
  RECT 16.614 0.000 16.894 0.720 ;
  LAYER ME2 ;
  RECT 16.614 0.000 16.894 0.720 ;
  LAYER ME1 ;
  RECT 16.614 0.000 16.894 0.720 ;
 END
 ANTENNAPARTIALMETALAREA                  0.805 LAYER ME1 ;
 ANTENNAGATEAREA                          0.072 LAYER ME1 ;
 ANTENNAGATEAREA                          0.072 LAYER ME2 ;
 ANTENNAGATEAREA                          0.072 LAYER ME3 ;
 ANTENNAGATEAREA                          0.072 LAYER ME4 ;
 ANTENNADIFFAREA                          0.218 LAYER ME1 ;
 ANTENNADIFFAREA                          0.218 LAYER ME2 ;
 ANTENNADIFFAREA                          0.218 LAYER ME3 ;
 ANTENNADIFFAREA                          0.218 LAYER ME4 ;
 ANTENNAMAXAREACAR                       13.984 LAYER ME1 ;
 ANTENNAMAXAREACAR                       16.784 LAYER ME2 ;
 ANTENNAMAXAREACAR                       19.584 LAYER ME3 ;
 ANTENNAMAXAREACAR                       22.384 LAYER ME4 ;
END DI1
PIN DO1
  DIRECTION OUTPUT ;
 PORT
  LAYER ME4 ;
  RECT 14.636 0.000 14.916 0.720 ;
  LAYER ME3 ;
  RECT 14.636 0.000 14.916 0.720 ;
  LAYER ME2 ;
  RECT 14.636 0.000 14.916 0.720 ;
  LAYER ME1 ;
  RECT 14.636 0.000 14.916 0.720 ;
 END
 ANTENNAPARTIALMETALAREA                  2.030 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME3 ;
 ANTENNADIFFAREA                          1.293 LAYER ME4 ;
END DO1
PIN DI0
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 8.606 0.000 8.886 0.720 ;
  LAYER ME3 ;
  RECT 8.606 0.000 8.886 0.720 ;
  LAYER ME2 ;
  RECT 8.606 0.000 8.886 0.720 ;
  LAYER ME1 ;
  RECT 8.606 0.000 8.886 0.720 ;
 END
 ANTENNAPARTIALMETALAREA                  0.805 LAYER ME1 ;
 ANTENNAGATEAREA                          0.072 LAYER ME1 ;
 ANTENNAGATEAREA                          0.072 LAYER ME2 ;
 ANTENNAGATEAREA                          0.072 LAYER ME3 ;
 ANTENNAGATEAREA                          0.072 LAYER ME4 ;
 ANTENNADIFFAREA                          0.218 LAYER ME1 ;
 ANTENNADIFFAREA                          0.218 LAYER ME2 ;
 ANTENNADIFFAREA                          0.218 LAYER ME3 ;
 ANTENNADIFFAREA                          0.218 LAYER ME4 ;
 ANTENNAMAXAREACAR                       13.984 LAYER ME1 ;
 ANTENNAMAXAREACAR                       16.784 LAYER ME2 ;
 ANTENNAMAXAREACAR                       19.584 LAYER ME3 ;
 ANTENNAMAXAREACAR                       22.384 LAYER ME4 ;
END DI0
PIN DO0
  DIRECTION OUTPUT ;
 PORT
  LAYER ME4 ;
  RECT 6.628 0.000 6.908 0.720 ;
  LAYER ME3 ;
  RECT 6.628 0.000 6.908 0.720 ;
  LAYER ME2 ;
  RECT 6.628 0.000 6.908 0.720 ;
  LAYER ME1 ;
  RECT 6.628 0.000 6.908 0.720 ;
 END
 ANTENNAPARTIALMETALAREA                  2.030 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME3 ;
 ANTENNADIFFAREA                          1.293 LAYER ME4 ;
END DO0
PIN A2
  DIRECTION INPUT ;
 PORT
  LAYER ME3 ;
  RECT 42.908 0.000 43.228 0.600 ;
  LAYER ME2 ;
  RECT 42.908 0.000 43.228 0.600 ;
  LAYER ME1 ;
  RECT 42.908 0.000 43.228 0.600 ;
 END
 ANTENNAPARTIALMETALAREA                  1.067 LAYER ME2 ;
 ANTENNAGATEAREA                          0.144 LAYER ME2 ;
 ANTENNAGATEAREA                          0.144 LAYER ME3 ;
 ANTENNADIFFAREA                          0.218 LAYER ME2 ;
 ANTENNADIFFAREA                          0.218 LAYER ME3 ;
 ANTENNAMAXAREACAR                        9.746 LAYER ME2 ;
 ANTENNAMAXAREACAR                       11.079 LAYER ME3 ;
END A2
PIN A3
  DIRECTION INPUT ;
 PORT
  LAYER ME3 ;
  RECT 43.495 0.000 43.815 0.600 ;
  LAYER ME2 ;
  RECT 43.495 0.000 43.815 0.600 ;
  LAYER ME1 ;
  RECT 43.495 0.000 43.815 0.600 ;
 END
 ANTENNAPARTIALMETALAREA                  1.188 LAYER ME2 ;
 ANTENNAGATEAREA                          0.144 LAYER ME2 ;
 ANTENNAGATEAREA                          0.144 LAYER ME3 ;
 ANTENNADIFFAREA                          0.218 LAYER ME2 ;
 ANTENNADIFFAREA                          0.218 LAYER ME3 ;
 ANTENNAMAXAREACAR                       10.582 LAYER ME2 ;
 ANTENNAMAXAREACAR                       11.915 LAYER ME3 ;
END A3
PIN A4
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 36.656 0.000 36.976 0.600 ;
  LAYER ME3 ;
  RECT 36.656 0.000 36.976 0.600 ;
  LAYER ME2 ;
  RECT 36.656 0.000 36.976 0.600 ;
  LAYER ME1 ;
  RECT 36.656 0.000 36.976 0.600 ;
 END
 ANTENNAPARTIALMETALAREA                  1.910 LAYER ME2 ;
 ANTENNAGATEAREA                          0.180 LAYER ME2 ;
 ANTENNAGATEAREA                          0.180 LAYER ME3 ;
 ANTENNAGATEAREA                          0.180 LAYER ME4 ;
 ANTENNADIFFAREA                          0.218 LAYER ME2 ;
 ANTENNADIFFAREA                          0.218 LAYER ME3 ;
 ANTENNADIFFAREA                          0.218 LAYER ME4 ;
 ANTENNAMAXAREACAR                       13.456 LAYER ME2 ;
 ANTENNAMAXAREACAR                       14.522 LAYER ME3 ;
 ANTENNAMAXAREACAR                       15.589 LAYER ME4 ;
END A4
PIN A5
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 36.036 0.000 36.356 0.600 ;
  LAYER ME3 ;
  RECT 36.036 0.000 36.356 0.600 ;
  LAYER ME2 ;
  RECT 36.036 0.000 36.356 0.600 ;
  LAYER ME1 ;
  RECT 36.036 0.000 36.356 0.600 ;
 END
 ANTENNAPARTIALMETALAREA                  1.447 LAYER ME2 ;
 ANTENNAGATEAREA                          0.180 LAYER ME2 ;
 ANTENNAGATEAREA                          0.180 LAYER ME3 ;
 ANTENNAGATEAREA                          0.180 LAYER ME4 ;
 ANTENNADIFFAREA                          0.218 LAYER ME2 ;
 ANTENNADIFFAREA                          0.218 LAYER ME3 ;
 ANTENNADIFFAREA                          0.218 LAYER ME4 ;
 ANTENNAMAXAREACAR                       12.818 LAYER ME2 ;
 ANTENNAMAXAREACAR                       13.884 LAYER ME3 ;
 ANTENNAMAXAREACAR                       14.951 LAYER ME4 ;
END A5
PIN A6
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 32.556 0.000 32.876 0.600 ;
  LAYER ME3 ;
  RECT 32.556 0.000 32.876 0.600 ;
  LAYER ME2 ;
  RECT 32.556 0.000 32.876 0.600 ;
  LAYER ME1 ;
  RECT 32.556 0.000 32.876 0.600 ;
 END
 ANTENNAPARTIALMETALAREA                  1.910 LAYER ME2 ;
 ANTENNAGATEAREA                          0.180 LAYER ME2 ;
 ANTENNAGATEAREA                          0.180 LAYER ME3 ;
 ANTENNAGATEAREA                          0.180 LAYER ME4 ;
 ANTENNADIFFAREA                          0.218 LAYER ME2 ;
 ANTENNADIFFAREA                          0.218 LAYER ME3 ;
 ANTENNADIFFAREA                          0.218 LAYER ME4 ;
 ANTENNAMAXAREACAR                       13.456 LAYER ME2 ;
 ANTENNAMAXAREACAR                       14.522 LAYER ME3 ;
 ANTENNAMAXAREACAR                       15.589 LAYER ME4 ;
END A6
PIN A1
  DIRECTION INPUT ;
 PORT
  LAYER ME3 ;
  RECT 47.781 0.000 48.101 0.712 ;
  LAYER ME2 ;
  RECT 47.781 0.000 48.101 0.712 ;
  LAYER ME1 ;
  RECT 47.781 0.000 48.101 0.712 ;
 END
 ANTENNAPARTIALMETALAREA                  3.219 LAYER ME2 ;
 ANTENNAGATEAREA                          0.108 LAYER ME2 ;
 ANTENNAGATEAREA                          0.108 LAYER ME3 ;
 ANTENNADIFFAREA                          0.218 LAYER ME2 ;
 ANTENNADIFFAREA                          0.218 LAYER ME3 ;
 ANTENNAMAXAREACAR                       33.245 LAYER ME2 ;
 ANTENNAMAXAREACAR                       35.355 LAYER ME3 ;
END A1
PIN A0
  DIRECTION INPUT ;
 PORT
  LAYER ME3 ;
  RECT 51.010 0.000 51.330 0.712 ;
  LAYER ME2 ;
  RECT 51.010 0.000 51.330 0.712 ;
  LAYER ME1 ;
  RECT 51.010 0.000 51.330 0.712 ;
 END
 ANTENNAPARTIALMETALAREA                  3.457 LAYER ME2 ;
 ANTENNAGATEAREA                          0.108 LAYER ME2 ;
 ANTENNAGATEAREA                          0.108 LAYER ME3 ;
 ANTENNADIFFAREA                          0.218 LAYER ME2 ;
 ANTENNADIFFAREA                          0.218 LAYER ME3 ;
 ANTENNAMAXAREACAR                       35.986 LAYER ME2 ;
 ANTENNAMAXAREACAR                       38.095 LAYER ME3 ;
END A0
PIN DVSE
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 63.601 0.000 63.921 0.717 ;
  LAYER ME3 ;
  RECT 63.601 0.000 63.921 0.717 ;
  LAYER ME3 ;
  RECT 63.601 0.000 63.921 0.717 ;
  LAYER ME2 ;
  RECT 63.601 0.000 63.921 0.717 ;
  LAYER ME2 ;
  RECT 63.601 0.000 63.921 0.717 ;
  LAYER ME1 ;
  RECT 63.601 0.000 63.921 0.717 ;
  LAYER ME1 ;
  RECT 63.601 0.000 63.921 0.717 ;
 END
 ANTENNAPARTIALMETALAREA                  5.305 LAYER ME2 ;
 ANTENNAGATEAREA                          0.612 LAYER ME2 ;
 ANTENNAGATEAREA                          0.612 LAYER ME3 ;
 ANTENNAGATEAREA                          0.612 LAYER ME4 ;
 ANTENNADIFFAREA                          0.218 LAYER ME2 ;
 ANTENNADIFFAREA                          0.218 LAYER ME3 ;
 ANTENNADIFFAREA                          0.218 LAYER ME4 ;
 ANTENNAMAXAREACAR                       53.132 LAYER ME2 ;
 ANTENNAMAXAREACAR                       55.256 LAYER ME3 ;
 ANTENNAMAXAREACAR                       57.381 LAYER ME4 ;
END DVSE
PIN DVS3
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 63.081 0.000 63.401 0.717 ;
  LAYER ME3 ;
  RECT 63.081 0.000 63.401 0.717 ;
  LAYER ME3 ;
  RECT 63.081 0.000 63.401 0.717 ;
  LAYER ME2 ;
  RECT 63.081 0.000 63.401 0.717 ;
  LAYER ME2 ;
  RECT 63.081 0.000 63.401 0.717 ;
  LAYER ME1 ;
  RECT 63.081 0.000 63.401 0.717 ;
  LAYER ME1 ;
  RECT 63.081 0.000 63.401 0.717 ;
 END
 ANTENNAPARTIALMETALAREA                  3.675 LAYER ME2 ;
 ANTENNAGATEAREA                          0.108 LAYER ME2 ;
 ANTENNAGATEAREA                          0.108 LAYER ME3 ;
 ANTENNAGATEAREA                          0.108 LAYER ME4 ;
 ANTENNADIFFAREA                          0.218 LAYER ME2 ;
 ANTENNADIFFAREA                          0.218 LAYER ME3 ;
 ANTENNADIFFAREA                          0.218 LAYER ME4 ;
 ANTENNAMAXAREACAR                       45.625 LAYER ME2 ;
 ANTENNAMAXAREACAR                       47.749 LAYER ME3 ;
 ANTENNAMAXAREACAR                       49.874 LAYER ME4 ;
END DVS3
PIN DVS2
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 64.121 0.000 64.441 0.717 ;
  LAYER ME3 ;
  RECT 64.121 0.000 64.441 0.717 ;
  LAYER ME3 ;
  RECT 64.121 0.000 64.441 0.717 ;
  LAYER ME2 ;
  RECT 64.121 0.000 64.441 0.717 ;
  LAYER ME2 ;
  RECT 64.121 0.000 64.441 0.717 ;
  LAYER ME1 ;
  RECT 64.121 0.000 64.441 0.717 ;
  LAYER ME1 ;
  RECT 64.121 0.000 64.441 0.717 ;
 END
 ANTENNAPARTIALMETALAREA                  5.371 LAYER ME2 ;
 ANTENNAGATEAREA                          0.108 LAYER ME2 ;
 ANTENNAGATEAREA                          0.108 LAYER ME3 ;
 ANTENNAGATEAREA                          0.108 LAYER ME4 ;
 ANTENNADIFFAREA                          0.218 LAYER ME2 ;
 ANTENNADIFFAREA                          0.218 LAYER ME3 ;
 ANTENNADIFFAREA                          0.218 LAYER ME4 ;
 ANTENNAMAXAREACAR                       60.060 LAYER ME2 ;
 ANTENNAMAXAREACAR                       62.184 LAYER ME3 ;
 ANTENNAMAXAREACAR                       64.309 LAYER ME4 ;
END DVS2
PIN DVS1
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 62.561 0.000 62.881 0.717 ;
  LAYER ME3 ;
  RECT 62.561 0.000 62.881 0.717 ;
  LAYER ME3 ;
  RECT 62.561 0.000 62.881 0.717 ;
  LAYER ME2 ;
  RECT 62.561 0.000 62.881 0.717 ;
  LAYER ME2 ;
  RECT 62.561 0.000 62.881 0.717 ;
  LAYER ME1 ;
  RECT 62.561 0.000 62.881 0.717 ;
  LAYER ME1 ;
  RECT 62.561 0.000 62.881 0.717 ;
 END
 ANTENNAPARTIALMETALAREA                  3.307 LAYER ME2 ;
 ANTENNAGATEAREA                          0.108 LAYER ME2 ;
 ANTENNAGATEAREA                          0.108 LAYER ME3 ;
 ANTENNAGATEAREA                          0.108 LAYER ME4 ;
 ANTENNADIFFAREA                          0.218 LAYER ME2 ;
 ANTENNADIFFAREA                          0.218 LAYER ME3 ;
 ANTENNADIFFAREA                          0.218 LAYER ME4 ;
 ANTENNAMAXAREACAR                       42.063 LAYER ME2 ;
 ANTENNAMAXAREACAR                       44.188 LAYER ME3 ;
 ANTENNAMAXAREACAR                       46.312 LAYER ME4 ;
END DVS1
PIN DVS0
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 64.641 0.000 64.961 0.693 ;
  LAYER ME3 ;
  RECT 64.641 0.000 64.961 0.693 ;
  LAYER ME3 ;
  RECT 64.641 0.000 64.961 0.693 ;
  LAYER ME2 ;
  RECT 64.641 0.000 64.961 0.693 ;
  LAYER ME2 ;
  RECT 64.641 0.000 64.961 0.693 ;
  LAYER ME1 ;
  RECT 64.641 0.000 64.961 0.693 ;
  LAYER ME1 ;
  RECT 64.641 0.000 64.961 0.693 ;
 END
 ANTENNAPARTIALMETALAREA                  4.376 LAYER ME2 ;
 ANTENNAGATEAREA                          0.108 LAYER ME2 ;
 ANTENNAGATEAREA                          0.108 LAYER ME3 ;
 ANTENNAGATEAREA                          0.108 LAYER ME4 ;
 ANTENNADIFFAREA                          0.218 LAYER ME2 ;
 ANTENNADIFFAREA                          0.218 LAYER ME3 ;
 ANTENNADIFFAREA                          0.218 LAYER ME4 ;
 ANTENNAMAXAREACAR                       53.260 LAYER ME2 ;
 ANTENNAMAXAREACAR                       55.313 LAYER ME3 ;
 ANTENNAMAXAREACAR                       57.367 LAYER ME4 ;
END DVS0
PIN CK
  DIRECTION INPUT ;
 PORT
  LAYER ME3 ;
  RECT 56.077 0.000 56.397 0.713 ;
  LAYER ME2 ;
  RECT 56.077 0.000 56.397 0.713 ;
  LAYER ME1 ;
  RECT 56.077 0.000 56.397 0.713 ;
 END
 ANTENNAPARTIALMETALAREA                  2.392 LAYER ME2 ;
 ANTENNAPARTIALMETALAREA                  7.363 LAYER ME3 ;
 ANTENNAGATEAREA                          0.072 LAYER ME2 ;
 ANTENNAGATEAREA                          1.260 LAYER ME3 ;
 ANTENNADIFFAREA                          0.218 LAYER ME2 ;
 ANTENNADIFFAREA                          0.218 LAYER ME3 ;
 ANTENNAMAXAREACAR                       46.148 LAYER ME2 ;
 ANTENNAMAXAREACAR                      151.587 LAYER ME3 ;
END CK
PIN CSB
  DIRECTION INPUT ;
 PORT
  LAYER ME3 ;
  RECT 49.289 0.000 49.609 0.712 ;
  LAYER ME2 ;
  RECT 49.289 0.000 49.609 0.712 ;
  LAYER ME1 ;
  RECT 49.289 0.000 49.609 0.712 ;
 END
 ANTENNAPARTIALMETALAREA                  3.350 LAYER ME2 ;
 ANTENNAPARTIALMETALAREA                  7.235 LAYER ME3 ;
 ANTENNAGATEAREA                          2.244 LAYER ME2 ;
 ANTENNAGATEAREA                          3.216 LAYER ME3 ;
 ANTENNADIFFAREA                          0.218 LAYER ME2 ;
 ANTENNADIFFAREA                          0.218 LAYER ME3 ;
 ANTENNAMAXAREACAR                       17.231 LAYER ME2 ;
 ANTENNAMAXAREACAR                       51.784 LAYER ME3 ;
END CSB
PIN WEB
  DIRECTION INPUT ;
 PORT
  LAYER ME3 ;
  RECT 59.788 0.000 60.108 0.717 ;
  LAYER ME2 ;
  RECT 59.788 0.000 60.108 0.717 ;
  LAYER ME1 ;
  RECT 59.788 0.000 60.108 0.717 ;
 END
 ANTENNAPARTIALMETALAREA                  0.681 LAYER ME2 ;
 ANTENNAPARTIALMETALAREA                 10.739 LAYER ME3 ;
 ANTENNAGATEAREA                          0.576 LAYER ME3 ;
 ANTENNADIFFAREA                          0.218 LAYER ME2 ;
 ANTENNADIFFAREA                          0.653 LAYER ME3 ;
 ANTENNAMAXAREACAR                       41.333 LAYER ME3 ;
END WEB
PIN DI6
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 94.331 0.000 94.611 0.720 ;
  LAYER ME3 ;
  RECT 94.331 0.000 94.611 0.720 ;
  LAYER ME2 ;
  RECT 94.331 0.000 94.611 0.720 ;
  LAYER ME1 ;
  RECT 94.331 0.000 94.611 0.720 ;
 END
 ANTENNAPARTIALMETALAREA                  0.805 LAYER ME1 ;
 ANTENNAGATEAREA                          0.072 LAYER ME1 ;
 ANTENNAGATEAREA                          0.072 LAYER ME2 ;
 ANTENNAGATEAREA                          0.072 LAYER ME3 ;
 ANTENNAGATEAREA                          0.072 LAYER ME4 ;
 ANTENNADIFFAREA                          0.218 LAYER ME1 ;
 ANTENNADIFFAREA                          0.218 LAYER ME2 ;
 ANTENNADIFFAREA                          0.218 LAYER ME3 ;
 ANTENNADIFFAREA                          0.218 LAYER ME4 ;
 ANTENNAMAXAREACAR                       13.984 LAYER ME1 ;
 ANTENNAMAXAREACAR                       16.784 LAYER ME2 ;
 ANTENNAMAXAREACAR                       19.584 LAYER ME3 ;
 ANTENNAMAXAREACAR                       22.384 LAYER ME4 ;
END DI6
PIN DO6
  DIRECTION OUTPUT ;
 PORT
  LAYER ME4 ;
  RECT 92.353 0.000 92.633 0.720 ;
  LAYER ME3 ;
  RECT 92.353 0.000 92.633 0.720 ;
  LAYER ME2 ;
  RECT 92.353 0.000 92.633 0.720 ;
  LAYER ME1 ;
  RECT 92.353 0.000 92.633 0.720 ;
 END
 ANTENNAPARTIALMETALAREA                  2.030 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME3 ;
 ANTENNADIFFAREA                          1.293 LAYER ME4 ;
END DO6
PIN DI5
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 86.323 0.000 86.603 0.720 ;
  LAYER ME3 ;
  RECT 86.323 0.000 86.603 0.720 ;
  LAYER ME2 ;
  RECT 86.323 0.000 86.603 0.720 ;
  LAYER ME1 ;
  RECT 86.323 0.000 86.603 0.720 ;
 END
 ANTENNAPARTIALMETALAREA                  0.805 LAYER ME1 ;
 ANTENNAGATEAREA                          0.072 LAYER ME1 ;
 ANTENNAGATEAREA                          0.072 LAYER ME2 ;
 ANTENNAGATEAREA                          0.072 LAYER ME3 ;
 ANTENNAGATEAREA                          0.072 LAYER ME4 ;
 ANTENNADIFFAREA                          0.218 LAYER ME1 ;
 ANTENNADIFFAREA                          0.218 LAYER ME2 ;
 ANTENNADIFFAREA                          0.218 LAYER ME3 ;
 ANTENNADIFFAREA                          0.218 LAYER ME4 ;
 ANTENNAMAXAREACAR                       13.984 LAYER ME1 ;
 ANTENNAMAXAREACAR                       16.784 LAYER ME2 ;
 ANTENNAMAXAREACAR                       19.584 LAYER ME3 ;
 ANTENNAMAXAREACAR                       22.384 LAYER ME4 ;
END DI5
PIN DO5
  DIRECTION OUTPUT ;
 PORT
  LAYER ME4 ;
  RECT 84.345 0.000 84.625 0.720 ;
  LAYER ME3 ;
  RECT 84.345 0.000 84.625 0.720 ;
  LAYER ME2 ;
  RECT 84.345 0.000 84.625 0.720 ;
  LAYER ME1 ;
  RECT 84.345 0.000 84.625 0.720 ;
 END
 ANTENNAPARTIALMETALAREA                  2.030 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME3 ;
 ANTENNADIFFAREA                          1.293 LAYER ME4 ;
END DO5
PIN DI4
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 78.315 0.000 78.595 0.720 ;
  LAYER ME3 ;
  RECT 78.315 0.000 78.595 0.720 ;
  LAYER ME2 ;
  RECT 78.315 0.000 78.595 0.720 ;
  LAYER ME1 ;
  RECT 78.315 0.000 78.595 0.720 ;
 END
 ANTENNAPARTIALMETALAREA                  0.805 LAYER ME1 ;
 ANTENNAGATEAREA                          0.072 LAYER ME1 ;
 ANTENNAGATEAREA                          0.072 LAYER ME2 ;
 ANTENNAGATEAREA                          0.072 LAYER ME3 ;
 ANTENNAGATEAREA                          0.072 LAYER ME4 ;
 ANTENNADIFFAREA                          0.218 LAYER ME1 ;
 ANTENNADIFFAREA                          0.218 LAYER ME2 ;
 ANTENNADIFFAREA                          0.218 LAYER ME3 ;
 ANTENNADIFFAREA                          0.218 LAYER ME4 ;
 ANTENNAMAXAREACAR                       13.984 LAYER ME1 ;
 ANTENNAMAXAREACAR                       16.784 LAYER ME2 ;
 ANTENNAMAXAREACAR                       19.584 LAYER ME3 ;
 ANTENNAMAXAREACAR                       22.384 LAYER ME4 ;
END DI4
PIN DO4
  DIRECTION OUTPUT ;
 PORT
  LAYER ME4 ;
  RECT 76.337 0.000 76.617 0.720 ;
  LAYER ME3 ;
  RECT 76.337 0.000 76.617 0.720 ;
  LAYER ME2 ;
  RECT 76.337 0.000 76.617 0.720 ;
  LAYER ME1 ;
  RECT 76.337 0.000 76.617 0.720 ;
 END
 ANTENNAPARTIALMETALAREA                  2.030 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME3 ;
 ANTENNADIFFAREA                          1.293 LAYER ME4 ;
END DO4
PIN DI3
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 70.307 0.000 70.587 0.720 ;
  LAYER ME3 ;
  RECT 70.307 0.000 70.587 0.720 ;
  LAYER ME2 ;
  RECT 70.307 0.000 70.587 0.720 ;
  LAYER ME1 ;
  RECT 70.307 0.000 70.587 0.720 ;
 END
 ANTENNAPARTIALMETALAREA                  0.522 LAYER ME1 ;
 ANTENNAGATEAREA                          0.072 LAYER ME1 ;
 ANTENNAGATEAREA                          0.072 LAYER ME2 ;
 ANTENNAGATEAREA                          0.072 LAYER ME3 ;
 ANTENNAGATEAREA                          0.072 LAYER ME4 ;
 ANTENNADIFFAREA                          0.218 LAYER ME1 ;
 ANTENNADIFFAREA                          0.218 LAYER ME2 ;
 ANTENNADIFFAREA                          0.218 LAYER ME3 ;
 ANTENNADIFFAREA                          0.218 LAYER ME4 ;
 ANTENNAMAXAREACAR                       10.048 LAYER ME1 ;
 ANTENNAMAXAREACAR                       12.848 LAYER ME2 ;
 ANTENNAMAXAREACAR                       15.648 LAYER ME3 ;
 ANTENNAMAXAREACAR                       18.448 LAYER ME4 ;
END DI3
PIN DO3
  DIRECTION OUTPUT ;
 PORT
  LAYER ME4 ;
  RECT 68.249 0.000 68.529 0.720 ;
  LAYER ME3 ;
  RECT 68.249 0.000 68.529 0.720 ;
  LAYER ME2 ;
  RECT 68.249 0.000 68.529 0.720 ;
  LAYER ME1 ;
  RECT 68.249 0.000 68.529 0.720 ;
 END
 ANTENNAPARTIALMETALAREA                  2.030 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME3 ;
 ANTENNADIFFAREA                          1.293 LAYER ME4 ;
END DO3
OBS
  LAYER ME3 ;
  RECT 0.000 0.000 99.555 68.179 ;
  LAYER ME2 ;
  RECT 0.000 0.000 99.555 68.179 ;
  LAYER ME1 ;
  RECT 0.000 0.000 99.555 68.179 ;
  LAYER ME4 ;
  RECT 0.000 0.000 39.766 68.179 ;
  LAYER ME4 ;
  RECT 41.420 0.000 42.540 68.179 ;
  LAYER ME4 ;
  RECT 44.135 0.000 44.855 68.179 ;
  LAYER ME4 ;
  RECT 45.585 0.000 46.305 68.179 ;
  LAYER ME4 ;
  RECT 48.365 0.000 48.965 68.179 ;
  LAYER ME4 ;
  RECT 51.579 0.000 53.265 68.179 ;
  LAYER ME4 ;
  RECT 54.655 0.000 55.775 68.179 ;
  LAYER ME4 ;
  RECT 57.050 0.000 57.770 68.179 ;
  LAYER ME4 ;
  RECT 58.765 0.000 59.485 68.179 ;
  LAYER ME4 ;
  RECT 60.685 0.000 99.555 68.179 ;
END
END SYKB110_128X7X1CM4
END LIBRARY





