# ________________________________________________________________________________________________
# 
# 
#             Synchronous One-Port Register File Compiler
# 
#                 UMC 0.11um LL AE Logic Process
# 
# ________________________________________________________________________________________________
# 
#               
#         Copyright (C) 2024 Faraday Technology Corporation. All Rights Reserved.       
#                
#         This source code is an unpublished work belongs to Faraday Technology Corporation       
#         It is considered a trade secret and is not to be divulged or       
#         used by parties who have not received written authorization from       
#         Faraday Technology Corporation       
#                
#         Faraday's home page can be found at: http://www.faraday-tech.com/       
#                
# ________________________________________________________________________________________________
# 
#        IP Name            :  FSR0K_B_SY                
#        IP Version         :  1.4.0                     
#        IP Release Status  :  Active                    
#        Word               :  128                       
#        Bit                :  7                         
#        Byte               :  6                         
#        Mux                :  4                         
#        Output Loading     :  0.01                      
#        Clock Input Slew   :  0.016                     
#        Data Input Slew    :  0.016                     
#        Ring Type          :  Ringless Model            
#        Ring Width         :  0                         
#        Bus Format         :  0                         
#        Memaker Path       :  /home/mem/Desktop/memlib  
#        GUI Version        :  m20230904                 
#        Date               :  2024/09/06 19:52:02       
# ________________________________________________________________________________________________
# 

VERSION 5.5 ;
NAMESCASESENSITIVE ON ;
MACRO SYKB110_128X7X6CM4
CLASS BLOCK ;
FOREIGN SYKB110_128X7X6CM4 0.000 0.000 ;
ORIGIN 0.000 0.000 ;
SIZE 379.835 BY 68.179 ;
SYMMETRY x y r90 ;
SITE core ;
PIN VCC
  DIRECTION INOUT ;
  USE POWER ;
 PORT
  LAYER ME4 ;
  RECT 213.401 0.000 214.121 33.870 ;
 END
 PORT
  LAYER ME4 ;
  RECT 209.397 0.000 210.117 33.870 ;
 END
 PORT
  LAYER ME4 ;
  RECT 221.409 0.000 222.129 33.870 ;
 END
 PORT
  LAYER ME4 ;
  RECT 217.405 0.000 218.125 33.870 ;
 END
 PORT
  LAYER ME4 ;
  RECT 229.417 0.000 230.137 33.870 ;
 END
 PORT
  LAYER ME4 ;
  RECT 225.413 0.000 226.133 33.870 ;
 END
 PORT
  LAYER ME4 ;
  RECT 237.425 0.000 238.145 33.870 ;
 END
 PORT
  LAYER ME4 ;
  RECT 233.421 0.000 234.141 33.870 ;
 END
 PORT
  LAYER ME4 ;
  RECT 245.433 0.000 246.153 33.870 ;
 END
 PORT
  LAYER ME4 ;
  RECT 241.429 0.000 242.149 33.870 ;
 END
 PORT
  LAYER ME4 ;
  RECT 253.441 0.000 254.161 33.870 ;
 END
 PORT
  LAYER ME4 ;
  RECT 249.437 0.000 250.157 33.870 ;
 END
 PORT
  LAYER ME4 ;
  RECT 261.449 0.000 262.169 33.870 ;
 END
 PORT
  LAYER ME4 ;
  RECT 257.445 0.000 258.165 33.870 ;
 END
 PORT
  LAYER ME4 ;
  RECT 269.457 0.000 270.177 33.870 ;
 END
 PORT
  LAYER ME4 ;
  RECT 265.453 0.000 266.173 33.870 ;
 END
 PORT
  LAYER ME4 ;
  RECT 277.465 0.000 278.185 33.870 ;
 END
 PORT
  LAYER ME4 ;
  RECT 273.461 0.000 274.181 33.870 ;
 END
 PORT
  LAYER ME4 ;
  RECT 285.473 0.000 286.193 33.870 ;
 END
 PORT
  LAYER ME4 ;
  RECT 281.469 0.000 282.189 33.870 ;
 END
 PORT
  LAYER ME4 ;
  RECT 293.481 0.000 294.201 33.870 ;
 END
 PORT
  LAYER ME4 ;
  RECT 289.477 0.000 290.197 33.870 ;
 END
 PORT
  LAYER ME4 ;
  RECT 301.489 0.000 302.209 33.870 ;
 END
 PORT
  LAYER ME4 ;
  RECT 297.485 0.000 298.205 33.870 ;
 END
 PORT
  LAYER ME4 ;
  RECT 309.497 0.000 310.217 33.870 ;
 END
 PORT
  LAYER ME4 ;
  RECT 305.493 0.000 306.213 33.870 ;
 END
 PORT
  LAYER ME4 ;
  RECT 317.505 0.000 318.225 33.870 ;
 END
 PORT
  LAYER ME4 ;
  RECT 313.501 0.000 314.221 33.870 ;
 END
 PORT
  LAYER ME4 ;
  RECT 325.513 0.000 326.233 33.870 ;
 END
 PORT
  LAYER ME4 ;
  RECT 321.509 0.000 322.229 33.870 ;
 END
 PORT
  LAYER ME4 ;
  RECT 333.521 0.000 334.241 33.870 ;
 END
 PORT
  LAYER ME4 ;
  RECT 329.517 0.000 330.237 33.870 ;
 END
 PORT
  LAYER ME4 ;
  RECT 341.529 0.000 342.249 33.870 ;
 END
 PORT
  LAYER ME4 ;
  RECT 337.525 0.000 338.245 33.870 ;
 END
 PORT
  LAYER ME4 ;
  RECT 349.537 0.000 350.257 33.870 ;
 END
 PORT
  LAYER ME4 ;
  RECT 345.533 0.000 346.253 33.870 ;
 END
 PORT
  LAYER ME4 ;
  RECT 357.545 0.000 358.265 33.870 ;
 END
 PORT
  LAYER ME4 ;
  RECT 353.541 0.000 354.261 33.870 ;
 END
 PORT
  LAYER ME4 ;
  RECT 365.553 0.000 366.273 33.870 ;
 END
 PORT
  LAYER ME4 ;
  RECT 361.549 0.000 362.269 33.870 ;
 END
 PORT
  LAYER ME4 ;
  RECT 373.561 0.000 374.281 33.870 ;
 END
 PORT
  LAYER ME4 ;
  RECT 369.557 0.000 370.277 33.870 ;
 END
 PORT
  LAYER ME4 ;
  RECT 378.535 0.000 378.915 68.179 ;
 END
 PORT
  LAYER ME4 ;
  RECT 192.509 0.000 193.109 68.179 ;
 END
 PORT
  LAYER ME4 ;
  RECT 196.689 0.000 197.409 68.179 ;
 END
 PORT
  LAYER ME4 ;
  RECT 198.799 0.000 199.919 68.179 ;
 END
 PORT
  LAYER ME4 ;
  RECT 204.829 0.000 205.549 68.179 ;
 END
 PORT
  LAYER ME4 ;
  RECT 206.765 0.921 207.145 68.179 ;
 END
 PORT
  LAYER ME4 ;
  RECT 185.564 0.000 186.684 68.179 ;
 END
 PORT
  LAYER ME4 ;
  RECT 188.279 0.000 188.999 68.179 ;
 END
 PORT
  LAYER ME4 ;
  RECT 183.190 0.000 183.910 67.420 ;
 END
 PORT
  LAYER ME4 ;
  RECT 181.150 0.921 181.870 68.179 ;
 END
 PORT
  LAYER ME4 ;
  RECT 179.030 0.000 179.750 68.179 ;
 END
 PORT
  LAYER ME4 ;
  RECT 176.990 0.921 177.710 68.179 ;
 END
 PORT
  LAYER ME4 ;
  RECT 0.920 0.000 1.300 68.179 ;
 END
 PORT
  LAYER ME4 ;
  RECT 7.556 0.000 8.276 33.870 ;
 END
 PORT
  LAYER ME4 ;
  RECT 3.552 0.000 4.272 33.870 ;
 END
 PORT
  LAYER ME4 ;
  RECT 15.564 0.000 16.284 33.870 ;
 END
 PORT
  LAYER ME4 ;
  RECT 11.560 0.000 12.280 33.870 ;
 END
 PORT
  LAYER ME4 ;
  RECT 23.572 0.000 24.292 33.870 ;
 END
 PORT
  LAYER ME4 ;
  RECT 19.568 0.000 20.288 33.870 ;
 END
 PORT
  LAYER ME4 ;
  RECT 31.580 0.000 32.300 33.870 ;
 END
 PORT
  LAYER ME4 ;
  RECT 27.576 0.000 28.296 33.870 ;
 END
 PORT
  LAYER ME4 ;
  RECT 39.588 0.000 40.308 33.870 ;
 END
 PORT
  LAYER ME4 ;
  RECT 35.584 0.000 36.304 33.870 ;
 END
 PORT
  LAYER ME4 ;
  RECT 47.596 0.000 48.316 33.870 ;
 END
 PORT
  LAYER ME4 ;
  RECT 43.592 0.000 44.312 33.870 ;
 END
 PORT
  LAYER ME4 ;
  RECT 55.604 0.000 56.324 33.870 ;
 END
 PORT
  LAYER ME4 ;
  RECT 51.600 0.000 52.320 33.870 ;
 END
 PORT
  LAYER ME4 ;
  RECT 63.612 0.000 64.332 33.870 ;
 END
 PORT
  LAYER ME4 ;
  RECT 59.608 0.000 60.328 33.870 ;
 END
 PORT
  LAYER ME4 ;
  RECT 71.620 0.000 72.340 33.870 ;
 END
 PORT
  LAYER ME4 ;
  RECT 67.616 0.000 68.336 33.870 ;
 END
 PORT
  LAYER ME4 ;
  RECT 79.628 0.000 80.348 33.870 ;
 END
 PORT
  LAYER ME4 ;
  RECT 75.624 0.000 76.344 33.870 ;
 END
 PORT
  LAYER ME4 ;
  RECT 87.636 0.000 88.356 33.870 ;
 END
 PORT
  LAYER ME4 ;
  RECT 83.632 0.000 84.352 33.870 ;
 END
 PORT
  LAYER ME4 ;
  RECT 95.644 0.000 96.364 33.870 ;
 END
 PORT
  LAYER ME4 ;
  RECT 91.640 0.000 92.360 33.870 ;
 END
 PORT
  LAYER ME4 ;
  RECT 103.652 0.000 104.372 33.870 ;
 END
 PORT
  LAYER ME4 ;
  RECT 99.648 0.000 100.368 33.870 ;
 END
 PORT
  LAYER ME4 ;
  RECT 111.660 0.000 112.380 33.870 ;
 END
 PORT
  LAYER ME4 ;
  RECT 107.656 0.000 108.376 33.870 ;
 END
 PORT
  LAYER ME4 ;
  RECT 119.668 0.000 120.388 33.870 ;
 END
 PORT
  LAYER ME4 ;
  RECT 115.664 0.000 116.384 33.870 ;
 END
 PORT
  LAYER ME4 ;
  RECT 127.676 0.000 128.396 33.870 ;
 END
 PORT
  LAYER ME4 ;
  RECT 123.672 0.000 124.392 33.870 ;
 END
 PORT
  LAYER ME4 ;
  RECT 135.684 0.000 136.404 33.870 ;
 END
 PORT
  LAYER ME4 ;
  RECT 131.680 0.000 132.400 33.870 ;
 END
 PORT
  LAYER ME4 ;
  RECT 143.692 0.000 144.412 33.870 ;
 END
 PORT
  LAYER ME4 ;
  RECT 139.688 0.000 140.408 33.870 ;
 END
 PORT
  LAYER ME4 ;
  RECT 151.700 0.000 152.420 33.870 ;
 END
 PORT
  LAYER ME4 ;
  RECT 147.696 0.000 148.416 33.870 ;
 END
 PORT
  LAYER ME4 ;
  RECT 159.708 0.000 160.428 33.870 ;
 END
 PORT
  LAYER ME4 ;
  RECT 155.704 0.000 156.424 33.870 ;
 END
 PORT
  LAYER ME4 ;
  RECT 167.716 0.000 168.436 33.870 ;
 END
 PORT
  LAYER ME4 ;
  RECT 163.712 0.000 164.432 33.870 ;
 END
 PORT
  LAYER ME4 ;
  RECT 174.870 0.000 175.590 68.179 ;
 END
 PORT
  LAYER ME4 ;
  RECT 172.690 0.000 173.070 68.179 ;
 END
 PORT
  LAYER ME4 ;
  RECT 215.593 35.220 215.933 68.179 ;
 END
 PORT
  LAYER ME4 ;
  RECT 213.591 35.220 213.931 68.179 ;
 END
 PORT
  LAYER ME4 ;
  RECT 211.589 35.220 211.929 68.179 ;
 END
 PORT
  LAYER ME4 ;
  RECT 209.587 35.220 209.927 68.179 ;
 END
 PORT
  LAYER ME4 ;
  RECT 223.601 35.220 223.941 68.179 ;
 END
 PORT
  LAYER ME4 ;
  RECT 221.599 35.220 221.939 68.179 ;
 END
 PORT
  LAYER ME4 ;
  RECT 219.597 35.220 219.937 68.179 ;
 END
 PORT
  LAYER ME4 ;
  RECT 217.595 35.220 217.935 68.179 ;
 END
 PORT
  LAYER ME4 ;
  RECT 231.609 35.220 231.949 68.179 ;
 END
 PORT
  LAYER ME4 ;
  RECT 229.607 35.220 229.947 68.179 ;
 END
 PORT
  LAYER ME4 ;
  RECT 227.605 35.220 227.945 68.179 ;
 END
 PORT
  LAYER ME4 ;
  RECT 225.603 35.220 225.943 68.179 ;
 END
 PORT
  LAYER ME4 ;
  RECT 239.617 35.220 239.957 68.179 ;
 END
 PORT
  LAYER ME4 ;
  RECT 237.615 35.220 237.955 68.179 ;
 END
 PORT
  LAYER ME4 ;
  RECT 235.613 35.220 235.953 68.179 ;
 END
 PORT
  LAYER ME4 ;
  RECT 233.611 35.220 233.951 68.179 ;
 END
 PORT
  LAYER ME4 ;
  RECT 247.625 35.220 247.965 68.179 ;
 END
 PORT
  LAYER ME4 ;
  RECT 245.623 35.220 245.963 68.179 ;
 END
 PORT
  LAYER ME4 ;
  RECT 243.621 35.220 243.961 68.179 ;
 END
 PORT
  LAYER ME4 ;
  RECT 241.619 35.220 241.959 68.179 ;
 END
 PORT
  LAYER ME4 ;
  RECT 255.633 35.220 255.973 68.179 ;
 END
 PORT
  LAYER ME4 ;
  RECT 253.631 35.220 253.971 68.179 ;
 END
 PORT
  LAYER ME4 ;
  RECT 251.629 35.220 251.969 68.179 ;
 END
 PORT
  LAYER ME4 ;
  RECT 249.627 35.220 249.967 68.179 ;
 END
 PORT
  LAYER ME4 ;
  RECT 263.641 35.220 263.981 68.179 ;
 END
 PORT
  LAYER ME4 ;
  RECT 261.639 35.220 261.979 68.179 ;
 END
 PORT
  LAYER ME4 ;
  RECT 259.637 35.220 259.977 68.179 ;
 END
 PORT
  LAYER ME4 ;
  RECT 257.635 35.220 257.975 68.179 ;
 END
 PORT
  LAYER ME4 ;
  RECT 271.649 35.220 271.989 68.179 ;
 END
 PORT
  LAYER ME4 ;
  RECT 269.647 35.220 269.987 68.179 ;
 END
 PORT
  LAYER ME4 ;
  RECT 267.645 35.220 267.985 68.179 ;
 END
 PORT
  LAYER ME4 ;
  RECT 265.643 35.220 265.983 68.179 ;
 END
 PORT
  LAYER ME4 ;
  RECT 279.657 35.220 279.997 68.179 ;
 END
 PORT
  LAYER ME4 ;
  RECT 277.655 35.220 277.995 68.179 ;
 END
 PORT
  LAYER ME4 ;
  RECT 275.653 35.220 275.993 68.179 ;
 END
 PORT
  LAYER ME4 ;
  RECT 273.651 35.220 273.991 68.179 ;
 END
 PORT
  LAYER ME4 ;
  RECT 287.665 35.220 288.005 68.179 ;
 END
 PORT
  LAYER ME4 ;
  RECT 285.663 35.220 286.003 68.179 ;
 END
 PORT
  LAYER ME4 ;
  RECT 283.661 35.220 284.001 68.179 ;
 END
 PORT
  LAYER ME4 ;
  RECT 281.659 35.220 281.999 68.179 ;
 END
 PORT
  LAYER ME4 ;
  RECT 295.673 35.220 296.013 68.179 ;
 END
 PORT
  LAYER ME4 ;
  RECT 293.671 35.220 294.011 68.179 ;
 END
 PORT
  LAYER ME4 ;
  RECT 291.669 35.220 292.009 68.179 ;
 END
 PORT
  LAYER ME4 ;
  RECT 289.667 35.220 290.007 68.179 ;
 END
 PORT
  LAYER ME4 ;
  RECT 303.681 35.220 304.021 68.179 ;
 END
 PORT
  LAYER ME4 ;
  RECT 301.679 35.220 302.019 68.179 ;
 END
 PORT
  LAYER ME4 ;
  RECT 299.677 35.220 300.017 68.179 ;
 END
 PORT
  LAYER ME4 ;
  RECT 297.675 35.220 298.015 68.179 ;
 END
 PORT
  LAYER ME4 ;
  RECT 311.689 35.220 312.029 68.179 ;
 END
 PORT
  LAYER ME4 ;
  RECT 309.687 35.220 310.027 68.179 ;
 END
 PORT
  LAYER ME4 ;
  RECT 307.685 35.220 308.025 68.179 ;
 END
 PORT
  LAYER ME4 ;
  RECT 305.683 35.220 306.023 68.179 ;
 END
 PORT
  LAYER ME4 ;
  RECT 319.697 35.220 320.037 68.179 ;
 END
 PORT
  LAYER ME4 ;
  RECT 317.695 35.220 318.035 68.179 ;
 END
 PORT
  LAYER ME4 ;
  RECT 315.693 35.220 316.033 68.179 ;
 END
 PORT
  LAYER ME4 ;
  RECT 313.691 35.220 314.031 68.179 ;
 END
 PORT
  LAYER ME4 ;
  RECT 327.705 35.220 328.045 68.179 ;
 END
 PORT
  LAYER ME4 ;
  RECT 325.703 35.220 326.043 68.179 ;
 END
 PORT
  LAYER ME4 ;
  RECT 323.701 35.220 324.041 68.179 ;
 END
 PORT
  LAYER ME4 ;
  RECT 321.699 35.220 322.039 68.179 ;
 END
 PORT
  LAYER ME4 ;
  RECT 335.713 35.220 336.053 68.179 ;
 END
 PORT
  LAYER ME4 ;
  RECT 333.711 35.220 334.051 68.179 ;
 END
 PORT
  LAYER ME4 ;
  RECT 331.709 35.220 332.049 68.179 ;
 END
 PORT
  LAYER ME4 ;
  RECT 329.707 35.220 330.047 68.179 ;
 END
 PORT
  LAYER ME4 ;
  RECT 343.721 35.220 344.061 68.179 ;
 END
 PORT
  LAYER ME4 ;
  RECT 341.719 35.220 342.059 68.179 ;
 END
 PORT
  LAYER ME4 ;
  RECT 339.717 35.220 340.057 68.179 ;
 END
 PORT
  LAYER ME4 ;
  RECT 337.715 35.220 338.055 68.179 ;
 END
 PORT
  LAYER ME4 ;
  RECT 351.729 35.220 352.069 68.179 ;
 END
 PORT
  LAYER ME4 ;
  RECT 349.727 35.220 350.067 68.179 ;
 END
 PORT
  LAYER ME4 ;
  RECT 347.725 35.220 348.065 68.179 ;
 END
 PORT
  LAYER ME4 ;
  RECT 345.723 35.220 346.063 68.179 ;
 END
 PORT
  LAYER ME4 ;
  RECT 359.737 35.220 360.077 68.179 ;
 END
 PORT
  LAYER ME4 ;
  RECT 357.735 35.220 358.075 68.179 ;
 END
 PORT
  LAYER ME4 ;
  RECT 355.733 35.220 356.073 68.179 ;
 END
 PORT
  LAYER ME4 ;
  RECT 353.731 35.220 354.071 68.179 ;
 END
 PORT
  LAYER ME4 ;
  RECT 367.745 35.220 368.085 68.179 ;
 END
 PORT
  LAYER ME4 ;
  RECT 365.743 35.220 366.083 68.179 ;
 END
 PORT
  LAYER ME4 ;
  RECT 363.741 35.220 364.081 68.179 ;
 END
 PORT
  LAYER ME4 ;
  RECT 361.739 35.220 362.079 68.179 ;
 END
 PORT
  LAYER ME4 ;
  RECT 375.753 35.220 376.093 68.179 ;
 END
 PORT
  LAYER ME4 ;
  RECT 373.751 35.220 374.091 68.179 ;
 END
 PORT
  LAYER ME4 ;
  RECT 371.749 35.220 372.089 68.179 ;
 END
 PORT
  LAYER ME4 ;
  RECT 369.747 35.220 370.087 68.179 ;
 END
 PORT
  LAYER ME4 ;
  RECT 9.748 35.220 10.088 68.179 ;
 END
 PORT
  LAYER ME4 ;
  RECT 7.746 35.220 8.086 68.179 ;
 END
 PORT
  LAYER ME4 ;
  RECT 5.744 35.220 6.084 68.179 ;
 END
 PORT
  LAYER ME4 ;
  RECT 3.742 35.220 4.082 68.179 ;
 END
 PORT
  LAYER ME4 ;
  RECT 17.756 35.220 18.096 68.179 ;
 END
 PORT
  LAYER ME4 ;
  RECT 15.754 35.220 16.094 68.179 ;
 END
 PORT
  LAYER ME4 ;
  RECT 13.752 35.220 14.092 68.179 ;
 END
 PORT
  LAYER ME4 ;
  RECT 11.750 35.220 12.090 68.179 ;
 END
 PORT
  LAYER ME4 ;
  RECT 25.764 35.220 26.104 68.179 ;
 END
 PORT
  LAYER ME4 ;
  RECT 23.762 35.220 24.102 68.179 ;
 END
 PORT
  LAYER ME4 ;
  RECT 21.760 35.220 22.100 68.179 ;
 END
 PORT
  LAYER ME4 ;
  RECT 19.758 35.220 20.098 68.179 ;
 END
 PORT
  LAYER ME4 ;
  RECT 33.772 35.220 34.112 68.179 ;
 END
 PORT
  LAYER ME4 ;
  RECT 31.770 35.220 32.110 68.179 ;
 END
 PORT
  LAYER ME4 ;
  RECT 29.768 35.220 30.108 68.179 ;
 END
 PORT
  LAYER ME4 ;
  RECT 27.766 35.220 28.106 68.179 ;
 END
 PORT
  LAYER ME4 ;
  RECT 41.780 35.220 42.120 68.179 ;
 END
 PORT
  LAYER ME4 ;
  RECT 39.778 35.220 40.118 68.179 ;
 END
 PORT
  LAYER ME4 ;
  RECT 37.776 35.220 38.116 68.179 ;
 END
 PORT
  LAYER ME4 ;
  RECT 35.774 35.220 36.114 68.179 ;
 END
 PORT
  LAYER ME4 ;
  RECT 49.788 35.220 50.128 68.179 ;
 END
 PORT
  LAYER ME4 ;
  RECT 47.786 35.220 48.126 68.179 ;
 END
 PORT
  LAYER ME4 ;
  RECT 45.784 35.220 46.124 68.179 ;
 END
 PORT
  LAYER ME4 ;
  RECT 43.782 35.220 44.122 68.179 ;
 END
 PORT
  LAYER ME4 ;
  RECT 57.796 35.220 58.136 68.179 ;
 END
 PORT
  LAYER ME4 ;
  RECT 55.794 35.220 56.134 68.179 ;
 END
 PORT
  LAYER ME4 ;
  RECT 53.792 35.220 54.132 68.179 ;
 END
 PORT
  LAYER ME4 ;
  RECT 51.790 35.220 52.130 68.179 ;
 END
 PORT
  LAYER ME4 ;
  RECT 65.804 35.220 66.144 68.179 ;
 END
 PORT
  LAYER ME4 ;
  RECT 63.802 35.220 64.142 68.179 ;
 END
 PORT
  LAYER ME4 ;
  RECT 61.800 35.220 62.140 68.179 ;
 END
 PORT
  LAYER ME4 ;
  RECT 59.798 35.220 60.138 68.179 ;
 END
 PORT
  LAYER ME4 ;
  RECT 73.812 35.220 74.152 68.179 ;
 END
 PORT
  LAYER ME4 ;
  RECT 71.810 35.220 72.150 68.179 ;
 END
 PORT
  LAYER ME4 ;
  RECT 69.808 35.220 70.148 68.179 ;
 END
 PORT
  LAYER ME4 ;
  RECT 67.806 35.220 68.146 68.179 ;
 END
 PORT
  LAYER ME4 ;
  RECT 81.820 35.220 82.160 68.179 ;
 END
 PORT
  LAYER ME4 ;
  RECT 79.818 35.220 80.158 68.179 ;
 END
 PORT
  LAYER ME4 ;
  RECT 77.816 35.220 78.156 68.179 ;
 END
 PORT
  LAYER ME4 ;
  RECT 75.814 35.220 76.154 68.179 ;
 END
 PORT
  LAYER ME4 ;
  RECT 89.828 35.220 90.168 68.179 ;
 END
 PORT
  LAYER ME4 ;
  RECT 87.826 35.220 88.166 68.179 ;
 END
 PORT
  LAYER ME4 ;
  RECT 85.824 35.220 86.164 68.179 ;
 END
 PORT
  LAYER ME4 ;
  RECT 83.822 35.220 84.162 68.179 ;
 END
 PORT
  LAYER ME4 ;
  RECT 97.836 35.220 98.176 68.179 ;
 END
 PORT
  LAYER ME4 ;
  RECT 95.834 35.220 96.174 68.179 ;
 END
 PORT
  LAYER ME4 ;
  RECT 93.832 35.220 94.172 68.179 ;
 END
 PORT
  LAYER ME4 ;
  RECT 91.830 35.220 92.170 68.179 ;
 END
 PORT
  LAYER ME4 ;
  RECT 105.844 35.220 106.184 68.179 ;
 END
 PORT
  LAYER ME4 ;
  RECT 103.842 35.220 104.182 68.179 ;
 END
 PORT
  LAYER ME4 ;
  RECT 101.840 35.220 102.180 68.179 ;
 END
 PORT
  LAYER ME4 ;
  RECT 99.838 35.220 100.178 68.179 ;
 END
 PORT
  LAYER ME4 ;
  RECT 113.852 35.220 114.192 68.179 ;
 END
 PORT
  LAYER ME4 ;
  RECT 111.850 35.220 112.190 68.179 ;
 END
 PORT
  LAYER ME4 ;
  RECT 109.848 35.220 110.188 68.179 ;
 END
 PORT
  LAYER ME4 ;
  RECT 107.846 35.220 108.186 68.179 ;
 END
 PORT
  LAYER ME4 ;
  RECT 121.860 35.220 122.200 68.179 ;
 END
 PORT
  LAYER ME4 ;
  RECT 119.858 35.220 120.198 68.179 ;
 END
 PORT
  LAYER ME4 ;
  RECT 117.856 35.220 118.196 68.179 ;
 END
 PORT
  LAYER ME4 ;
  RECT 115.854 35.220 116.194 68.179 ;
 END
 PORT
  LAYER ME4 ;
  RECT 129.868 35.220 130.208 68.179 ;
 END
 PORT
  LAYER ME4 ;
  RECT 127.866 35.220 128.206 68.179 ;
 END
 PORT
  LAYER ME4 ;
  RECT 125.864 35.220 126.204 68.179 ;
 END
 PORT
  LAYER ME4 ;
  RECT 123.862 35.220 124.202 68.179 ;
 END
 PORT
  LAYER ME4 ;
  RECT 137.876 35.220 138.216 68.179 ;
 END
 PORT
  LAYER ME4 ;
  RECT 135.874 35.220 136.214 68.179 ;
 END
 PORT
  LAYER ME4 ;
  RECT 133.872 35.220 134.212 68.179 ;
 END
 PORT
  LAYER ME4 ;
  RECT 131.870 35.220 132.210 68.179 ;
 END
 PORT
  LAYER ME4 ;
  RECT 145.884 35.220 146.224 68.179 ;
 END
 PORT
  LAYER ME4 ;
  RECT 143.882 35.220 144.222 68.179 ;
 END
 PORT
  LAYER ME4 ;
  RECT 141.880 35.220 142.220 68.179 ;
 END
 PORT
  LAYER ME4 ;
  RECT 139.878 35.220 140.218 68.179 ;
 END
 PORT
  LAYER ME4 ;
  RECT 153.892 35.220 154.232 68.179 ;
 END
 PORT
  LAYER ME4 ;
  RECT 151.890 35.220 152.230 68.179 ;
 END
 PORT
  LAYER ME4 ;
  RECT 149.888 35.220 150.228 68.179 ;
 END
 PORT
  LAYER ME4 ;
  RECT 147.886 35.220 148.226 68.179 ;
 END
 PORT
  LAYER ME4 ;
  RECT 161.900 35.220 162.240 68.179 ;
 END
 PORT
  LAYER ME4 ;
  RECT 159.898 35.220 160.238 68.179 ;
 END
 PORT
  LAYER ME4 ;
  RECT 157.896 35.220 158.236 68.179 ;
 END
 PORT
  LAYER ME4 ;
  RECT 155.894 35.220 156.234 68.179 ;
 END
 PORT
  LAYER ME4 ;
  RECT 169.908 35.220 170.248 68.179 ;
 END
 PORT
  LAYER ME4 ;
  RECT 167.906 35.220 168.246 68.179 ;
 END
 PORT
  LAYER ME4 ;
  RECT 165.904 35.220 166.244 68.179 ;
 END
 PORT
  LAYER ME4 ;
  RECT 163.902 35.220 164.242 68.179 ;
 END
END VCC
PIN GND
  DIRECTION INOUT ;
  USE GROUND ;
 PORT
  LAYER ME4 ;
  RECT 208.586 0.921 208.926 68.179 ;
 END
 PORT
  LAYER ME4 ;
  RECT 215.403 0.000 216.123 31.570 ;
 END
 PORT
  LAYER ME4 ;
  RECT 216.594 0.000 216.934 68.179 ;
 END
 PORT
  LAYER ME4 ;
  RECT 210.588 0.000 210.928 68.179 ;
 END
 PORT
  LAYER ME4 ;
  RECT 211.399 0.000 212.119 31.570 ;
 END
 PORT
  LAYER ME4 ;
  RECT 212.590 0.921 212.930 68.179 ;
 END
 PORT
  LAYER ME4 ;
  RECT 214.592 0.921 214.932 68.179 ;
 END
 PORT
  LAYER ME4 ;
  RECT 223.411 0.000 224.131 31.570 ;
 END
 PORT
  LAYER ME4 ;
  RECT 224.602 0.000 224.942 68.179 ;
 END
 PORT
  LAYER ME4 ;
  RECT 218.596 0.000 218.936 68.179 ;
 END
 PORT
  LAYER ME4 ;
  RECT 219.407 0.000 220.127 31.570 ;
 END
 PORT
  LAYER ME4 ;
  RECT 220.598 0.921 220.938 68.179 ;
 END
 PORT
  LAYER ME4 ;
  RECT 222.600 0.921 222.940 68.179 ;
 END
 PORT
  LAYER ME4 ;
  RECT 231.419 0.000 232.139 31.570 ;
 END
 PORT
  LAYER ME4 ;
  RECT 232.610 0.000 232.950 68.179 ;
 END
 PORT
  LAYER ME4 ;
  RECT 226.604 0.000 226.944 68.179 ;
 END
 PORT
  LAYER ME4 ;
  RECT 227.415 0.000 228.135 31.570 ;
 END
 PORT
  LAYER ME4 ;
  RECT 228.606 0.921 228.946 68.179 ;
 END
 PORT
  LAYER ME4 ;
  RECT 230.608 0.921 230.948 68.179 ;
 END
 PORT
  LAYER ME4 ;
  RECT 239.427 0.000 240.147 31.570 ;
 END
 PORT
  LAYER ME4 ;
  RECT 240.618 0.000 240.958 68.179 ;
 END
 PORT
  LAYER ME4 ;
  RECT 234.612 0.000 234.952 68.179 ;
 END
 PORT
  LAYER ME4 ;
  RECT 235.423 0.000 236.143 31.570 ;
 END
 PORT
  LAYER ME4 ;
  RECT 236.614 0.921 236.954 68.179 ;
 END
 PORT
  LAYER ME4 ;
  RECT 238.616 0.921 238.956 68.179 ;
 END
 PORT
  LAYER ME4 ;
  RECT 247.435 0.000 248.155 31.570 ;
 END
 PORT
  LAYER ME4 ;
  RECT 248.626 0.000 248.966 68.179 ;
 END
 PORT
  LAYER ME4 ;
  RECT 242.620 0.000 242.960 68.179 ;
 END
 PORT
  LAYER ME4 ;
  RECT 243.431 0.000 244.151 31.570 ;
 END
 PORT
  LAYER ME4 ;
  RECT 244.622 0.921 244.962 68.179 ;
 END
 PORT
  LAYER ME4 ;
  RECT 246.624 0.921 246.964 68.179 ;
 END
 PORT
  LAYER ME4 ;
  RECT 255.443 0.000 256.163 31.570 ;
 END
 PORT
  LAYER ME4 ;
  RECT 256.634 0.000 256.974 68.179 ;
 END
 PORT
  LAYER ME4 ;
  RECT 250.628 0.000 250.968 68.179 ;
 END
 PORT
  LAYER ME4 ;
  RECT 251.439 0.000 252.159 31.570 ;
 END
 PORT
  LAYER ME4 ;
  RECT 252.630 0.921 252.970 68.179 ;
 END
 PORT
  LAYER ME4 ;
  RECT 254.632 0.921 254.972 68.179 ;
 END
 PORT
  LAYER ME4 ;
  RECT 263.451 0.000 264.171 31.570 ;
 END
 PORT
  LAYER ME4 ;
  RECT 264.642 0.000 264.982 68.179 ;
 END
 PORT
  LAYER ME4 ;
  RECT 258.636 0.000 258.976 68.179 ;
 END
 PORT
  LAYER ME4 ;
  RECT 259.447 0.000 260.167 31.570 ;
 END
 PORT
  LAYER ME4 ;
  RECT 260.638 0.921 260.978 68.179 ;
 END
 PORT
  LAYER ME4 ;
  RECT 262.640 0.921 262.980 68.179 ;
 END
 PORT
  LAYER ME4 ;
  RECT 271.459 0.000 272.179 31.570 ;
 END
 PORT
  LAYER ME4 ;
  RECT 272.650 0.000 272.990 68.179 ;
 END
 PORT
  LAYER ME4 ;
  RECT 266.644 0.000 266.984 68.179 ;
 END
 PORT
  LAYER ME4 ;
  RECT 267.455 0.000 268.175 31.570 ;
 END
 PORT
  LAYER ME4 ;
  RECT 268.646 0.921 268.986 68.179 ;
 END
 PORT
  LAYER ME4 ;
  RECT 270.648 0.921 270.988 68.179 ;
 END
 PORT
  LAYER ME4 ;
  RECT 279.467 0.000 280.187 31.570 ;
 END
 PORT
  LAYER ME4 ;
  RECT 280.658 0.000 280.998 68.179 ;
 END
 PORT
  LAYER ME4 ;
  RECT 274.652 0.000 274.992 68.179 ;
 END
 PORT
  LAYER ME4 ;
  RECT 275.463 0.000 276.183 31.570 ;
 END
 PORT
  LAYER ME4 ;
  RECT 276.654 0.921 276.994 68.179 ;
 END
 PORT
  LAYER ME4 ;
  RECT 278.656 0.921 278.996 68.179 ;
 END
 PORT
  LAYER ME4 ;
  RECT 287.475 0.000 288.195 31.570 ;
 END
 PORT
  LAYER ME4 ;
  RECT 288.666 0.000 289.006 68.179 ;
 END
 PORT
  LAYER ME4 ;
  RECT 282.660 0.000 283.000 68.179 ;
 END
 PORT
  LAYER ME4 ;
  RECT 283.471 0.000 284.191 31.570 ;
 END
 PORT
  LAYER ME4 ;
  RECT 284.662 0.921 285.002 68.179 ;
 END
 PORT
  LAYER ME4 ;
  RECT 286.664 0.921 287.004 68.179 ;
 END
 PORT
  LAYER ME4 ;
  RECT 295.483 0.000 296.203 31.570 ;
 END
 PORT
  LAYER ME4 ;
  RECT 296.674 0.000 297.014 68.179 ;
 END
 PORT
  LAYER ME4 ;
  RECT 290.668 0.000 291.008 68.179 ;
 END
 PORT
  LAYER ME4 ;
  RECT 291.479 0.000 292.199 31.570 ;
 END
 PORT
  LAYER ME4 ;
  RECT 292.670 0.921 293.010 68.179 ;
 END
 PORT
  LAYER ME4 ;
  RECT 294.672 0.921 295.012 68.179 ;
 END
 PORT
  LAYER ME4 ;
  RECT 303.491 0.000 304.211 31.570 ;
 END
 PORT
  LAYER ME4 ;
  RECT 304.682 0.000 305.022 68.179 ;
 END
 PORT
  LAYER ME4 ;
  RECT 298.676 0.000 299.016 68.179 ;
 END
 PORT
  LAYER ME4 ;
  RECT 299.487 0.000 300.207 31.570 ;
 END
 PORT
  LAYER ME4 ;
  RECT 300.678 0.921 301.018 68.179 ;
 END
 PORT
  LAYER ME4 ;
  RECT 302.680 0.921 303.020 68.179 ;
 END
 PORT
  LAYER ME4 ;
  RECT 311.499 0.000 312.219 31.570 ;
 END
 PORT
  LAYER ME4 ;
  RECT 312.690 0.000 313.030 68.179 ;
 END
 PORT
  LAYER ME4 ;
  RECT 306.684 0.000 307.024 68.179 ;
 END
 PORT
  LAYER ME4 ;
  RECT 307.495 0.000 308.215 31.570 ;
 END
 PORT
  LAYER ME4 ;
  RECT 308.686 0.921 309.026 68.179 ;
 END
 PORT
  LAYER ME4 ;
  RECT 310.688 0.921 311.028 68.179 ;
 END
 PORT
  LAYER ME4 ;
  RECT 319.507 0.000 320.227 31.570 ;
 END
 PORT
  LAYER ME4 ;
  RECT 320.698 0.000 321.038 68.179 ;
 END
 PORT
  LAYER ME4 ;
  RECT 314.692 0.000 315.032 68.179 ;
 END
 PORT
  LAYER ME4 ;
  RECT 315.503 0.000 316.223 31.570 ;
 END
 PORT
  LAYER ME4 ;
  RECT 316.694 0.921 317.034 68.179 ;
 END
 PORT
  LAYER ME4 ;
  RECT 318.696 0.921 319.036 68.179 ;
 END
 PORT
  LAYER ME4 ;
  RECT 327.515 0.000 328.235 31.570 ;
 END
 PORT
  LAYER ME4 ;
  RECT 328.706 0.000 329.046 68.179 ;
 END
 PORT
  LAYER ME4 ;
  RECT 322.700 0.000 323.040 68.179 ;
 END
 PORT
  LAYER ME4 ;
  RECT 323.511 0.000 324.231 31.570 ;
 END
 PORT
  LAYER ME4 ;
  RECT 324.702 0.921 325.042 68.179 ;
 END
 PORT
  LAYER ME4 ;
  RECT 326.704 0.921 327.044 68.179 ;
 END
 PORT
  LAYER ME4 ;
  RECT 335.523 0.000 336.243 31.570 ;
 END
 PORT
  LAYER ME4 ;
  RECT 336.714 0.000 337.054 68.179 ;
 END
 PORT
  LAYER ME4 ;
  RECT 330.708 0.000 331.048 68.179 ;
 END
 PORT
  LAYER ME4 ;
  RECT 331.519 0.000 332.239 31.570 ;
 END
 PORT
  LAYER ME4 ;
  RECT 332.710 0.921 333.050 68.179 ;
 END
 PORT
  LAYER ME4 ;
  RECT 334.712 0.921 335.052 68.179 ;
 END
 PORT
  LAYER ME4 ;
  RECT 343.531 0.000 344.251 31.570 ;
 END
 PORT
  LAYER ME4 ;
  RECT 344.722 0.000 345.062 68.179 ;
 END
 PORT
  LAYER ME4 ;
  RECT 338.716 0.000 339.056 68.179 ;
 END
 PORT
  LAYER ME4 ;
  RECT 339.527 0.000 340.247 31.570 ;
 END
 PORT
  LAYER ME4 ;
  RECT 340.718 0.921 341.058 68.179 ;
 END
 PORT
  LAYER ME4 ;
  RECT 342.720 0.921 343.060 68.179 ;
 END
 PORT
  LAYER ME4 ;
  RECT 351.539 0.000 352.259 31.570 ;
 END
 PORT
  LAYER ME4 ;
  RECT 352.730 0.000 353.070 68.179 ;
 END
 PORT
  LAYER ME4 ;
  RECT 346.724 0.000 347.064 68.179 ;
 END
 PORT
  LAYER ME4 ;
  RECT 347.535 0.000 348.255 31.570 ;
 END
 PORT
  LAYER ME4 ;
  RECT 348.726 0.921 349.066 68.179 ;
 END
 PORT
  LAYER ME4 ;
  RECT 350.728 0.921 351.068 68.179 ;
 END
 PORT
  LAYER ME4 ;
  RECT 359.547 0.000 360.267 31.570 ;
 END
 PORT
  LAYER ME4 ;
  RECT 360.738 0.000 361.078 68.179 ;
 END
 PORT
  LAYER ME4 ;
  RECT 354.732 0.000 355.072 68.179 ;
 END
 PORT
  LAYER ME4 ;
  RECT 355.543 0.000 356.263 31.570 ;
 END
 PORT
  LAYER ME4 ;
  RECT 356.734 0.921 357.074 68.179 ;
 END
 PORT
  LAYER ME4 ;
  RECT 358.736 0.921 359.076 68.179 ;
 END
 PORT
  LAYER ME4 ;
  RECT 367.555 0.000 368.275 31.570 ;
 END
 PORT
  LAYER ME4 ;
  RECT 368.746 0.000 369.086 68.179 ;
 END
 PORT
  LAYER ME4 ;
  RECT 362.740 0.000 363.080 68.179 ;
 END
 PORT
  LAYER ME4 ;
  RECT 363.551 0.000 364.271 31.570 ;
 END
 PORT
  LAYER ME4 ;
  RECT 364.742 0.921 365.082 68.179 ;
 END
 PORT
  LAYER ME4 ;
  RECT 366.744 0.921 367.084 68.179 ;
 END
 PORT
  LAYER ME4 ;
  RECT 375.563 0.000 376.283 31.570 ;
 END
 PORT
  LAYER ME4 ;
  RECT 376.754 0.000 377.094 68.179 ;
 END
 PORT
  LAYER ME4 ;
  RECT 370.748 0.000 371.088 68.179 ;
 END
 PORT
  LAYER ME4 ;
  RECT 371.559 0.000 372.279 31.570 ;
 END
 PORT
  LAYER ME4 ;
  RECT 372.750 0.921 373.090 68.179 ;
 END
 PORT
  LAYER ME4 ;
  RECT 374.752 0.921 375.092 68.179 ;
 END
 PORT
  LAYER ME4 ;
  RECT 377.755 0.000 378.095 68.179 ;
 END
 PORT
  LAYER ME4 ;
  RECT 189.729 0.000 190.449 68.179 ;
 END
 PORT
  LAYER ME4 ;
  RECT 195.723 0.000 196.443 68.179 ;
 END
 PORT
  LAYER ME4 ;
  RECT 201.194 0.000 201.914 68.179 ;
 END
 PORT
  LAYER ME4 ;
  RECT 202.909 0.000 203.629 68.179 ;
 END
 PORT
  LAYER ME4 ;
  RECT 205.905 0.000 206.505 68.179 ;
 END
 PORT
  LAYER ME4 ;
  RECT 207.585 0.921 207.925 68.179 ;
 END
 PORT
  LAYER ME4 ;
  RECT 182.170 0.000 182.890 68.179 ;
 END
 PORT
  LAYER ME4 ;
  RECT 180.130 0.921 180.850 67.420 ;
 END
 PORT
  LAYER ME4 ;
  RECT 178.010 0.000 178.730 68.179 ;
 END
 PORT
  LAYER ME4 ;
  RECT 175.970 0.921 176.690 68.179 ;
 END
 PORT
  LAYER ME4 ;
  RECT 1.740 0.000 2.080 68.179 ;
 END
 PORT
  LAYER ME4 ;
  RECT 2.741 0.921 3.081 68.179 ;
 END
 PORT
  LAYER ME4 ;
  RECT 9.558 0.000 10.278 31.570 ;
 END
 PORT
  LAYER ME4 ;
  RECT 10.749 0.000 11.089 68.179 ;
 END
 PORT
  LAYER ME4 ;
  RECT 4.743 0.000 5.083 68.179 ;
 END
 PORT
  LAYER ME4 ;
  RECT 5.554 0.000 6.274 31.570 ;
 END
 PORT
  LAYER ME4 ;
  RECT 6.745 0.921 7.085 68.179 ;
 END
 PORT
  LAYER ME4 ;
  RECT 8.747 0.921 9.087 68.179 ;
 END
 PORT
  LAYER ME4 ;
  RECT 17.566 0.000 18.286 31.570 ;
 END
 PORT
  LAYER ME4 ;
  RECT 18.757 0.000 19.097 68.179 ;
 END
 PORT
  LAYER ME4 ;
  RECT 12.751 0.000 13.091 68.179 ;
 END
 PORT
  LAYER ME4 ;
  RECT 13.562 0.000 14.282 31.570 ;
 END
 PORT
  LAYER ME4 ;
  RECT 14.753 0.921 15.093 68.179 ;
 END
 PORT
  LAYER ME4 ;
  RECT 16.755 0.921 17.095 68.179 ;
 END
 PORT
  LAYER ME4 ;
  RECT 25.574 0.000 26.294 31.570 ;
 END
 PORT
  LAYER ME4 ;
  RECT 26.765 0.000 27.105 68.179 ;
 END
 PORT
  LAYER ME4 ;
  RECT 20.759 0.000 21.099 68.179 ;
 END
 PORT
  LAYER ME4 ;
  RECT 21.570 0.000 22.290 31.570 ;
 END
 PORT
  LAYER ME4 ;
  RECT 22.761 0.921 23.101 68.179 ;
 END
 PORT
  LAYER ME4 ;
  RECT 24.763 0.921 25.103 68.179 ;
 END
 PORT
  LAYER ME4 ;
  RECT 33.582 0.000 34.302 31.570 ;
 END
 PORT
  LAYER ME4 ;
  RECT 34.773 0.000 35.113 68.179 ;
 END
 PORT
  LAYER ME4 ;
  RECT 28.767 0.000 29.107 68.179 ;
 END
 PORT
  LAYER ME4 ;
  RECT 29.578 0.000 30.298 31.570 ;
 END
 PORT
  LAYER ME4 ;
  RECT 30.769 0.921 31.109 68.179 ;
 END
 PORT
  LAYER ME4 ;
  RECT 32.771 0.921 33.111 68.179 ;
 END
 PORT
  LAYER ME4 ;
  RECT 41.590 0.000 42.310 31.570 ;
 END
 PORT
  LAYER ME4 ;
  RECT 42.781 0.000 43.121 68.179 ;
 END
 PORT
  LAYER ME4 ;
  RECT 36.775 0.000 37.115 68.179 ;
 END
 PORT
  LAYER ME4 ;
  RECT 37.586 0.000 38.306 31.570 ;
 END
 PORT
  LAYER ME4 ;
  RECT 38.777 0.921 39.117 68.179 ;
 END
 PORT
  LAYER ME4 ;
  RECT 40.779 0.921 41.119 68.179 ;
 END
 PORT
  LAYER ME4 ;
  RECT 49.598 0.000 50.318 31.570 ;
 END
 PORT
  LAYER ME4 ;
  RECT 50.789 0.000 51.129 68.179 ;
 END
 PORT
  LAYER ME4 ;
  RECT 44.783 0.000 45.123 68.179 ;
 END
 PORT
  LAYER ME4 ;
  RECT 45.594 0.000 46.314 31.570 ;
 END
 PORT
  LAYER ME4 ;
  RECT 46.785 0.921 47.125 68.179 ;
 END
 PORT
  LAYER ME4 ;
  RECT 48.787 0.921 49.127 68.179 ;
 END
 PORT
  LAYER ME4 ;
  RECT 57.606 0.000 58.326 31.570 ;
 END
 PORT
  LAYER ME4 ;
  RECT 58.797 0.000 59.137 68.179 ;
 END
 PORT
  LAYER ME4 ;
  RECT 52.791 0.000 53.131 68.179 ;
 END
 PORT
  LAYER ME4 ;
  RECT 53.602 0.000 54.322 31.570 ;
 END
 PORT
  LAYER ME4 ;
  RECT 54.793 0.921 55.133 68.179 ;
 END
 PORT
  LAYER ME4 ;
  RECT 56.795 0.921 57.135 68.179 ;
 END
 PORT
  LAYER ME4 ;
  RECT 65.614 0.000 66.334 31.570 ;
 END
 PORT
  LAYER ME4 ;
  RECT 66.805 0.000 67.145 68.179 ;
 END
 PORT
  LAYER ME4 ;
  RECT 60.799 0.000 61.139 68.179 ;
 END
 PORT
  LAYER ME4 ;
  RECT 61.610 0.000 62.330 31.570 ;
 END
 PORT
  LAYER ME4 ;
  RECT 62.801 0.921 63.141 68.179 ;
 END
 PORT
  LAYER ME4 ;
  RECT 64.803 0.921 65.143 68.179 ;
 END
 PORT
  LAYER ME4 ;
  RECT 73.622 0.000 74.342 31.570 ;
 END
 PORT
  LAYER ME4 ;
  RECT 74.813 0.000 75.153 68.179 ;
 END
 PORT
  LAYER ME4 ;
  RECT 68.807 0.000 69.147 68.179 ;
 END
 PORT
  LAYER ME4 ;
  RECT 69.618 0.000 70.338 31.570 ;
 END
 PORT
  LAYER ME4 ;
  RECT 70.809 0.921 71.149 68.179 ;
 END
 PORT
  LAYER ME4 ;
  RECT 72.811 0.921 73.151 68.179 ;
 END
 PORT
  LAYER ME4 ;
  RECT 81.630 0.000 82.350 31.570 ;
 END
 PORT
  LAYER ME4 ;
  RECT 82.821 0.000 83.161 68.179 ;
 END
 PORT
  LAYER ME4 ;
  RECT 76.815 0.000 77.155 68.179 ;
 END
 PORT
  LAYER ME4 ;
  RECT 77.626 0.000 78.346 31.570 ;
 END
 PORT
  LAYER ME4 ;
  RECT 78.817 0.921 79.157 68.179 ;
 END
 PORT
  LAYER ME4 ;
  RECT 80.819 0.921 81.159 68.179 ;
 END
 PORT
  LAYER ME4 ;
  RECT 89.638 0.000 90.358 31.570 ;
 END
 PORT
  LAYER ME4 ;
  RECT 90.829 0.000 91.169 68.179 ;
 END
 PORT
  LAYER ME4 ;
  RECT 84.823 0.000 85.163 68.179 ;
 END
 PORT
  LAYER ME4 ;
  RECT 85.634 0.000 86.354 31.570 ;
 END
 PORT
  LAYER ME4 ;
  RECT 86.825 0.921 87.165 68.179 ;
 END
 PORT
  LAYER ME4 ;
  RECT 88.827 0.921 89.167 68.179 ;
 END
 PORT
  LAYER ME4 ;
  RECT 97.646 0.000 98.366 31.570 ;
 END
 PORT
  LAYER ME4 ;
  RECT 98.837 0.000 99.177 68.179 ;
 END
 PORT
  LAYER ME4 ;
  RECT 92.831 0.000 93.171 68.179 ;
 END
 PORT
  LAYER ME4 ;
  RECT 93.642 0.000 94.362 31.570 ;
 END
 PORT
  LAYER ME4 ;
  RECT 94.833 0.921 95.173 68.179 ;
 END
 PORT
  LAYER ME4 ;
  RECT 96.835 0.921 97.175 68.179 ;
 END
 PORT
  LAYER ME4 ;
  RECT 105.654 0.000 106.374 31.570 ;
 END
 PORT
  LAYER ME4 ;
  RECT 106.845 0.000 107.185 68.179 ;
 END
 PORT
  LAYER ME4 ;
  RECT 100.839 0.000 101.179 68.179 ;
 END
 PORT
  LAYER ME4 ;
  RECT 101.650 0.000 102.370 31.570 ;
 END
 PORT
  LAYER ME4 ;
  RECT 102.841 0.921 103.181 68.179 ;
 END
 PORT
  LAYER ME4 ;
  RECT 104.843 0.921 105.183 68.179 ;
 END
 PORT
  LAYER ME4 ;
  RECT 113.662 0.000 114.382 31.570 ;
 END
 PORT
  LAYER ME4 ;
  RECT 114.853 0.000 115.193 68.179 ;
 END
 PORT
  LAYER ME4 ;
  RECT 108.847 0.000 109.187 68.179 ;
 END
 PORT
  LAYER ME4 ;
  RECT 109.658 0.000 110.378 31.570 ;
 END
 PORT
  LAYER ME4 ;
  RECT 110.849 0.921 111.189 68.179 ;
 END
 PORT
  LAYER ME4 ;
  RECT 112.851 0.921 113.191 68.179 ;
 END
 PORT
  LAYER ME4 ;
  RECT 121.670 0.000 122.390 31.570 ;
 END
 PORT
  LAYER ME4 ;
  RECT 122.861 0.000 123.201 68.179 ;
 END
 PORT
  LAYER ME4 ;
  RECT 116.855 0.000 117.195 68.179 ;
 END
 PORT
  LAYER ME4 ;
  RECT 117.666 0.000 118.386 31.570 ;
 END
 PORT
  LAYER ME4 ;
  RECT 118.857 0.921 119.197 68.179 ;
 END
 PORT
  LAYER ME4 ;
  RECT 120.859 0.921 121.199 68.179 ;
 END
 PORT
  LAYER ME4 ;
  RECT 129.678 0.000 130.398 31.570 ;
 END
 PORT
  LAYER ME4 ;
  RECT 130.869 0.000 131.209 68.179 ;
 END
 PORT
  LAYER ME4 ;
  RECT 124.863 0.000 125.203 68.179 ;
 END
 PORT
  LAYER ME4 ;
  RECT 125.674 0.000 126.394 31.570 ;
 END
 PORT
  LAYER ME4 ;
  RECT 126.865 0.921 127.205 68.179 ;
 END
 PORT
  LAYER ME4 ;
  RECT 128.867 0.921 129.207 68.179 ;
 END
 PORT
  LAYER ME4 ;
  RECT 137.686 0.000 138.406 31.570 ;
 END
 PORT
  LAYER ME4 ;
  RECT 138.877 0.000 139.217 68.179 ;
 END
 PORT
  LAYER ME4 ;
  RECT 132.871 0.000 133.211 68.179 ;
 END
 PORT
  LAYER ME4 ;
  RECT 133.682 0.000 134.402 31.570 ;
 END
 PORT
  LAYER ME4 ;
  RECT 134.873 0.921 135.213 68.179 ;
 END
 PORT
  LAYER ME4 ;
  RECT 136.875 0.921 137.215 68.179 ;
 END
 PORT
  LAYER ME4 ;
  RECT 145.694 0.000 146.414 31.570 ;
 END
 PORT
  LAYER ME4 ;
  RECT 146.885 0.000 147.225 68.179 ;
 END
 PORT
  LAYER ME4 ;
  RECT 140.879 0.000 141.219 68.179 ;
 END
 PORT
  LAYER ME4 ;
  RECT 141.690 0.000 142.410 31.570 ;
 END
 PORT
  LAYER ME4 ;
  RECT 142.881 0.921 143.221 68.179 ;
 END
 PORT
  LAYER ME4 ;
  RECT 144.883 0.921 145.223 68.179 ;
 END
 PORT
  LAYER ME4 ;
  RECT 153.702 0.000 154.422 31.570 ;
 END
 PORT
  LAYER ME4 ;
  RECT 154.893 0.000 155.233 68.179 ;
 END
 PORT
  LAYER ME4 ;
  RECT 148.887 0.000 149.227 68.179 ;
 END
 PORT
  LAYER ME4 ;
  RECT 149.698 0.000 150.418 31.570 ;
 END
 PORT
  LAYER ME4 ;
  RECT 150.889 0.921 151.229 68.179 ;
 END
 PORT
  LAYER ME4 ;
  RECT 152.891 0.921 153.231 68.179 ;
 END
 PORT
  LAYER ME4 ;
  RECT 161.710 0.000 162.430 31.570 ;
 END
 PORT
  LAYER ME4 ;
  RECT 162.901 0.000 163.241 68.179 ;
 END
 PORT
  LAYER ME4 ;
  RECT 156.895 0.000 157.235 68.179 ;
 END
 PORT
  LAYER ME4 ;
  RECT 157.706 0.000 158.426 31.570 ;
 END
 PORT
  LAYER ME4 ;
  RECT 158.897 0.921 159.237 68.179 ;
 END
 PORT
  LAYER ME4 ;
  RECT 160.899 0.921 161.239 68.179 ;
 END
 PORT
  LAYER ME4 ;
  RECT 169.718 0.000 170.438 31.570 ;
 END
 PORT
  LAYER ME4 ;
  RECT 170.909 0.000 171.249 68.179 ;
 END
 PORT
  LAYER ME4 ;
  RECT 164.903 0.000 165.243 68.179 ;
 END
 PORT
  LAYER ME4 ;
  RECT 165.714 0.000 166.434 31.570 ;
 END
 PORT
  LAYER ME4 ;
  RECT 166.905 0.921 167.245 68.179 ;
 END
 PORT
  LAYER ME4 ;
  RECT 168.907 0.921 169.247 68.179 ;
 END
 PORT
  LAYER ME4 ;
  RECT 173.850 0.000 174.570 68.179 ;
 END
 PORT
  LAYER ME4 ;
  RECT 171.910 0.000 172.250 68.179 ;
 END
END GND
PIN DI20
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 168.766 0.000 169.046 0.720 ;
  LAYER ME3 ;
  RECT 168.766 0.000 169.046 0.720 ;
  LAYER ME2 ;
  RECT 168.766 0.000 169.046 0.720 ;
  LAYER ME1 ;
  RECT 168.766 0.000 169.046 0.720 ;
 END
 ANTENNAPARTIALMETALAREA                  0.805 LAYER ME1 ;
 ANTENNAGATEAREA                          0.072 LAYER ME1 ;
 ANTENNAGATEAREA                          0.072 LAYER ME2 ;
 ANTENNAGATEAREA                          0.072 LAYER ME3 ;
 ANTENNAGATEAREA                          0.072 LAYER ME4 ;
 ANTENNADIFFAREA                          0.218 LAYER ME1 ;
 ANTENNADIFFAREA                          0.218 LAYER ME2 ;
 ANTENNADIFFAREA                          0.218 LAYER ME3 ;
 ANTENNADIFFAREA                          0.218 LAYER ME4 ;
 ANTENNAMAXAREACAR                       13.984 LAYER ME1 ;
 ANTENNAMAXAREACAR                       16.784 LAYER ME2 ;
 ANTENNAMAXAREACAR                       19.584 LAYER ME3 ;
 ANTENNAMAXAREACAR                       22.384 LAYER ME4 ;
END DI20
PIN DO20
  DIRECTION OUTPUT ;
 PORT
  LAYER ME4 ;
  RECT 166.788 0.000 167.068 0.720 ;
  LAYER ME3 ;
  RECT 166.788 0.000 167.068 0.720 ;
  LAYER ME2 ;
  RECT 166.788 0.000 167.068 0.720 ;
  LAYER ME1 ;
  RECT 166.788 0.000 167.068 0.720 ;
 END
 ANTENNAPARTIALMETALAREA                  2.030 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME3 ;
 ANTENNADIFFAREA                          1.293 LAYER ME4 ;
END DO20
PIN DI19
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 160.758 0.000 161.038 0.720 ;
  LAYER ME3 ;
  RECT 160.758 0.000 161.038 0.720 ;
  LAYER ME2 ;
  RECT 160.758 0.000 161.038 0.720 ;
  LAYER ME1 ;
  RECT 160.758 0.000 161.038 0.720 ;
 END
 ANTENNAPARTIALMETALAREA                  0.805 LAYER ME1 ;
 ANTENNAGATEAREA                          0.072 LAYER ME1 ;
 ANTENNAGATEAREA                          0.072 LAYER ME2 ;
 ANTENNAGATEAREA                          0.072 LAYER ME3 ;
 ANTENNAGATEAREA                          0.072 LAYER ME4 ;
 ANTENNADIFFAREA                          0.218 LAYER ME1 ;
 ANTENNADIFFAREA                          0.218 LAYER ME2 ;
 ANTENNADIFFAREA                          0.218 LAYER ME3 ;
 ANTENNADIFFAREA                          0.218 LAYER ME4 ;
 ANTENNAMAXAREACAR                       13.984 LAYER ME1 ;
 ANTENNAMAXAREACAR                       16.784 LAYER ME2 ;
 ANTENNAMAXAREACAR                       19.584 LAYER ME3 ;
 ANTENNAMAXAREACAR                       22.384 LAYER ME4 ;
END DI19
PIN DO19
  DIRECTION OUTPUT ;
 PORT
  LAYER ME4 ;
  RECT 158.780 0.000 159.060 0.720 ;
  LAYER ME3 ;
  RECT 158.780 0.000 159.060 0.720 ;
  LAYER ME2 ;
  RECT 158.780 0.000 159.060 0.720 ;
  LAYER ME1 ;
  RECT 158.780 0.000 159.060 0.720 ;
 END
 ANTENNAPARTIALMETALAREA                  2.030 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME3 ;
 ANTENNADIFFAREA                          1.293 LAYER ME4 ;
END DO19
PIN DI18
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 152.750 0.000 153.030 0.720 ;
  LAYER ME3 ;
  RECT 152.750 0.000 153.030 0.720 ;
  LAYER ME2 ;
  RECT 152.750 0.000 153.030 0.720 ;
  LAYER ME1 ;
  RECT 152.750 0.000 153.030 0.720 ;
 END
 ANTENNAPARTIALMETALAREA                  0.805 LAYER ME1 ;
 ANTENNAGATEAREA                          0.072 LAYER ME1 ;
 ANTENNAGATEAREA                          0.072 LAYER ME2 ;
 ANTENNAGATEAREA                          0.072 LAYER ME3 ;
 ANTENNAGATEAREA                          0.072 LAYER ME4 ;
 ANTENNADIFFAREA                          0.218 LAYER ME1 ;
 ANTENNADIFFAREA                          0.218 LAYER ME2 ;
 ANTENNADIFFAREA                          0.218 LAYER ME3 ;
 ANTENNADIFFAREA                          0.218 LAYER ME4 ;
 ANTENNAMAXAREACAR                       13.984 LAYER ME1 ;
 ANTENNAMAXAREACAR                       16.784 LAYER ME2 ;
 ANTENNAMAXAREACAR                       19.584 LAYER ME3 ;
 ANTENNAMAXAREACAR                       22.384 LAYER ME4 ;
END DI18
PIN DO18
  DIRECTION OUTPUT ;
 PORT
  LAYER ME4 ;
  RECT 150.772 0.000 151.052 0.720 ;
  LAYER ME3 ;
  RECT 150.772 0.000 151.052 0.720 ;
  LAYER ME2 ;
  RECT 150.772 0.000 151.052 0.720 ;
  LAYER ME1 ;
  RECT 150.772 0.000 151.052 0.720 ;
 END
 ANTENNAPARTIALMETALAREA                  2.030 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME3 ;
 ANTENNADIFFAREA                          1.293 LAYER ME4 ;
END DO18
PIN DI17
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 144.742 0.000 145.022 0.720 ;
  LAYER ME3 ;
  RECT 144.742 0.000 145.022 0.720 ;
  LAYER ME2 ;
  RECT 144.742 0.000 145.022 0.720 ;
  LAYER ME1 ;
  RECT 144.742 0.000 145.022 0.720 ;
 END
 ANTENNAPARTIALMETALAREA                  0.805 LAYER ME1 ;
 ANTENNAGATEAREA                          0.072 LAYER ME1 ;
 ANTENNAGATEAREA                          0.072 LAYER ME2 ;
 ANTENNAGATEAREA                          0.072 LAYER ME3 ;
 ANTENNAGATEAREA                          0.072 LAYER ME4 ;
 ANTENNADIFFAREA                          0.218 LAYER ME1 ;
 ANTENNADIFFAREA                          0.218 LAYER ME2 ;
 ANTENNADIFFAREA                          0.218 LAYER ME3 ;
 ANTENNADIFFAREA                          0.218 LAYER ME4 ;
 ANTENNAMAXAREACAR                       13.984 LAYER ME1 ;
 ANTENNAMAXAREACAR                       16.784 LAYER ME2 ;
 ANTENNAMAXAREACAR                       19.584 LAYER ME3 ;
 ANTENNAMAXAREACAR                       22.384 LAYER ME4 ;
END DI17
PIN DO17
  DIRECTION OUTPUT ;
 PORT
  LAYER ME4 ;
  RECT 142.764 0.000 143.044 0.720 ;
  LAYER ME3 ;
  RECT 142.764 0.000 143.044 0.720 ;
  LAYER ME2 ;
  RECT 142.764 0.000 143.044 0.720 ;
  LAYER ME1 ;
  RECT 142.764 0.000 143.044 0.720 ;
 END
 ANTENNAPARTIALMETALAREA                  2.030 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME3 ;
 ANTENNADIFFAREA                          1.293 LAYER ME4 ;
END DO17
PIN DI16
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 136.734 0.000 137.014 0.720 ;
  LAYER ME3 ;
  RECT 136.734 0.000 137.014 0.720 ;
  LAYER ME2 ;
  RECT 136.734 0.000 137.014 0.720 ;
  LAYER ME1 ;
  RECT 136.734 0.000 137.014 0.720 ;
 END
 ANTENNAPARTIALMETALAREA                  0.805 LAYER ME1 ;
 ANTENNAGATEAREA                          0.072 LAYER ME1 ;
 ANTENNAGATEAREA                          0.072 LAYER ME2 ;
 ANTENNAGATEAREA                          0.072 LAYER ME3 ;
 ANTENNAGATEAREA                          0.072 LAYER ME4 ;
 ANTENNADIFFAREA                          0.218 LAYER ME1 ;
 ANTENNADIFFAREA                          0.218 LAYER ME2 ;
 ANTENNADIFFAREA                          0.218 LAYER ME3 ;
 ANTENNADIFFAREA                          0.218 LAYER ME4 ;
 ANTENNAMAXAREACAR                       13.984 LAYER ME1 ;
 ANTENNAMAXAREACAR                       16.784 LAYER ME2 ;
 ANTENNAMAXAREACAR                       19.584 LAYER ME3 ;
 ANTENNAMAXAREACAR                       22.384 LAYER ME4 ;
END DI16
PIN DO16
  DIRECTION OUTPUT ;
 PORT
  LAYER ME4 ;
  RECT 134.756 0.000 135.036 0.720 ;
  LAYER ME3 ;
  RECT 134.756 0.000 135.036 0.720 ;
  LAYER ME2 ;
  RECT 134.756 0.000 135.036 0.720 ;
  LAYER ME1 ;
  RECT 134.756 0.000 135.036 0.720 ;
 END
 ANTENNAPARTIALMETALAREA                  2.030 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME3 ;
 ANTENNADIFFAREA                          1.293 LAYER ME4 ;
END DO16
PIN DI15
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 128.726 0.000 129.006 0.720 ;
  LAYER ME3 ;
  RECT 128.726 0.000 129.006 0.720 ;
  LAYER ME2 ;
  RECT 128.726 0.000 129.006 0.720 ;
  LAYER ME1 ;
  RECT 128.726 0.000 129.006 0.720 ;
 END
 ANTENNAPARTIALMETALAREA                  0.805 LAYER ME1 ;
 ANTENNAGATEAREA                          0.072 LAYER ME1 ;
 ANTENNAGATEAREA                          0.072 LAYER ME2 ;
 ANTENNAGATEAREA                          0.072 LAYER ME3 ;
 ANTENNAGATEAREA                          0.072 LAYER ME4 ;
 ANTENNADIFFAREA                          0.218 LAYER ME1 ;
 ANTENNADIFFAREA                          0.218 LAYER ME2 ;
 ANTENNADIFFAREA                          0.218 LAYER ME3 ;
 ANTENNADIFFAREA                          0.218 LAYER ME4 ;
 ANTENNAMAXAREACAR                       13.984 LAYER ME1 ;
 ANTENNAMAXAREACAR                       16.784 LAYER ME2 ;
 ANTENNAMAXAREACAR                       19.584 LAYER ME3 ;
 ANTENNAMAXAREACAR                       22.384 LAYER ME4 ;
END DI15
PIN DO15
  DIRECTION OUTPUT ;
 PORT
  LAYER ME4 ;
  RECT 126.748 0.000 127.028 0.720 ;
  LAYER ME3 ;
  RECT 126.748 0.000 127.028 0.720 ;
  LAYER ME2 ;
  RECT 126.748 0.000 127.028 0.720 ;
  LAYER ME1 ;
  RECT 126.748 0.000 127.028 0.720 ;
 END
 ANTENNAPARTIALMETALAREA                  2.030 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME3 ;
 ANTENNADIFFAREA                          1.293 LAYER ME4 ;
END DO15
PIN DI14
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 120.718 0.000 120.998 0.720 ;
  LAYER ME3 ;
  RECT 120.718 0.000 120.998 0.720 ;
  LAYER ME2 ;
  RECT 120.718 0.000 120.998 0.720 ;
  LAYER ME1 ;
  RECT 120.718 0.000 120.998 0.720 ;
 END
 ANTENNAPARTIALMETALAREA                  0.522 LAYER ME1 ;
 ANTENNAGATEAREA                          0.072 LAYER ME1 ;
 ANTENNAGATEAREA                          0.072 LAYER ME2 ;
 ANTENNAGATEAREA                          0.072 LAYER ME3 ;
 ANTENNAGATEAREA                          0.072 LAYER ME4 ;
 ANTENNADIFFAREA                          0.218 LAYER ME1 ;
 ANTENNADIFFAREA                          0.218 LAYER ME2 ;
 ANTENNADIFFAREA                          0.218 LAYER ME3 ;
 ANTENNADIFFAREA                          0.218 LAYER ME4 ;
 ANTENNAMAXAREACAR                       10.048 LAYER ME1 ;
 ANTENNAMAXAREACAR                       12.848 LAYER ME2 ;
 ANTENNAMAXAREACAR                       15.648 LAYER ME3 ;
 ANTENNAMAXAREACAR                       18.448 LAYER ME4 ;
END DI14
PIN DO14
  DIRECTION OUTPUT ;
 PORT
  LAYER ME4 ;
  RECT 118.660 0.000 118.940 0.720 ;
  LAYER ME3 ;
  RECT 118.660 0.000 118.940 0.720 ;
  LAYER ME2 ;
  RECT 118.660 0.000 118.940 0.720 ;
  LAYER ME1 ;
  RECT 118.660 0.000 118.940 0.720 ;
 END
 ANTENNAPARTIALMETALAREA                  2.030 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME3 ;
 ANTENNADIFFAREA                          1.293 LAYER ME4 ;
END DO14
PIN WEB2
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 119.140 0.000 119.420 0.720 ;
  LAYER ME3 ;
  RECT 119.140 0.000 119.420 0.720 ;
  LAYER ME2 ;
  RECT 119.140 0.000 119.420 0.720 ;
  LAYER ME1 ;
  RECT 119.140 0.000 119.420 0.720 ;
 END
 ANTENNAPARTIALMETALAREA                  0.436 LAYER ME2 ;
 ANTENNAGATEAREA                          0.288 LAYER ME2 ;
 ANTENNAGATEAREA                          0.288 LAYER ME3 ;
 ANTENNAGATEAREA                          0.288 LAYER ME4 ;
 ANTENNADIFFAREA                          0.218 LAYER ME2 ;
 ANTENNADIFFAREA                          0.218 LAYER ME3 ;
 ANTENNADIFFAREA                          0.218 LAYER ME4 ;
 ANTENNAMAXAREACAR                        4.602 LAYER ME2 ;
 ANTENNAMAXAREACAR                        5.302 LAYER ME3 ;
 ANTENNAMAXAREACAR                        6.002 LAYER ME4 ;
END WEB2
PIN DI13
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 112.710 0.000 112.990 0.720 ;
  LAYER ME3 ;
  RECT 112.710 0.000 112.990 0.720 ;
  LAYER ME2 ;
  RECT 112.710 0.000 112.990 0.720 ;
  LAYER ME1 ;
  RECT 112.710 0.000 112.990 0.720 ;
 END
 ANTENNAPARTIALMETALAREA                  0.805 LAYER ME1 ;
 ANTENNAGATEAREA                          0.072 LAYER ME1 ;
 ANTENNAGATEAREA                          0.072 LAYER ME2 ;
 ANTENNAGATEAREA                          0.072 LAYER ME3 ;
 ANTENNAGATEAREA                          0.072 LAYER ME4 ;
 ANTENNADIFFAREA                          0.218 LAYER ME1 ;
 ANTENNADIFFAREA                          0.218 LAYER ME2 ;
 ANTENNADIFFAREA                          0.218 LAYER ME3 ;
 ANTENNADIFFAREA                          0.218 LAYER ME4 ;
 ANTENNAMAXAREACAR                       13.984 LAYER ME1 ;
 ANTENNAMAXAREACAR                       16.784 LAYER ME2 ;
 ANTENNAMAXAREACAR                       19.584 LAYER ME3 ;
 ANTENNAMAXAREACAR                       22.384 LAYER ME4 ;
END DI13
PIN DO13
  DIRECTION OUTPUT ;
 PORT
  LAYER ME4 ;
  RECT 110.732 0.000 111.012 0.720 ;
  LAYER ME3 ;
  RECT 110.732 0.000 111.012 0.720 ;
  LAYER ME2 ;
  RECT 110.732 0.000 111.012 0.720 ;
  LAYER ME1 ;
  RECT 110.732 0.000 111.012 0.720 ;
 END
 ANTENNAPARTIALMETALAREA                  2.030 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME3 ;
 ANTENNADIFFAREA                          1.293 LAYER ME4 ;
END DO13
PIN DI12
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 104.702 0.000 104.982 0.720 ;
  LAYER ME3 ;
  RECT 104.702 0.000 104.982 0.720 ;
  LAYER ME2 ;
  RECT 104.702 0.000 104.982 0.720 ;
  LAYER ME1 ;
  RECT 104.702 0.000 104.982 0.720 ;
 END
 ANTENNAPARTIALMETALAREA                  0.805 LAYER ME1 ;
 ANTENNAGATEAREA                          0.072 LAYER ME1 ;
 ANTENNAGATEAREA                          0.072 LAYER ME2 ;
 ANTENNAGATEAREA                          0.072 LAYER ME3 ;
 ANTENNAGATEAREA                          0.072 LAYER ME4 ;
 ANTENNADIFFAREA                          0.218 LAYER ME1 ;
 ANTENNADIFFAREA                          0.218 LAYER ME2 ;
 ANTENNADIFFAREA                          0.218 LAYER ME3 ;
 ANTENNADIFFAREA                          0.218 LAYER ME4 ;
 ANTENNAMAXAREACAR                       13.984 LAYER ME1 ;
 ANTENNAMAXAREACAR                       16.784 LAYER ME2 ;
 ANTENNAMAXAREACAR                       19.584 LAYER ME3 ;
 ANTENNAMAXAREACAR                       22.384 LAYER ME4 ;
END DI12
PIN DO12
  DIRECTION OUTPUT ;
 PORT
  LAYER ME4 ;
  RECT 102.724 0.000 103.004 0.720 ;
  LAYER ME3 ;
  RECT 102.724 0.000 103.004 0.720 ;
  LAYER ME2 ;
  RECT 102.724 0.000 103.004 0.720 ;
  LAYER ME1 ;
  RECT 102.724 0.000 103.004 0.720 ;
 END
 ANTENNAPARTIALMETALAREA                  2.030 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME3 ;
 ANTENNADIFFAREA                          1.293 LAYER ME4 ;
END DO12
PIN DI11
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 96.694 0.000 96.974 0.720 ;
  LAYER ME3 ;
  RECT 96.694 0.000 96.974 0.720 ;
  LAYER ME2 ;
  RECT 96.694 0.000 96.974 0.720 ;
  LAYER ME1 ;
  RECT 96.694 0.000 96.974 0.720 ;
 END
 ANTENNAPARTIALMETALAREA                  0.805 LAYER ME1 ;
 ANTENNAGATEAREA                          0.072 LAYER ME1 ;
 ANTENNAGATEAREA                          0.072 LAYER ME2 ;
 ANTENNAGATEAREA                          0.072 LAYER ME3 ;
 ANTENNAGATEAREA                          0.072 LAYER ME4 ;
 ANTENNADIFFAREA                          0.218 LAYER ME1 ;
 ANTENNADIFFAREA                          0.218 LAYER ME2 ;
 ANTENNADIFFAREA                          0.218 LAYER ME3 ;
 ANTENNADIFFAREA                          0.218 LAYER ME4 ;
 ANTENNAMAXAREACAR                       13.984 LAYER ME1 ;
 ANTENNAMAXAREACAR                       16.784 LAYER ME2 ;
 ANTENNAMAXAREACAR                       19.584 LAYER ME3 ;
 ANTENNAMAXAREACAR                       22.384 LAYER ME4 ;
END DI11
PIN DO11
  DIRECTION OUTPUT ;
 PORT
  LAYER ME4 ;
  RECT 94.716 0.000 94.996 0.720 ;
  LAYER ME3 ;
  RECT 94.716 0.000 94.996 0.720 ;
  LAYER ME2 ;
  RECT 94.716 0.000 94.996 0.720 ;
  LAYER ME1 ;
  RECT 94.716 0.000 94.996 0.720 ;
 END
 ANTENNAPARTIALMETALAREA                  2.030 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME3 ;
 ANTENNADIFFAREA                          1.293 LAYER ME4 ;
END DO11
PIN DI10
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 88.686 0.000 88.966 0.720 ;
  LAYER ME3 ;
  RECT 88.686 0.000 88.966 0.720 ;
  LAYER ME2 ;
  RECT 88.686 0.000 88.966 0.720 ;
  LAYER ME1 ;
  RECT 88.686 0.000 88.966 0.720 ;
 END
 ANTENNAPARTIALMETALAREA                  0.805 LAYER ME1 ;
 ANTENNAGATEAREA                          0.072 LAYER ME1 ;
 ANTENNAGATEAREA                          0.072 LAYER ME2 ;
 ANTENNAGATEAREA                          0.072 LAYER ME3 ;
 ANTENNAGATEAREA                          0.072 LAYER ME4 ;
 ANTENNADIFFAREA                          0.218 LAYER ME1 ;
 ANTENNADIFFAREA                          0.218 LAYER ME2 ;
 ANTENNADIFFAREA                          0.218 LAYER ME3 ;
 ANTENNADIFFAREA                          0.218 LAYER ME4 ;
 ANTENNAMAXAREACAR                       13.984 LAYER ME1 ;
 ANTENNAMAXAREACAR                       16.784 LAYER ME2 ;
 ANTENNAMAXAREACAR                       19.584 LAYER ME3 ;
 ANTENNAMAXAREACAR                       22.384 LAYER ME4 ;
END DI10
PIN DO10
  DIRECTION OUTPUT ;
 PORT
  LAYER ME4 ;
  RECT 86.708 0.000 86.988 0.720 ;
  LAYER ME3 ;
  RECT 86.708 0.000 86.988 0.720 ;
  LAYER ME2 ;
  RECT 86.708 0.000 86.988 0.720 ;
  LAYER ME1 ;
  RECT 86.708 0.000 86.988 0.720 ;
 END
 ANTENNAPARTIALMETALAREA                  2.030 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME3 ;
 ANTENNADIFFAREA                          1.293 LAYER ME4 ;
END DO10
PIN DI9
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 80.678 0.000 80.958 0.720 ;
  LAYER ME3 ;
  RECT 80.678 0.000 80.958 0.720 ;
  LAYER ME2 ;
  RECT 80.678 0.000 80.958 0.720 ;
  LAYER ME1 ;
  RECT 80.678 0.000 80.958 0.720 ;
 END
 ANTENNAPARTIALMETALAREA                  0.805 LAYER ME1 ;
 ANTENNAGATEAREA                          0.072 LAYER ME1 ;
 ANTENNAGATEAREA                          0.072 LAYER ME2 ;
 ANTENNAGATEAREA                          0.072 LAYER ME3 ;
 ANTENNAGATEAREA                          0.072 LAYER ME4 ;
 ANTENNADIFFAREA                          0.218 LAYER ME1 ;
 ANTENNADIFFAREA                          0.218 LAYER ME2 ;
 ANTENNADIFFAREA                          0.218 LAYER ME3 ;
 ANTENNADIFFAREA                          0.218 LAYER ME4 ;
 ANTENNAMAXAREACAR                       13.984 LAYER ME1 ;
 ANTENNAMAXAREACAR                       16.784 LAYER ME2 ;
 ANTENNAMAXAREACAR                       19.584 LAYER ME3 ;
 ANTENNAMAXAREACAR                       22.384 LAYER ME4 ;
END DI9
PIN DO9
  DIRECTION OUTPUT ;
 PORT
  LAYER ME4 ;
  RECT 78.700 0.000 78.980 0.720 ;
  LAYER ME3 ;
  RECT 78.700 0.000 78.980 0.720 ;
  LAYER ME2 ;
  RECT 78.700 0.000 78.980 0.720 ;
  LAYER ME1 ;
  RECT 78.700 0.000 78.980 0.720 ;
 END
 ANTENNAPARTIALMETALAREA                  2.030 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME3 ;
 ANTENNADIFFAREA                          1.293 LAYER ME4 ;
END DO9
PIN DI8
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 72.670 0.000 72.950 0.720 ;
  LAYER ME3 ;
  RECT 72.670 0.000 72.950 0.720 ;
  LAYER ME2 ;
  RECT 72.670 0.000 72.950 0.720 ;
  LAYER ME1 ;
  RECT 72.670 0.000 72.950 0.720 ;
 END
 ANTENNAPARTIALMETALAREA                  0.805 LAYER ME1 ;
 ANTENNAGATEAREA                          0.072 LAYER ME1 ;
 ANTENNAGATEAREA                          0.072 LAYER ME2 ;
 ANTENNAGATEAREA                          0.072 LAYER ME3 ;
 ANTENNAGATEAREA                          0.072 LAYER ME4 ;
 ANTENNADIFFAREA                          0.218 LAYER ME1 ;
 ANTENNADIFFAREA                          0.218 LAYER ME2 ;
 ANTENNADIFFAREA                          0.218 LAYER ME3 ;
 ANTENNADIFFAREA                          0.218 LAYER ME4 ;
 ANTENNAMAXAREACAR                       13.984 LAYER ME1 ;
 ANTENNAMAXAREACAR                       16.784 LAYER ME2 ;
 ANTENNAMAXAREACAR                       19.584 LAYER ME3 ;
 ANTENNAMAXAREACAR                       22.384 LAYER ME4 ;
END DI8
PIN DO8
  DIRECTION OUTPUT ;
 PORT
  LAYER ME4 ;
  RECT 70.692 0.000 70.972 0.720 ;
  LAYER ME3 ;
  RECT 70.692 0.000 70.972 0.720 ;
  LAYER ME2 ;
  RECT 70.692 0.000 70.972 0.720 ;
  LAYER ME1 ;
  RECT 70.692 0.000 70.972 0.720 ;
 END
 ANTENNAPARTIALMETALAREA                  2.030 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME3 ;
 ANTENNADIFFAREA                          1.293 LAYER ME4 ;
END DO8
PIN DI7
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 64.662 0.000 64.942 0.720 ;
  LAYER ME3 ;
  RECT 64.662 0.000 64.942 0.720 ;
  LAYER ME2 ;
  RECT 64.662 0.000 64.942 0.720 ;
  LAYER ME1 ;
  RECT 64.662 0.000 64.942 0.720 ;
 END
 ANTENNAPARTIALMETALAREA                  0.522 LAYER ME1 ;
 ANTENNAGATEAREA                          0.072 LAYER ME1 ;
 ANTENNAGATEAREA                          0.072 LAYER ME2 ;
 ANTENNAGATEAREA                          0.072 LAYER ME3 ;
 ANTENNAGATEAREA                          0.072 LAYER ME4 ;
 ANTENNADIFFAREA                          0.218 LAYER ME1 ;
 ANTENNADIFFAREA                          0.218 LAYER ME2 ;
 ANTENNADIFFAREA                          0.218 LAYER ME3 ;
 ANTENNADIFFAREA                          0.218 LAYER ME4 ;
 ANTENNAMAXAREACAR                       10.048 LAYER ME1 ;
 ANTENNAMAXAREACAR                       12.848 LAYER ME2 ;
 ANTENNAMAXAREACAR                       15.648 LAYER ME3 ;
 ANTENNAMAXAREACAR                       18.448 LAYER ME4 ;
END DI7
PIN DO7
  DIRECTION OUTPUT ;
 PORT
  LAYER ME4 ;
  RECT 62.604 0.000 62.884 0.720 ;
  LAYER ME3 ;
  RECT 62.604 0.000 62.884 0.720 ;
  LAYER ME2 ;
  RECT 62.604 0.000 62.884 0.720 ;
  LAYER ME1 ;
  RECT 62.604 0.000 62.884 0.720 ;
 END
 ANTENNAPARTIALMETALAREA                  2.030 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME3 ;
 ANTENNADIFFAREA                          1.293 LAYER ME4 ;
END DO7
PIN WEB1
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 63.084 0.000 63.364 0.720 ;
  LAYER ME3 ;
  RECT 63.084 0.000 63.364 0.720 ;
  LAYER ME2 ;
  RECT 63.084 0.000 63.364 0.720 ;
  LAYER ME1 ;
  RECT 63.084 0.000 63.364 0.720 ;
 END
 ANTENNAPARTIALMETALAREA                  0.436 LAYER ME2 ;
 ANTENNAGATEAREA                          0.288 LAYER ME2 ;
 ANTENNAGATEAREA                          0.288 LAYER ME3 ;
 ANTENNAGATEAREA                          0.288 LAYER ME4 ;
 ANTENNADIFFAREA                          0.218 LAYER ME2 ;
 ANTENNADIFFAREA                          0.218 LAYER ME3 ;
 ANTENNADIFFAREA                          0.218 LAYER ME4 ;
 ANTENNAMAXAREACAR                        4.602 LAYER ME2 ;
 ANTENNAMAXAREACAR                        5.302 LAYER ME3 ;
 ANTENNAMAXAREACAR                        6.002 LAYER ME4 ;
END WEB1
PIN DI6
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 56.654 0.000 56.934 0.720 ;
  LAYER ME3 ;
  RECT 56.654 0.000 56.934 0.720 ;
  LAYER ME2 ;
  RECT 56.654 0.000 56.934 0.720 ;
  LAYER ME1 ;
  RECT 56.654 0.000 56.934 0.720 ;
 END
 ANTENNAPARTIALMETALAREA                  0.805 LAYER ME1 ;
 ANTENNAGATEAREA                          0.072 LAYER ME1 ;
 ANTENNAGATEAREA                          0.072 LAYER ME2 ;
 ANTENNAGATEAREA                          0.072 LAYER ME3 ;
 ANTENNAGATEAREA                          0.072 LAYER ME4 ;
 ANTENNADIFFAREA                          0.218 LAYER ME1 ;
 ANTENNADIFFAREA                          0.218 LAYER ME2 ;
 ANTENNADIFFAREA                          0.218 LAYER ME3 ;
 ANTENNADIFFAREA                          0.218 LAYER ME4 ;
 ANTENNAMAXAREACAR                       13.984 LAYER ME1 ;
 ANTENNAMAXAREACAR                       16.784 LAYER ME2 ;
 ANTENNAMAXAREACAR                       19.584 LAYER ME3 ;
 ANTENNAMAXAREACAR                       22.384 LAYER ME4 ;
END DI6
PIN DO6
  DIRECTION OUTPUT ;
 PORT
  LAYER ME4 ;
  RECT 54.676 0.000 54.956 0.720 ;
  LAYER ME3 ;
  RECT 54.676 0.000 54.956 0.720 ;
  LAYER ME2 ;
  RECT 54.676 0.000 54.956 0.720 ;
  LAYER ME1 ;
  RECT 54.676 0.000 54.956 0.720 ;
 END
 ANTENNAPARTIALMETALAREA                  2.030 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME3 ;
 ANTENNADIFFAREA                          1.293 LAYER ME4 ;
END DO6
PIN DI5
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 48.646 0.000 48.926 0.720 ;
  LAYER ME3 ;
  RECT 48.646 0.000 48.926 0.720 ;
  LAYER ME2 ;
  RECT 48.646 0.000 48.926 0.720 ;
  LAYER ME1 ;
  RECT 48.646 0.000 48.926 0.720 ;
 END
 ANTENNAPARTIALMETALAREA                  0.805 LAYER ME1 ;
 ANTENNAGATEAREA                          0.072 LAYER ME1 ;
 ANTENNAGATEAREA                          0.072 LAYER ME2 ;
 ANTENNAGATEAREA                          0.072 LAYER ME3 ;
 ANTENNAGATEAREA                          0.072 LAYER ME4 ;
 ANTENNADIFFAREA                          0.218 LAYER ME1 ;
 ANTENNADIFFAREA                          0.218 LAYER ME2 ;
 ANTENNADIFFAREA                          0.218 LAYER ME3 ;
 ANTENNADIFFAREA                          0.218 LAYER ME4 ;
 ANTENNAMAXAREACAR                       13.984 LAYER ME1 ;
 ANTENNAMAXAREACAR                       16.784 LAYER ME2 ;
 ANTENNAMAXAREACAR                       19.584 LAYER ME3 ;
 ANTENNAMAXAREACAR                       22.384 LAYER ME4 ;
END DI5
PIN DO5
  DIRECTION OUTPUT ;
 PORT
  LAYER ME4 ;
  RECT 46.668 0.000 46.948 0.720 ;
  LAYER ME3 ;
  RECT 46.668 0.000 46.948 0.720 ;
  LAYER ME2 ;
  RECT 46.668 0.000 46.948 0.720 ;
  LAYER ME1 ;
  RECT 46.668 0.000 46.948 0.720 ;
 END
 ANTENNAPARTIALMETALAREA                  2.030 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME3 ;
 ANTENNADIFFAREA                          1.293 LAYER ME4 ;
END DO5
PIN DI4
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 40.638 0.000 40.918 0.720 ;
  LAYER ME3 ;
  RECT 40.638 0.000 40.918 0.720 ;
  LAYER ME2 ;
  RECT 40.638 0.000 40.918 0.720 ;
  LAYER ME1 ;
  RECT 40.638 0.000 40.918 0.720 ;
 END
 ANTENNAPARTIALMETALAREA                  0.805 LAYER ME1 ;
 ANTENNAGATEAREA                          0.072 LAYER ME1 ;
 ANTENNAGATEAREA                          0.072 LAYER ME2 ;
 ANTENNAGATEAREA                          0.072 LAYER ME3 ;
 ANTENNAGATEAREA                          0.072 LAYER ME4 ;
 ANTENNADIFFAREA                          0.218 LAYER ME1 ;
 ANTENNADIFFAREA                          0.218 LAYER ME2 ;
 ANTENNADIFFAREA                          0.218 LAYER ME3 ;
 ANTENNADIFFAREA                          0.218 LAYER ME4 ;
 ANTENNAMAXAREACAR                       13.984 LAYER ME1 ;
 ANTENNAMAXAREACAR                       16.784 LAYER ME2 ;
 ANTENNAMAXAREACAR                       19.584 LAYER ME3 ;
 ANTENNAMAXAREACAR                       22.384 LAYER ME4 ;
END DI4
PIN DO4
  DIRECTION OUTPUT ;
 PORT
  LAYER ME4 ;
  RECT 38.660 0.000 38.940 0.720 ;
  LAYER ME3 ;
  RECT 38.660 0.000 38.940 0.720 ;
  LAYER ME2 ;
  RECT 38.660 0.000 38.940 0.720 ;
  LAYER ME1 ;
  RECT 38.660 0.000 38.940 0.720 ;
 END
 ANTENNAPARTIALMETALAREA                  2.030 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME3 ;
 ANTENNADIFFAREA                          1.293 LAYER ME4 ;
END DO4
PIN DI3
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 32.630 0.000 32.910 0.720 ;
  LAYER ME3 ;
  RECT 32.630 0.000 32.910 0.720 ;
  LAYER ME2 ;
  RECT 32.630 0.000 32.910 0.720 ;
  LAYER ME1 ;
  RECT 32.630 0.000 32.910 0.720 ;
 END
 ANTENNAPARTIALMETALAREA                  0.805 LAYER ME1 ;
 ANTENNAGATEAREA                          0.072 LAYER ME1 ;
 ANTENNAGATEAREA                          0.072 LAYER ME2 ;
 ANTENNAGATEAREA                          0.072 LAYER ME3 ;
 ANTENNAGATEAREA                          0.072 LAYER ME4 ;
 ANTENNADIFFAREA                          0.218 LAYER ME1 ;
 ANTENNADIFFAREA                          0.218 LAYER ME2 ;
 ANTENNADIFFAREA                          0.218 LAYER ME3 ;
 ANTENNADIFFAREA                          0.218 LAYER ME4 ;
 ANTENNAMAXAREACAR                       13.984 LAYER ME1 ;
 ANTENNAMAXAREACAR                       16.784 LAYER ME2 ;
 ANTENNAMAXAREACAR                       19.584 LAYER ME3 ;
 ANTENNAMAXAREACAR                       22.384 LAYER ME4 ;
END DI3
PIN DO3
  DIRECTION OUTPUT ;
 PORT
  LAYER ME4 ;
  RECT 30.652 0.000 30.932 0.720 ;
  LAYER ME3 ;
  RECT 30.652 0.000 30.932 0.720 ;
  LAYER ME2 ;
  RECT 30.652 0.000 30.932 0.720 ;
  LAYER ME1 ;
  RECT 30.652 0.000 30.932 0.720 ;
 END
 ANTENNAPARTIALMETALAREA                  2.030 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME3 ;
 ANTENNADIFFAREA                          1.293 LAYER ME4 ;
END DO3
PIN DI2
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 24.622 0.000 24.902 0.720 ;
  LAYER ME3 ;
  RECT 24.622 0.000 24.902 0.720 ;
  LAYER ME2 ;
  RECT 24.622 0.000 24.902 0.720 ;
  LAYER ME1 ;
  RECT 24.622 0.000 24.902 0.720 ;
 END
 ANTENNAPARTIALMETALAREA                  0.805 LAYER ME1 ;
 ANTENNAGATEAREA                          0.072 LAYER ME1 ;
 ANTENNAGATEAREA                          0.072 LAYER ME2 ;
 ANTENNAGATEAREA                          0.072 LAYER ME3 ;
 ANTENNAGATEAREA                          0.072 LAYER ME4 ;
 ANTENNADIFFAREA                          0.218 LAYER ME1 ;
 ANTENNADIFFAREA                          0.218 LAYER ME2 ;
 ANTENNADIFFAREA                          0.218 LAYER ME3 ;
 ANTENNADIFFAREA                          0.218 LAYER ME4 ;
 ANTENNAMAXAREACAR                       13.984 LAYER ME1 ;
 ANTENNAMAXAREACAR                       16.784 LAYER ME2 ;
 ANTENNAMAXAREACAR                       19.584 LAYER ME3 ;
 ANTENNAMAXAREACAR                       22.384 LAYER ME4 ;
END DI2
PIN DO2
  DIRECTION OUTPUT ;
 PORT
  LAYER ME4 ;
  RECT 22.644 0.000 22.924 0.720 ;
  LAYER ME3 ;
  RECT 22.644 0.000 22.924 0.720 ;
  LAYER ME2 ;
  RECT 22.644 0.000 22.924 0.720 ;
  LAYER ME1 ;
  RECT 22.644 0.000 22.924 0.720 ;
 END
 ANTENNAPARTIALMETALAREA                  2.030 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME3 ;
 ANTENNADIFFAREA                          1.293 LAYER ME4 ;
END DO2
PIN DI1
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 16.614 0.000 16.894 0.720 ;
  LAYER ME3 ;
  RECT 16.614 0.000 16.894 0.720 ;
  LAYER ME2 ;
  RECT 16.614 0.000 16.894 0.720 ;
  LAYER ME1 ;
  RECT 16.614 0.000 16.894 0.720 ;
 END
 ANTENNAPARTIALMETALAREA                  0.805 LAYER ME1 ;
 ANTENNAGATEAREA                          0.072 LAYER ME1 ;
 ANTENNAGATEAREA                          0.072 LAYER ME2 ;
 ANTENNAGATEAREA                          0.072 LAYER ME3 ;
 ANTENNAGATEAREA                          0.072 LAYER ME4 ;
 ANTENNADIFFAREA                          0.218 LAYER ME1 ;
 ANTENNADIFFAREA                          0.218 LAYER ME2 ;
 ANTENNADIFFAREA                          0.218 LAYER ME3 ;
 ANTENNADIFFAREA                          0.218 LAYER ME4 ;
 ANTENNAMAXAREACAR                       13.984 LAYER ME1 ;
 ANTENNAMAXAREACAR                       16.784 LAYER ME2 ;
 ANTENNAMAXAREACAR                       19.584 LAYER ME3 ;
 ANTENNAMAXAREACAR                       22.384 LAYER ME4 ;
END DI1
PIN DO1
  DIRECTION OUTPUT ;
 PORT
  LAYER ME4 ;
  RECT 14.636 0.000 14.916 0.720 ;
  LAYER ME3 ;
  RECT 14.636 0.000 14.916 0.720 ;
  LAYER ME2 ;
  RECT 14.636 0.000 14.916 0.720 ;
  LAYER ME1 ;
  RECT 14.636 0.000 14.916 0.720 ;
 END
 ANTENNAPARTIALMETALAREA                  2.030 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME3 ;
 ANTENNADIFFAREA                          1.293 LAYER ME4 ;
END DO1
PIN DI0
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 8.606 0.000 8.886 0.720 ;
  LAYER ME3 ;
  RECT 8.606 0.000 8.886 0.720 ;
  LAYER ME2 ;
  RECT 8.606 0.000 8.886 0.720 ;
  LAYER ME1 ;
  RECT 8.606 0.000 8.886 0.720 ;
 END
 ANTENNAPARTIALMETALAREA                  0.522 LAYER ME1 ;
 ANTENNAGATEAREA                          0.072 LAYER ME1 ;
 ANTENNAGATEAREA                          0.072 LAYER ME2 ;
 ANTENNAGATEAREA                          0.072 LAYER ME3 ;
 ANTENNAGATEAREA                          0.072 LAYER ME4 ;
 ANTENNADIFFAREA                          0.218 LAYER ME1 ;
 ANTENNADIFFAREA                          0.218 LAYER ME2 ;
 ANTENNADIFFAREA                          0.218 LAYER ME3 ;
 ANTENNADIFFAREA                          0.218 LAYER ME4 ;
 ANTENNAMAXAREACAR                       10.048 LAYER ME1 ;
 ANTENNAMAXAREACAR                       12.848 LAYER ME2 ;
 ANTENNAMAXAREACAR                       15.648 LAYER ME3 ;
 ANTENNAMAXAREACAR                       18.448 LAYER ME4 ;
END DI0
PIN DO0
  DIRECTION OUTPUT ;
 PORT
  LAYER ME4 ;
  RECT 6.548 0.000 6.828 0.720 ;
  LAYER ME3 ;
  RECT 6.548 0.000 6.828 0.720 ;
  LAYER ME2 ;
  RECT 6.548 0.000 6.828 0.720 ;
  LAYER ME1 ;
  RECT 6.548 0.000 6.828 0.720 ;
 END
 ANTENNAPARTIALMETALAREA                  2.030 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME3 ;
 ANTENNADIFFAREA                          1.293 LAYER ME4 ;
END DO0
PIN WEB0
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 7.028 0.000 7.308 0.720 ;
  LAYER ME3 ;
  RECT 7.028 0.000 7.308 0.720 ;
  LAYER ME2 ;
  RECT 7.028 0.000 7.308 0.720 ;
  LAYER ME1 ;
  RECT 7.028 0.000 7.308 0.720 ;
 END
 ANTENNAPARTIALMETALAREA                  0.436 LAYER ME2 ;
 ANTENNAGATEAREA                          0.288 LAYER ME2 ;
 ANTENNAGATEAREA                          0.288 LAYER ME3 ;
 ANTENNAGATEAREA                          0.288 LAYER ME4 ;
 ANTENNADIFFAREA                          0.218 LAYER ME2 ;
 ANTENNADIFFAREA                          0.218 LAYER ME3 ;
 ANTENNADIFFAREA                          0.218 LAYER ME4 ;
 ANTENNAMAXAREACAR                        4.602 LAYER ME2 ;
 ANTENNAMAXAREACAR                        5.302 LAYER ME3 ;
 ANTENNAMAXAREACAR                        6.002 LAYER ME4 ;
END WEB0
PIN A2
  DIRECTION INPUT ;
 PORT
  LAYER ME3 ;
  RECT 187.052 0.000 187.372 0.600 ;
  LAYER ME2 ;
  RECT 187.052 0.000 187.372 0.600 ;
  LAYER ME1 ;
  RECT 187.052 0.000 187.372 0.600 ;
 END
 ANTENNAPARTIALMETALAREA                  1.067 LAYER ME2 ;
 ANTENNAGATEAREA                          0.144 LAYER ME2 ;
 ANTENNAGATEAREA                          0.144 LAYER ME3 ;
 ANTENNADIFFAREA                          0.218 LAYER ME2 ;
 ANTENNADIFFAREA                          0.218 LAYER ME3 ;
 ANTENNAMAXAREACAR                        9.746 LAYER ME2 ;
 ANTENNAMAXAREACAR                       11.079 LAYER ME3 ;
END A2
PIN A3
  DIRECTION INPUT ;
 PORT
  LAYER ME3 ;
  RECT 187.639 0.000 187.959 0.600 ;
  LAYER ME2 ;
  RECT 187.639 0.000 187.959 0.600 ;
  LAYER ME1 ;
  RECT 187.639 0.000 187.959 0.600 ;
 END
 ANTENNAPARTIALMETALAREA                  1.188 LAYER ME2 ;
 ANTENNAGATEAREA                          0.144 LAYER ME2 ;
 ANTENNAGATEAREA                          0.144 LAYER ME3 ;
 ANTENNADIFFAREA                          0.218 LAYER ME2 ;
 ANTENNADIFFAREA                          0.218 LAYER ME3 ;
 ANTENNAMAXAREACAR                       10.582 LAYER ME2 ;
 ANTENNAMAXAREACAR                       11.915 LAYER ME3 ;
END A3
PIN A4
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 180.800 0.000 181.120 0.600 ;
  LAYER ME3 ;
  RECT 180.800 0.000 181.120 0.600 ;
  LAYER ME2 ;
  RECT 180.800 0.000 181.120 0.600 ;
  LAYER ME1 ;
  RECT 180.800 0.000 181.120 0.600 ;
 END
 ANTENNAPARTIALMETALAREA                  1.910 LAYER ME2 ;
 ANTENNAGATEAREA                          0.180 LAYER ME2 ;
 ANTENNAGATEAREA                          0.180 LAYER ME3 ;
 ANTENNAGATEAREA                          0.180 LAYER ME4 ;
 ANTENNADIFFAREA                          0.218 LAYER ME2 ;
 ANTENNADIFFAREA                          0.218 LAYER ME3 ;
 ANTENNADIFFAREA                          0.218 LAYER ME4 ;
 ANTENNAMAXAREACAR                       13.456 LAYER ME2 ;
 ANTENNAMAXAREACAR                       14.522 LAYER ME3 ;
 ANTENNAMAXAREACAR                       15.589 LAYER ME4 ;
END A4
PIN A5
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 180.180 0.000 180.500 0.600 ;
  LAYER ME3 ;
  RECT 180.180 0.000 180.500 0.600 ;
  LAYER ME2 ;
  RECT 180.180 0.000 180.500 0.600 ;
  LAYER ME1 ;
  RECT 180.180 0.000 180.500 0.600 ;
 END
 ANTENNAPARTIALMETALAREA                  1.447 LAYER ME2 ;
 ANTENNAGATEAREA                          0.180 LAYER ME2 ;
 ANTENNAGATEAREA                          0.180 LAYER ME3 ;
 ANTENNAGATEAREA                          0.180 LAYER ME4 ;
 ANTENNADIFFAREA                          0.218 LAYER ME2 ;
 ANTENNADIFFAREA                          0.218 LAYER ME3 ;
 ANTENNADIFFAREA                          0.218 LAYER ME4 ;
 ANTENNAMAXAREACAR                       12.818 LAYER ME2 ;
 ANTENNAMAXAREACAR                       13.884 LAYER ME3 ;
 ANTENNAMAXAREACAR                       14.951 LAYER ME4 ;
END A5
PIN A6
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 176.700 0.000 177.020 0.600 ;
  LAYER ME3 ;
  RECT 176.700 0.000 177.020 0.600 ;
  LAYER ME2 ;
  RECT 176.700 0.000 177.020 0.600 ;
  LAYER ME1 ;
  RECT 176.700 0.000 177.020 0.600 ;
 END
 ANTENNAPARTIALMETALAREA                  1.910 LAYER ME2 ;
 ANTENNAGATEAREA                          0.180 LAYER ME2 ;
 ANTENNAGATEAREA                          0.180 LAYER ME3 ;
 ANTENNAGATEAREA                          0.180 LAYER ME4 ;
 ANTENNADIFFAREA                          0.218 LAYER ME2 ;
 ANTENNADIFFAREA                          0.218 LAYER ME3 ;
 ANTENNADIFFAREA                          0.218 LAYER ME4 ;
 ANTENNAMAXAREACAR                       13.456 LAYER ME2 ;
 ANTENNAMAXAREACAR                       14.522 LAYER ME3 ;
 ANTENNAMAXAREACAR                       15.589 LAYER ME4 ;
END A6
PIN A1
  DIRECTION INPUT ;
 PORT
  LAYER ME3 ;
  RECT 191.925 0.000 192.245 0.712 ;
  LAYER ME2 ;
  RECT 191.925 0.000 192.245 0.712 ;
  LAYER ME1 ;
  RECT 191.925 0.000 192.245 0.712 ;
 END
 ANTENNAPARTIALMETALAREA                  3.219 LAYER ME2 ;
 ANTENNAGATEAREA                          0.108 LAYER ME2 ;
 ANTENNAGATEAREA                          0.108 LAYER ME3 ;
 ANTENNADIFFAREA                          0.218 LAYER ME2 ;
 ANTENNADIFFAREA                          0.218 LAYER ME3 ;
 ANTENNAMAXAREACAR                       33.245 LAYER ME2 ;
 ANTENNAMAXAREACAR                       35.355 LAYER ME3 ;
END A1
PIN A0
  DIRECTION INPUT ;
 PORT
  LAYER ME3 ;
  RECT 195.154 0.000 195.474 0.712 ;
  LAYER ME2 ;
  RECT 195.154 0.000 195.474 0.712 ;
  LAYER ME1 ;
  RECT 195.154 0.000 195.474 0.712 ;
 END
 ANTENNAPARTIALMETALAREA                  3.457 LAYER ME2 ;
 ANTENNAGATEAREA                          0.108 LAYER ME2 ;
 ANTENNAGATEAREA                          0.108 LAYER ME3 ;
 ANTENNADIFFAREA                          0.218 LAYER ME2 ;
 ANTENNADIFFAREA                          0.218 LAYER ME3 ;
 ANTENNAMAXAREACAR                       35.986 LAYER ME2 ;
 ANTENNAMAXAREACAR                       38.095 LAYER ME3 ;
END A0
PIN DVSE
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 207.745 0.000 208.065 0.717 ;
  LAYER ME3 ;
  RECT 207.745 0.000 208.065 0.717 ;
  LAYER ME3 ;
  RECT 207.745 0.000 208.065 0.717 ;
  LAYER ME2 ;
  RECT 207.745 0.000 208.065 0.717 ;
  LAYER ME2 ;
  RECT 207.745 0.000 208.065 0.717 ;
  LAYER ME1 ;
  RECT 207.745 0.000 208.065 0.717 ;
  LAYER ME1 ;
  RECT 207.745 0.000 208.065 0.717 ;
 END
 ANTENNAPARTIALMETALAREA                  5.305 LAYER ME2 ;
 ANTENNAGATEAREA                          0.612 LAYER ME2 ;
 ANTENNAGATEAREA                          0.612 LAYER ME3 ;
 ANTENNAGATEAREA                          0.612 LAYER ME4 ;
 ANTENNADIFFAREA                          0.218 LAYER ME2 ;
 ANTENNADIFFAREA                          0.218 LAYER ME3 ;
 ANTENNADIFFAREA                          0.218 LAYER ME4 ;
 ANTENNAMAXAREACAR                       53.132 LAYER ME2 ;
 ANTENNAMAXAREACAR                       55.256 LAYER ME3 ;
 ANTENNAMAXAREACAR                       57.381 LAYER ME4 ;
END DVSE
PIN DVS3
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 207.225 0.000 207.545 0.717 ;
  LAYER ME3 ;
  RECT 207.225 0.000 207.545 0.717 ;
  LAYER ME3 ;
  RECT 207.225 0.000 207.545 0.717 ;
  LAYER ME2 ;
  RECT 207.225 0.000 207.545 0.717 ;
  LAYER ME2 ;
  RECT 207.225 0.000 207.545 0.717 ;
  LAYER ME1 ;
  RECT 207.225 0.000 207.545 0.717 ;
  LAYER ME1 ;
  RECT 207.225 0.000 207.545 0.717 ;
 END
 ANTENNAPARTIALMETALAREA                  3.675 LAYER ME2 ;
 ANTENNAGATEAREA                          0.108 LAYER ME2 ;
 ANTENNAGATEAREA                          0.108 LAYER ME3 ;
 ANTENNAGATEAREA                          0.108 LAYER ME4 ;
 ANTENNADIFFAREA                          0.218 LAYER ME2 ;
 ANTENNADIFFAREA                          0.218 LAYER ME3 ;
 ANTENNADIFFAREA                          0.218 LAYER ME4 ;
 ANTENNAMAXAREACAR                       45.625 LAYER ME2 ;
 ANTENNAMAXAREACAR                       47.749 LAYER ME3 ;
 ANTENNAMAXAREACAR                       49.874 LAYER ME4 ;
END DVS3
PIN DVS2
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 208.265 0.000 208.585 0.717 ;
  LAYER ME3 ;
  RECT 208.265 0.000 208.585 0.717 ;
  LAYER ME3 ;
  RECT 208.265 0.000 208.585 0.717 ;
  LAYER ME2 ;
  RECT 208.265 0.000 208.585 0.717 ;
  LAYER ME2 ;
  RECT 208.265 0.000 208.585 0.717 ;
  LAYER ME1 ;
  RECT 208.265 0.000 208.585 0.717 ;
  LAYER ME1 ;
  RECT 208.265 0.000 208.585 0.717 ;
 END
 ANTENNAPARTIALMETALAREA                  5.371 LAYER ME2 ;
 ANTENNAGATEAREA                          0.108 LAYER ME2 ;
 ANTENNAGATEAREA                          0.108 LAYER ME3 ;
 ANTENNAGATEAREA                          0.108 LAYER ME4 ;
 ANTENNADIFFAREA                          0.218 LAYER ME2 ;
 ANTENNADIFFAREA                          0.218 LAYER ME3 ;
 ANTENNADIFFAREA                          0.218 LAYER ME4 ;
 ANTENNAMAXAREACAR                       60.060 LAYER ME2 ;
 ANTENNAMAXAREACAR                       62.184 LAYER ME3 ;
 ANTENNAMAXAREACAR                       64.309 LAYER ME4 ;
END DVS2
PIN DVS1
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 206.705 0.000 207.025 0.717 ;
  LAYER ME3 ;
  RECT 206.705 0.000 207.025 0.717 ;
  LAYER ME3 ;
  RECT 206.705 0.000 207.025 0.717 ;
  LAYER ME2 ;
  RECT 206.705 0.000 207.025 0.717 ;
  LAYER ME2 ;
  RECT 206.705 0.000 207.025 0.717 ;
  LAYER ME1 ;
  RECT 206.705 0.000 207.025 0.717 ;
  LAYER ME1 ;
  RECT 206.705 0.000 207.025 0.717 ;
 END
 ANTENNAPARTIALMETALAREA                  3.307 LAYER ME2 ;
 ANTENNAGATEAREA                          0.108 LAYER ME2 ;
 ANTENNAGATEAREA                          0.108 LAYER ME3 ;
 ANTENNAGATEAREA                          0.108 LAYER ME4 ;
 ANTENNADIFFAREA                          0.218 LAYER ME2 ;
 ANTENNADIFFAREA                          0.218 LAYER ME3 ;
 ANTENNADIFFAREA                          0.218 LAYER ME4 ;
 ANTENNAMAXAREACAR                       42.063 LAYER ME2 ;
 ANTENNAMAXAREACAR                       44.188 LAYER ME3 ;
 ANTENNAMAXAREACAR                       46.312 LAYER ME4 ;
END DVS1
PIN DVS0
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 208.785 0.000 209.105 0.693 ;
  LAYER ME3 ;
  RECT 208.785 0.000 209.105 0.693 ;
  LAYER ME3 ;
  RECT 208.785 0.000 209.105 0.693 ;
  LAYER ME2 ;
  RECT 208.785 0.000 209.105 0.693 ;
  LAYER ME2 ;
  RECT 208.785 0.000 209.105 0.693 ;
  LAYER ME1 ;
  RECT 208.785 0.000 209.105 0.693 ;
  LAYER ME1 ;
  RECT 208.785 0.000 209.105 0.693 ;
 END
 ANTENNAPARTIALMETALAREA                  4.376 LAYER ME2 ;
 ANTENNAGATEAREA                          0.108 LAYER ME2 ;
 ANTENNAGATEAREA                          0.108 LAYER ME3 ;
 ANTENNAGATEAREA                          0.108 LAYER ME4 ;
 ANTENNADIFFAREA                          0.218 LAYER ME2 ;
 ANTENNADIFFAREA                          0.218 LAYER ME3 ;
 ANTENNADIFFAREA                          0.218 LAYER ME4 ;
 ANTENNAMAXAREACAR                       53.260 LAYER ME2 ;
 ANTENNAMAXAREACAR                       55.313 LAYER ME3 ;
 ANTENNAMAXAREACAR                       57.367 LAYER ME4 ;
END DVS0
PIN CK
  DIRECTION INPUT ;
 PORT
  LAYER ME3 ;
  RECT 200.221 0.000 200.541 0.713 ;
  LAYER ME2 ;
  RECT 200.221 0.000 200.541 0.713 ;
  LAYER ME1 ;
  RECT 200.221 0.000 200.541 0.713 ;
 END
 ANTENNAPARTIALMETALAREA                  2.392 LAYER ME2 ;
 ANTENNAPARTIALMETALAREA                  7.363 LAYER ME3 ;
 ANTENNAGATEAREA                          0.072 LAYER ME2 ;
 ANTENNAGATEAREA                          1.260 LAYER ME3 ;
 ANTENNADIFFAREA                          0.218 LAYER ME2 ;
 ANTENNADIFFAREA                          0.218 LAYER ME3 ;
 ANTENNAMAXAREACAR                       46.148 LAYER ME2 ;
 ANTENNAMAXAREACAR                      151.587 LAYER ME3 ;
END CK
PIN CSB
  DIRECTION INPUT ;
 PORT
  LAYER ME3 ;
  RECT 193.433 0.000 193.753 0.712 ;
  LAYER ME2 ;
  RECT 193.433 0.000 193.753 0.712 ;
  LAYER ME1 ;
  RECT 193.433 0.000 193.753 0.712 ;
 END
 ANTENNAPARTIALMETALAREA                  3.350 LAYER ME2 ;
 ANTENNAPARTIALMETALAREA                  7.235 LAYER ME3 ;
 ANTENNAGATEAREA                          2.244 LAYER ME2 ;
 ANTENNAGATEAREA                          3.216 LAYER ME3 ;
 ANTENNADIFFAREA                          0.218 LAYER ME2 ;
 ANTENNADIFFAREA                          0.218 LAYER ME3 ;
 ANTENNAMAXAREACAR                       17.231 LAYER ME2 ;
 ANTENNAMAXAREACAR                       51.784 LAYER ME3 ;
END CSB
PIN DI41
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 374.611 0.000 374.891 0.720 ;
  LAYER ME3 ;
  RECT 374.611 0.000 374.891 0.720 ;
  LAYER ME2 ;
  RECT 374.611 0.000 374.891 0.720 ;
  LAYER ME1 ;
  RECT 374.611 0.000 374.891 0.720 ;
 END
 ANTENNAPARTIALMETALAREA                  0.805 LAYER ME1 ;
 ANTENNAGATEAREA                          0.072 LAYER ME1 ;
 ANTENNAGATEAREA                          0.072 LAYER ME2 ;
 ANTENNAGATEAREA                          0.072 LAYER ME3 ;
 ANTENNAGATEAREA                          0.072 LAYER ME4 ;
 ANTENNADIFFAREA                          0.218 LAYER ME1 ;
 ANTENNADIFFAREA                          0.218 LAYER ME2 ;
 ANTENNADIFFAREA                          0.218 LAYER ME3 ;
 ANTENNADIFFAREA                          0.218 LAYER ME4 ;
 ANTENNAMAXAREACAR                       13.984 LAYER ME1 ;
 ANTENNAMAXAREACAR                       16.784 LAYER ME2 ;
 ANTENNAMAXAREACAR                       19.584 LAYER ME3 ;
 ANTENNAMAXAREACAR                       22.384 LAYER ME4 ;
END DI41
PIN DO41
  DIRECTION OUTPUT ;
 PORT
  LAYER ME4 ;
  RECT 372.633 0.000 372.913 0.720 ;
  LAYER ME3 ;
  RECT 372.633 0.000 372.913 0.720 ;
  LAYER ME2 ;
  RECT 372.633 0.000 372.913 0.720 ;
  LAYER ME1 ;
  RECT 372.633 0.000 372.913 0.720 ;
 END
 ANTENNAPARTIALMETALAREA                  2.030 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME3 ;
 ANTENNADIFFAREA                          1.293 LAYER ME4 ;
END DO41
PIN DI40
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 366.603 0.000 366.883 0.720 ;
  LAYER ME3 ;
  RECT 366.603 0.000 366.883 0.720 ;
  LAYER ME2 ;
  RECT 366.603 0.000 366.883 0.720 ;
  LAYER ME1 ;
  RECT 366.603 0.000 366.883 0.720 ;
 END
 ANTENNAPARTIALMETALAREA                  0.805 LAYER ME1 ;
 ANTENNAGATEAREA                          0.072 LAYER ME1 ;
 ANTENNAGATEAREA                          0.072 LAYER ME2 ;
 ANTENNAGATEAREA                          0.072 LAYER ME3 ;
 ANTENNAGATEAREA                          0.072 LAYER ME4 ;
 ANTENNADIFFAREA                          0.218 LAYER ME1 ;
 ANTENNADIFFAREA                          0.218 LAYER ME2 ;
 ANTENNADIFFAREA                          0.218 LAYER ME3 ;
 ANTENNADIFFAREA                          0.218 LAYER ME4 ;
 ANTENNAMAXAREACAR                       13.984 LAYER ME1 ;
 ANTENNAMAXAREACAR                       16.784 LAYER ME2 ;
 ANTENNAMAXAREACAR                       19.584 LAYER ME3 ;
 ANTENNAMAXAREACAR                       22.384 LAYER ME4 ;
END DI40
PIN DO40
  DIRECTION OUTPUT ;
 PORT
  LAYER ME4 ;
  RECT 364.625 0.000 364.905 0.720 ;
  LAYER ME3 ;
  RECT 364.625 0.000 364.905 0.720 ;
  LAYER ME2 ;
  RECT 364.625 0.000 364.905 0.720 ;
  LAYER ME1 ;
  RECT 364.625 0.000 364.905 0.720 ;
 END
 ANTENNAPARTIALMETALAREA                  2.030 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME3 ;
 ANTENNADIFFAREA                          1.293 LAYER ME4 ;
END DO40
PIN DI39
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 358.595 0.000 358.875 0.720 ;
  LAYER ME3 ;
  RECT 358.595 0.000 358.875 0.720 ;
  LAYER ME2 ;
  RECT 358.595 0.000 358.875 0.720 ;
  LAYER ME1 ;
  RECT 358.595 0.000 358.875 0.720 ;
 END
 ANTENNAPARTIALMETALAREA                  0.805 LAYER ME1 ;
 ANTENNAGATEAREA                          0.072 LAYER ME1 ;
 ANTENNAGATEAREA                          0.072 LAYER ME2 ;
 ANTENNAGATEAREA                          0.072 LAYER ME3 ;
 ANTENNAGATEAREA                          0.072 LAYER ME4 ;
 ANTENNADIFFAREA                          0.218 LAYER ME1 ;
 ANTENNADIFFAREA                          0.218 LAYER ME2 ;
 ANTENNADIFFAREA                          0.218 LAYER ME3 ;
 ANTENNADIFFAREA                          0.218 LAYER ME4 ;
 ANTENNAMAXAREACAR                       13.984 LAYER ME1 ;
 ANTENNAMAXAREACAR                       16.784 LAYER ME2 ;
 ANTENNAMAXAREACAR                       19.584 LAYER ME3 ;
 ANTENNAMAXAREACAR                       22.384 LAYER ME4 ;
END DI39
PIN DO39
  DIRECTION OUTPUT ;
 PORT
  LAYER ME4 ;
  RECT 356.617 0.000 356.897 0.720 ;
  LAYER ME3 ;
  RECT 356.617 0.000 356.897 0.720 ;
  LAYER ME2 ;
  RECT 356.617 0.000 356.897 0.720 ;
  LAYER ME1 ;
  RECT 356.617 0.000 356.897 0.720 ;
 END
 ANTENNAPARTIALMETALAREA                  2.030 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME3 ;
 ANTENNADIFFAREA                          1.293 LAYER ME4 ;
END DO39
PIN DI38
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 350.587 0.000 350.867 0.720 ;
  LAYER ME3 ;
  RECT 350.587 0.000 350.867 0.720 ;
  LAYER ME2 ;
  RECT 350.587 0.000 350.867 0.720 ;
  LAYER ME1 ;
  RECT 350.587 0.000 350.867 0.720 ;
 END
 ANTENNAPARTIALMETALAREA                  0.805 LAYER ME1 ;
 ANTENNAGATEAREA                          0.072 LAYER ME1 ;
 ANTENNAGATEAREA                          0.072 LAYER ME2 ;
 ANTENNAGATEAREA                          0.072 LAYER ME3 ;
 ANTENNAGATEAREA                          0.072 LAYER ME4 ;
 ANTENNADIFFAREA                          0.218 LAYER ME1 ;
 ANTENNADIFFAREA                          0.218 LAYER ME2 ;
 ANTENNADIFFAREA                          0.218 LAYER ME3 ;
 ANTENNADIFFAREA                          0.218 LAYER ME4 ;
 ANTENNAMAXAREACAR                       13.984 LAYER ME1 ;
 ANTENNAMAXAREACAR                       16.784 LAYER ME2 ;
 ANTENNAMAXAREACAR                       19.584 LAYER ME3 ;
 ANTENNAMAXAREACAR                       22.384 LAYER ME4 ;
END DI38
PIN DO38
  DIRECTION OUTPUT ;
 PORT
  LAYER ME4 ;
  RECT 348.609 0.000 348.889 0.720 ;
  LAYER ME3 ;
  RECT 348.609 0.000 348.889 0.720 ;
  LAYER ME2 ;
  RECT 348.609 0.000 348.889 0.720 ;
  LAYER ME1 ;
  RECT 348.609 0.000 348.889 0.720 ;
 END
 ANTENNAPARTIALMETALAREA                  2.030 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME3 ;
 ANTENNADIFFAREA                          1.293 LAYER ME4 ;
END DO38
PIN DI37
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 342.579 0.000 342.859 0.720 ;
  LAYER ME3 ;
  RECT 342.579 0.000 342.859 0.720 ;
  LAYER ME2 ;
  RECT 342.579 0.000 342.859 0.720 ;
  LAYER ME1 ;
  RECT 342.579 0.000 342.859 0.720 ;
 END
 ANTENNAPARTIALMETALAREA                  0.805 LAYER ME1 ;
 ANTENNAGATEAREA                          0.072 LAYER ME1 ;
 ANTENNAGATEAREA                          0.072 LAYER ME2 ;
 ANTENNAGATEAREA                          0.072 LAYER ME3 ;
 ANTENNAGATEAREA                          0.072 LAYER ME4 ;
 ANTENNADIFFAREA                          0.218 LAYER ME1 ;
 ANTENNADIFFAREA                          0.218 LAYER ME2 ;
 ANTENNADIFFAREA                          0.218 LAYER ME3 ;
 ANTENNADIFFAREA                          0.218 LAYER ME4 ;
 ANTENNAMAXAREACAR                       13.984 LAYER ME1 ;
 ANTENNAMAXAREACAR                       16.784 LAYER ME2 ;
 ANTENNAMAXAREACAR                       19.584 LAYER ME3 ;
 ANTENNAMAXAREACAR                       22.384 LAYER ME4 ;
END DI37
PIN DO37
  DIRECTION OUTPUT ;
 PORT
  LAYER ME4 ;
  RECT 340.601 0.000 340.881 0.720 ;
  LAYER ME3 ;
  RECT 340.601 0.000 340.881 0.720 ;
  LAYER ME2 ;
  RECT 340.601 0.000 340.881 0.720 ;
  LAYER ME1 ;
  RECT 340.601 0.000 340.881 0.720 ;
 END
 ANTENNAPARTIALMETALAREA                  2.030 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME3 ;
 ANTENNADIFFAREA                          1.293 LAYER ME4 ;
END DO37
PIN DI36
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 334.571 0.000 334.851 0.720 ;
  LAYER ME3 ;
  RECT 334.571 0.000 334.851 0.720 ;
  LAYER ME2 ;
  RECT 334.571 0.000 334.851 0.720 ;
  LAYER ME1 ;
  RECT 334.571 0.000 334.851 0.720 ;
 END
 ANTENNAPARTIALMETALAREA                  0.805 LAYER ME1 ;
 ANTENNAGATEAREA                          0.072 LAYER ME1 ;
 ANTENNAGATEAREA                          0.072 LAYER ME2 ;
 ANTENNAGATEAREA                          0.072 LAYER ME3 ;
 ANTENNAGATEAREA                          0.072 LAYER ME4 ;
 ANTENNADIFFAREA                          0.218 LAYER ME1 ;
 ANTENNADIFFAREA                          0.218 LAYER ME2 ;
 ANTENNADIFFAREA                          0.218 LAYER ME3 ;
 ANTENNADIFFAREA                          0.218 LAYER ME4 ;
 ANTENNAMAXAREACAR                       13.984 LAYER ME1 ;
 ANTENNAMAXAREACAR                       16.784 LAYER ME2 ;
 ANTENNAMAXAREACAR                       19.584 LAYER ME3 ;
 ANTENNAMAXAREACAR                       22.384 LAYER ME4 ;
END DI36
PIN DO36
  DIRECTION OUTPUT ;
 PORT
  LAYER ME4 ;
  RECT 332.593 0.000 332.873 0.720 ;
  LAYER ME3 ;
  RECT 332.593 0.000 332.873 0.720 ;
  LAYER ME2 ;
  RECT 332.593 0.000 332.873 0.720 ;
  LAYER ME1 ;
  RECT 332.593 0.000 332.873 0.720 ;
 END
 ANTENNAPARTIALMETALAREA                  2.030 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME3 ;
 ANTENNADIFFAREA                          1.293 LAYER ME4 ;
END DO36
PIN DI35
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 326.563 0.000 326.843 0.720 ;
  LAYER ME3 ;
  RECT 326.563 0.000 326.843 0.720 ;
  LAYER ME2 ;
  RECT 326.563 0.000 326.843 0.720 ;
  LAYER ME1 ;
  RECT 326.563 0.000 326.843 0.720 ;
 END
 ANTENNAPARTIALMETALAREA                  0.522 LAYER ME1 ;
 ANTENNAGATEAREA                          0.072 LAYER ME1 ;
 ANTENNAGATEAREA                          0.072 LAYER ME2 ;
 ANTENNAGATEAREA                          0.072 LAYER ME3 ;
 ANTENNAGATEAREA                          0.072 LAYER ME4 ;
 ANTENNADIFFAREA                          0.218 LAYER ME1 ;
 ANTENNADIFFAREA                          0.218 LAYER ME2 ;
 ANTENNADIFFAREA                          0.218 LAYER ME3 ;
 ANTENNADIFFAREA                          0.218 LAYER ME4 ;
 ANTENNAMAXAREACAR                       10.048 LAYER ME1 ;
 ANTENNAMAXAREACAR                       12.848 LAYER ME2 ;
 ANTENNAMAXAREACAR                       15.648 LAYER ME3 ;
 ANTENNAMAXAREACAR                       18.448 LAYER ME4 ;
END DI35
PIN DO35
  DIRECTION OUTPUT ;
 PORT
  LAYER ME4 ;
  RECT 324.505 0.000 324.785 0.720 ;
  LAYER ME3 ;
  RECT 324.505 0.000 324.785 0.720 ;
  LAYER ME2 ;
  RECT 324.505 0.000 324.785 0.720 ;
  LAYER ME1 ;
  RECT 324.505 0.000 324.785 0.720 ;
 END
 ANTENNAPARTIALMETALAREA                  2.030 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME3 ;
 ANTENNADIFFAREA                          1.293 LAYER ME4 ;
END DO35
PIN WEB5
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 324.985 0.000 325.265 0.720 ;
  LAYER ME3 ;
  RECT 324.985 0.000 325.265 0.720 ;
  LAYER ME2 ;
  RECT 324.985 0.000 325.265 0.720 ;
  LAYER ME1 ;
  RECT 324.985 0.000 325.265 0.720 ;
 END
 ANTENNAPARTIALMETALAREA                  0.436 LAYER ME2 ;
 ANTENNAGATEAREA                          0.288 LAYER ME2 ;
 ANTENNAGATEAREA                          0.288 LAYER ME3 ;
 ANTENNAGATEAREA                          0.288 LAYER ME4 ;
 ANTENNADIFFAREA                          0.218 LAYER ME2 ;
 ANTENNADIFFAREA                          0.218 LAYER ME3 ;
 ANTENNADIFFAREA                          0.218 LAYER ME4 ;
 ANTENNAMAXAREACAR                        4.602 LAYER ME2 ;
 ANTENNAMAXAREACAR                        5.302 LAYER ME3 ;
 ANTENNAMAXAREACAR                        6.002 LAYER ME4 ;
END WEB5
PIN DI34
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 318.555 0.000 318.835 0.720 ;
  LAYER ME3 ;
  RECT 318.555 0.000 318.835 0.720 ;
  LAYER ME2 ;
  RECT 318.555 0.000 318.835 0.720 ;
  LAYER ME1 ;
  RECT 318.555 0.000 318.835 0.720 ;
 END
 ANTENNAPARTIALMETALAREA                  0.805 LAYER ME1 ;
 ANTENNAGATEAREA                          0.072 LAYER ME1 ;
 ANTENNAGATEAREA                          0.072 LAYER ME2 ;
 ANTENNAGATEAREA                          0.072 LAYER ME3 ;
 ANTENNAGATEAREA                          0.072 LAYER ME4 ;
 ANTENNADIFFAREA                          0.218 LAYER ME1 ;
 ANTENNADIFFAREA                          0.218 LAYER ME2 ;
 ANTENNADIFFAREA                          0.218 LAYER ME3 ;
 ANTENNADIFFAREA                          0.218 LAYER ME4 ;
 ANTENNAMAXAREACAR                       13.984 LAYER ME1 ;
 ANTENNAMAXAREACAR                       16.784 LAYER ME2 ;
 ANTENNAMAXAREACAR                       19.584 LAYER ME3 ;
 ANTENNAMAXAREACAR                       22.384 LAYER ME4 ;
END DI34
PIN DO34
  DIRECTION OUTPUT ;
 PORT
  LAYER ME4 ;
  RECT 316.577 0.000 316.857 0.720 ;
  LAYER ME3 ;
  RECT 316.577 0.000 316.857 0.720 ;
  LAYER ME2 ;
  RECT 316.577 0.000 316.857 0.720 ;
  LAYER ME1 ;
  RECT 316.577 0.000 316.857 0.720 ;
 END
 ANTENNAPARTIALMETALAREA                  2.030 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME3 ;
 ANTENNADIFFAREA                          1.293 LAYER ME4 ;
END DO34
PIN DI33
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 310.547 0.000 310.827 0.720 ;
  LAYER ME3 ;
  RECT 310.547 0.000 310.827 0.720 ;
  LAYER ME2 ;
  RECT 310.547 0.000 310.827 0.720 ;
  LAYER ME1 ;
  RECT 310.547 0.000 310.827 0.720 ;
 END
 ANTENNAPARTIALMETALAREA                  0.805 LAYER ME1 ;
 ANTENNAGATEAREA                          0.072 LAYER ME1 ;
 ANTENNAGATEAREA                          0.072 LAYER ME2 ;
 ANTENNAGATEAREA                          0.072 LAYER ME3 ;
 ANTENNAGATEAREA                          0.072 LAYER ME4 ;
 ANTENNADIFFAREA                          0.218 LAYER ME1 ;
 ANTENNADIFFAREA                          0.218 LAYER ME2 ;
 ANTENNADIFFAREA                          0.218 LAYER ME3 ;
 ANTENNADIFFAREA                          0.218 LAYER ME4 ;
 ANTENNAMAXAREACAR                       13.984 LAYER ME1 ;
 ANTENNAMAXAREACAR                       16.784 LAYER ME2 ;
 ANTENNAMAXAREACAR                       19.584 LAYER ME3 ;
 ANTENNAMAXAREACAR                       22.384 LAYER ME4 ;
END DI33
PIN DO33
  DIRECTION OUTPUT ;
 PORT
  LAYER ME4 ;
  RECT 308.569 0.000 308.849 0.720 ;
  LAYER ME3 ;
  RECT 308.569 0.000 308.849 0.720 ;
  LAYER ME2 ;
  RECT 308.569 0.000 308.849 0.720 ;
  LAYER ME1 ;
  RECT 308.569 0.000 308.849 0.720 ;
 END
 ANTENNAPARTIALMETALAREA                  2.030 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME3 ;
 ANTENNADIFFAREA                          1.293 LAYER ME4 ;
END DO33
PIN DI32
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 302.539 0.000 302.819 0.720 ;
  LAYER ME3 ;
  RECT 302.539 0.000 302.819 0.720 ;
  LAYER ME2 ;
  RECT 302.539 0.000 302.819 0.720 ;
  LAYER ME1 ;
  RECT 302.539 0.000 302.819 0.720 ;
 END
 ANTENNAPARTIALMETALAREA                  0.805 LAYER ME1 ;
 ANTENNAGATEAREA                          0.072 LAYER ME1 ;
 ANTENNAGATEAREA                          0.072 LAYER ME2 ;
 ANTENNAGATEAREA                          0.072 LAYER ME3 ;
 ANTENNAGATEAREA                          0.072 LAYER ME4 ;
 ANTENNADIFFAREA                          0.218 LAYER ME1 ;
 ANTENNADIFFAREA                          0.218 LAYER ME2 ;
 ANTENNADIFFAREA                          0.218 LAYER ME3 ;
 ANTENNADIFFAREA                          0.218 LAYER ME4 ;
 ANTENNAMAXAREACAR                       13.984 LAYER ME1 ;
 ANTENNAMAXAREACAR                       16.784 LAYER ME2 ;
 ANTENNAMAXAREACAR                       19.584 LAYER ME3 ;
 ANTENNAMAXAREACAR                       22.384 LAYER ME4 ;
END DI32
PIN DO32
  DIRECTION OUTPUT ;
 PORT
  LAYER ME4 ;
  RECT 300.561 0.000 300.841 0.720 ;
  LAYER ME3 ;
  RECT 300.561 0.000 300.841 0.720 ;
  LAYER ME2 ;
  RECT 300.561 0.000 300.841 0.720 ;
  LAYER ME1 ;
  RECT 300.561 0.000 300.841 0.720 ;
 END
 ANTENNAPARTIALMETALAREA                  2.030 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME3 ;
 ANTENNADIFFAREA                          1.293 LAYER ME4 ;
END DO32
PIN DI31
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 294.531 0.000 294.811 0.720 ;
  LAYER ME3 ;
  RECT 294.531 0.000 294.811 0.720 ;
  LAYER ME2 ;
  RECT 294.531 0.000 294.811 0.720 ;
  LAYER ME1 ;
  RECT 294.531 0.000 294.811 0.720 ;
 END
 ANTENNAPARTIALMETALAREA                  0.805 LAYER ME1 ;
 ANTENNAGATEAREA                          0.072 LAYER ME1 ;
 ANTENNAGATEAREA                          0.072 LAYER ME2 ;
 ANTENNAGATEAREA                          0.072 LAYER ME3 ;
 ANTENNAGATEAREA                          0.072 LAYER ME4 ;
 ANTENNADIFFAREA                          0.218 LAYER ME1 ;
 ANTENNADIFFAREA                          0.218 LAYER ME2 ;
 ANTENNADIFFAREA                          0.218 LAYER ME3 ;
 ANTENNADIFFAREA                          0.218 LAYER ME4 ;
 ANTENNAMAXAREACAR                       13.984 LAYER ME1 ;
 ANTENNAMAXAREACAR                       16.784 LAYER ME2 ;
 ANTENNAMAXAREACAR                       19.584 LAYER ME3 ;
 ANTENNAMAXAREACAR                       22.384 LAYER ME4 ;
END DI31
PIN DO31
  DIRECTION OUTPUT ;
 PORT
  LAYER ME4 ;
  RECT 292.553 0.000 292.833 0.720 ;
  LAYER ME3 ;
  RECT 292.553 0.000 292.833 0.720 ;
  LAYER ME2 ;
  RECT 292.553 0.000 292.833 0.720 ;
  LAYER ME1 ;
  RECT 292.553 0.000 292.833 0.720 ;
 END
 ANTENNAPARTIALMETALAREA                  2.030 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME3 ;
 ANTENNADIFFAREA                          1.293 LAYER ME4 ;
END DO31
PIN DI30
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 286.523 0.000 286.803 0.720 ;
  LAYER ME3 ;
  RECT 286.523 0.000 286.803 0.720 ;
  LAYER ME2 ;
  RECT 286.523 0.000 286.803 0.720 ;
  LAYER ME1 ;
  RECT 286.523 0.000 286.803 0.720 ;
 END
 ANTENNAPARTIALMETALAREA                  0.805 LAYER ME1 ;
 ANTENNAGATEAREA                          0.072 LAYER ME1 ;
 ANTENNAGATEAREA                          0.072 LAYER ME2 ;
 ANTENNAGATEAREA                          0.072 LAYER ME3 ;
 ANTENNAGATEAREA                          0.072 LAYER ME4 ;
 ANTENNADIFFAREA                          0.218 LAYER ME1 ;
 ANTENNADIFFAREA                          0.218 LAYER ME2 ;
 ANTENNADIFFAREA                          0.218 LAYER ME3 ;
 ANTENNADIFFAREA                          0.218 LAYER ME4 ;
 ANTENNAMAXAREACAR                       13.984 LAYER ME1 ;
 ANTENNAMAXAREACAR                       16.784 LAYER ME2 ;
 ANTENNAMAXAREACAR                       19.584 LAYER ME3 ;
 ANTENNAMAXAREACAR                       22.384 LAYER ME4 ;
END DI30
PIN DO30
  DIRECTION OUTPUT ;
 PORT
  LAYER ME4 ;
  RECT 284.545 0.000 284.825 0.720 ;
  LAYER ME3 ;
  RECT 284.545 0.000 284.825 0.720 ;
  LAYER ME2 ;
  RECT 284.545 0.000 284.825 0.720 ;
  LAYER ME1 ;
  RECT 284.545 0.000 284.825 0.720 ;
 END
 ANTENNAPARTIALMETALAREA                  2.030 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME3 ;
 ANTENNADIFFAREA                          1.293 LAYER ME4 ;
END DO30
PIN DI29
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 278.515 0.000 278.795 0.720 ;
  LAYER ME3 ;
  RECT 278.515 0.000 278.795 0.720 ;
  LAYER ME2 ;
  RECT 278.515 0.000 278.795 0.720 ;
  LAYER ME1 ;
  RECT 278.515 0.000 278.795 0.720 ;
 END
 ANTENNAPARTIALMETALAREA                  0.805 LAYER ME1 ;
 ANTENNAGATEAREA                          0.072 LAYER ME1 ;
 ANTENNAGATEAREA                          0.072 LAYER ME2 ;
 ANTENNAGATEAREA                          0.072 LAYER ME3 ;
 ANTENNAGATEAREA                          0.072 LAYER ME4 ;
 ANTENNADIFFAREA                          0.218 LAYER ME1 ;
 ANTENNADIFFAREA                          0.218 LAYER ME2 ;
 ANTENNADIFFAREA                          0.218 LAYER ME3 ;
 ANTENNADIFFAREA                          0.218 LAYER ME4 ;
 ANTENNAMAXAREACAR                       13.984 LAYER ME1 ;
 ANTENNAMAXAREACAR                       16.784 LAYER ME2 ;
 ANTENNAMAXAREACAR                       19.584 LAYER ME3 ;
 ANTENNAMAXAREACAR                       22.384 LAYER ME4 ;
END DI29
PIN DO29
  DIRECTION OUTPUT ;
 PORT
  LAYER ME4 ;
  RECT 276.537 0.000 276.817 0.720 ;
  LAYER ME3 ;
  RECT 276.537 0.000 276.817 0.720 ;
  LAYER ME2 ;
  RECT 276.537 0.000 276.817 0.720 ;
  LAYER ME1 ;
  RECT 276.537 0.000 276.817 0.720 ;
 END
 ANTENNAPARTIALMETALAREA                  2.030 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME3 ;
 ANTENNADIFFAREA                          1.293 LAYER ME4 ;
END DO29
PIN DI28
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 270.507 0.000 270.787 0.720 ;
  LAYER ME3 ;
  RECT 270.507 0.000 270.787 0.720 ;
  LAYER ME2 ;
  RECT 270.507 0.000 270.787 0.720 ;
  LAYER ME1 ;
  RECT 270.507 0.000 270.787 0.720 ;
 END
 ANTENNAPARTIALMETALAREA                  0.522 LAYER ME1 ;
 ANTENNAGATEAREA                          0.072 LAYER ME1 ;
 ANTENNAGATEAREA                          0.072 LAYER ME2 ;
 ANTENNAGATEAREA                          0.072 LAYER ME3 ;
 ANTENNAGATEAREA                          0.072 LAYER ME4 ;
 ANTENNADIFFAREA                          0.218 LAYER ME1 ;
 ANTENNADIFFAREA                          0.218 LAYER ME2 ;
 ANTENNADIFFAREA                          0.218 LAYER ME3 ;
 ANTENNADIFFAREA                          0.218 LAYER ME4 ;
 ANTENNAMAXAREACAR                       10.048 LAYER ME1 ;
 ANTENNAMAXAREACAR                       12.848 LAYER ME2 ;
 ANTENNAMAXAREACAR                       15.648 LAYER ME3 ;
 ANTENNAMAXAREACAR                       18.448 LAYER ME4 ;
END DI28
PIN DO28
  DIRECTION OUTPUT ;
 PORT
  LAYER ME4 ;
  RECT 268.449 0.000 268.729 0.720 ;
  LAYER ME3 ;
  RECT 268.449 0.000 268.729 0.720 ;
  LAYER ME2 ;
  RECT 268.449 0.000 268.729 0.720 ;
  LAYER ME1 ;
  RECT 268.449 0.000 268.729 0.720 ;
 END
 ANTENNAPARTIALMETALAREA                  2.030 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME3 ;
 ANTENNADIFFAREA                          1.293 LAYER ME4 ;
END DO28
PIN WEB4
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 268.929 0.000 269.209 0.720 ;
  LAYER ME3 ;
  RECT 268.929 0.000 269.209 0.720 ;
  LAYER ME2 ;
  RECT 268.929 0.000 269.209 0.720 ;
  LAYER ME1 ;
  RECT 268.929 0.000 269.209 0.720 ;
 END
 ANTENNAPARTIALMETALAREA                  0.436 LAYER ME2 ;
 ANTENNAGATEAREA                          0.288 LAYER ME2 ;
 ANTENNAGATEAREA                          0.288 LAYER ME3 ;
 ANTENNAGATEAREA                          0.288 LAYER ME4 ;
 ANTENNADIFFAREA                          0.218 LAYER ME2 ;
 ANTENNADIFFAREA                          0.218 LAYER ME3 ;
 ANTENNADIFFAREA                          0.218 LAYER ME4 ;
 ANTENNAMAXAREACAR                        4.602 LAYER ME2 ;
 ANTENNAMAXAREACAR                        5.302 LAYER ME3 ;
 ANTENNAMAXAREACAR                        6.002 LAYER ME4 ;
END WEB4
PIN DI27
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 262.499 0.000 262.779 0.720 ;
  LAYER ME3 ;
  RECT 262.499 0.000 262.779 0.720 ;
  LAYER ME2 ;
  RECT 262.499 0.000 262.779 0.720 ;
  LAYER ME1 ;
  RECT 262.499 0.000 262.779 0.720 ;
 END
 ANTENNAPARTIALMETALAREA                  0.805 LAYER ME1 ;
 ANTENNAGATEAREA                          0.072 LAYER ME1 ;
 ANTENNAGATEAREA                          0.072 LAYER ME2 ;
 ANTENNAGATEAREA                          0.072 LAYER ME3 ;
 ANTENNAGATEAREA                          0.072 LAYER ME4 ;
 ANTENNADIFFAREA                          0.218 LAYER ME1 ;
 ANTENNADIFFAREA                          0.218 LAYER ME2 ;
 ANTENNADIFFAREA                          0.218 LAYER ME3 ;
 ANTENNADIFFAREA                          0.218 LAYER ME4 ;
 ANTENNAMAXAREACAR                       13.984 LAYER ME1 ;
 ANTENNAMAXAREACAR                       16.784 LAYER ME2 ;
 ANTENNAMAXAREACAR                       19.584 LAYER ME3 ;
 ANTENNAMAXAREACAR                       22.384 LAYER ME4 ;
END DI27
PIN DO27
  DIRECTION OUTPUT ;
 PORT
  LAYER ME4 ;
  RECT 260.521 0.000 260.801 0.720 ;
  LAYER ME3 ;
  RECT 260.521 0.000 260.801 0.720 ;
  LAYER ME2 ;
  RECT 260.521 0.000 260.801 0.720 ;
  LAYER ME1 ;
  RECT 260.521 0.000 260.801 0.720 ;
 END
 ANTENNAPARTIALMETALAREA                  2.030 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME3 ;
 ANTENNADIFFAREA                          1.293 LAYER ME4 ;
END DO27
PIN DI26
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 254.491 0.000 254.771 0.720 ;
  LAYER ME3 ;
  RECT 254.491 0.000 254.771 0.720 ;
  LAYER ME2 ;
  RECT 254.491 0.000 254.771 0.720 ;
  LAYER ME1 ;
  RECT 254.491 0.000 254.771 0.720 ;
 END
 ANTENNAPARTIALMETALAREA                  0.805 LAYER ME1 ;
 ANTENNAGATEAREA                          0.072 LAYER ME1 ;
 ANTENNAGATEAREA                          0.072 LAYER ME2 ;
 ANTENNAGATEAREA                          0.072 LAYER ME3 ;
 ANTENNAGATEAREA                          0.072 LAYER ME4 ;
 ANTENNADIFFAREA                          0.218 LAYER ME1 ;
 ANTENNADIFFAREA                          0.218 LAYER ME2 ;
 ANTENNADIFFAREA                          0.218 LAYER ME3 ;
 ANTENNADIFFAREA                          0.218 LAYER ME4 ;
 ANTENNAMAXAREACAR                       13.984 LAYER ME1 ;
 ANTENNAMAXAREACAR                       16.784 LAYER ME2 ;
 ANTENNAMAXAREACAR                       19.584 LAYER ME3 ;
 ANTENNAMAXAREACAR                       22.384 LAYER ME4 ;
END DI26
PIN DO26
  DIRECTION OUTPUT ;
 PORT
  LAYER ME4 ;
  RECT 252.513 0.000 252.793 0.720 ;
  LAYER ME3 ;
  RECT 252.513 0.000 252.793 0.720 ;
  LAYER ME2 ;
  RECT 252.513 0.000 252.793 0.720 ;
  LAYER ME1 ;
  RECT 252.513 0.000 252.793 0.720 ;
 END
 ANTENNAPARTIALMETALAREA                  2.030 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME3 ;
 ANTENNADIFFAREA                          1.293 LAYER ME4 ;
END DO26
PIN DI25
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 246.483 0.000 246.763 0.720 ;
  LAYER ME3 ;
  RECT 246.483 0.000 246.763 0.720 ;
  LAYER ME2 ;
  RECT 246.483 0.000 246.763 0.720 ;
  LAYER ME1 ;
  RECT 246.483 0.000 246.763 0.720 ;
 END
 ANTENNAPARTIALMETALAREA                  0.805 LAYER ME1 ;
 ANTENNAGATEAREA                          0.072 LAYER ME1 ;
 ANTENNAGATEAREA                          0.072 LAYER ME2 ;
 ANTENNAGATEAREA                          0.072 LAYER ME3 ;
 ANTENNAGATEAREA                          0.072 LAYER ME4 ;
 ANTENNADIFFAREA                          0.218 LAYER ME1 ;
 ANTENNADIFFAREA                          0.218 LAYER ME2 ;
 ANTENNADIFFAREA                          0.218 LAYER ME3 ;
 ANTENNADIFFAREA                          0.218 LAYER ME4 ;
 ANTENNAMAXAREACAR                       13.984 LAYER ME1 ;
 ANTENNAMAXAREACAR                       16.784 LAYER ME2 ;
 ANTENNAMAXAREACAR                       19.584 LAYER ME3 ;
 ANTENNAMAXAREACAR                       22.384 LAYER ME4 ;
END DI25
PIN DO25
  DIRECTION OUTPUT ;
 PORT
  LAYER ME4 ;
  RECT 244.505 0.000 244.785 0.720 ;
  LAYER ME3 ;
  RECT 244.505 0.000 244.785 0.720 ;
  LAYER ME2 ;
  RECT 244.505 0.000 244.785 0.720 ;
  LAYER ME1 ;
  RECT 244.505 0.000 244.785 0.720 ;
 END
 ANTENNAPARTIALMETALAREA                  2.030 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME3 ;
 ANTENNADIFFAREA                          1.293 LAYER ME4 ;
END DO25
PIN DI24
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 238.475 0.000 238.755 0.720 ;
  LAYER ME3 ;
  RECT 238.475 0.000 238.755 0.720 ;
  LAYER ME2 ;
  RECT 238.475 0.000 238.755 0.720 ;
  LAYER ME1 ;
  RECT 238.475 0.000 238.755 0.720 ;
 END
 ANTENNAPARTIALMETALAREA                  0.805 LAYER ME1 ;
 ANTENNAGATEAREA                          0.072 LAYER ME1 ;
 ANTENNAGATEAREA                          0.072 LAYER ME2 ;
 ANTENNAGATEAREA                          0.072 LAYER ME3 ;
 ANTENNAGATEAREA                          0.072 LAYER ME4 ;
 ANTENNADIFFAREA                          0.218 LAYER ME1 ;
 ANTENNADIFFAREA                          0.218 LAYER ME2 ;
 ANTENNADIFFAREA                          0.218 LAYER ME3 ;
 ANTENNADIFFAREA                          0.218 LAYER ME4 ;
 ANTENNAMAXAREACAR                       13.984 LAYER ME1 ;
 ANTENNAMAXAREACAR                       16.784 LAYER ME2 ;
 ANTENNAMAXAREACAR                       19.584 LAYER ME3 ;
 ANTENNAMAXAREACAR                       22.384 LAYER ME4 ;
END DI24
PIN DO24
  DIRECTION OUTPUT ;
 PORT
  LAYER ME4 ;
  RECT 236.497 0.000 236.777 0.720 ;
  LAYER ME3 ;
  RECT 236.497 0.000 236.777 0.720 ;
  LAYER ME2 ;
  RECT 236.497 0.000 236.777 0.720 ;
  LAYER ME1 ;
  RECT 236.497 0.000 236.777 0.720 ;
 END
 ANTENNAPARTIALMETALAREA                  2.030 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME3 ;
 ANTENNADIFFAREA                          1.293 LAYER ME4 ;
END DO24
PIN DI23
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 230.467 0.000 230.747 0.720 ;
  LAYER ME3 ;
  RECT 230.467 0.000 230.747 0.720 ;
  LAYER ME2 ;
  RECT 230.467 0.000 230.747 0.720 ;
  LAYER ME1 ;
  RECT 230.467 0.000 230.747 0.720 ;
 END
 ANTENNAPARTIALMETALAREA                  0.805 LAYER ME1 ;
 ANTENNAGATEAREA                          0.072 LAYER ME1 ;
 ANTENNAGATEAREA                          0.072 LAYER ME2 ;
 ANTENNAGATEAREA                          0.072 LAYER ME3 ;
 ANTENNAGATEAREA                          0.072 LAYER ME4 ;
 ANTENNADIFFAREA                          0.218 LAYER ME1 ;
 ANTENNADIFFAREA                          0.218 LAYER ME2 ;
 ANTENNADIFFAREA                          0.218 LAYER ME3 ;
 ANTENNADIFFAREA                          0.218 LAYER ME4 ;
 ANTENNAMAXAREACAR                       13.984 LAYER ME1 ;
 ANTENNAMAXAREACAR                       16.784 LAYER ME2 ;
 ANTENNAMAXAREACAR                       19.584 LAYER ME3 ;
 ANTENNAMAXAREACAR                       22.384 LAYER ME4 ;
END DI23
PIN DO23
  DIRECTION OUTPUT ;
 PORT
  LAYER ME4 ;
  RECT 228.489 0.000 228.769 0.720 ;
  LAYER ME3 ;
  RECT 228.489 0.000 228.769 0.720 ;
  LAYER ME2 ;
  RECT 228.489 0.000 228.769 0.720 ;
  LAYER ME1 ;
  RECT 228.489 0.000 228.769 0.720 ;
 END
 ANTENNAPARTIALMETALAREA                  2.030 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME3 ;
 ANTENNADIFFAREA                          1.293 LAYER ME4 ;
END DO23
PIN DI22
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 222.459 0.000 222.739 0.720 ;
  LAYER ME3 ;
  RECT 222.459 0.000 222.739 0.720 ;
  LAYER ME2 ;
  RECT 222.459 0.000 222.739 0.720 ;
  LAYER ME1 ;
  RECT 222.459 0.000 222.739 0.720 ;
 END
 ANTENNAPARTIALMETALAREA                  0.805 LAYER ME1 ;
 ANTENNAGATEAREA                          0.072 LAYER ME1 ;
 ANTENNAGATEAREA                          0.072 LAYER ME2 ;
 ANTENNAGATEAREA                          0.072 LAYER ME3 ;
 ANTENNAGATEAREA                          0.072 LAYER ME4 ;
 ANTENNADIFFAREA                          0.218 LAYER ME1 ;
 ANTENNADIFFAREA                          0.218 LAYER ME2 ;
 ANTENNADIFFAREA                          0.218 LAYER ME3 ;
 ANTENNADIFFAREA                          0.218 LAYER ME4 ;
 ANTENNAMAXAREACAR                       13.984 LAYER ME1 ;
 ANTENNAMAXAREACAR                       16.784 LAYER ME2 ;
 ANTENNAMAXAREACAR                       19.584 LAYER ME3 ;
 ANTENNAMAXAREACAR                       22.384 LAYER ME4 ;
END DI22
PIN DO22
  DIRECTION OUTPUT ;
 PORT
  LAYER ME4 ;
  RECT 220.481 0.000 220.761 0.720 ;
  LAYER ME3 ;
  RECT 220.481 0.000 220.761 0.720 ;
  LAYER ME2 ;
  RECT 220.481 0.000 220.761 0.720 ;
  LAYER ME1 ;
  RECT 220.481 0.000 220.761 0.720 ;
 END
 ANTENNAPARTIALMETALAREA                  2.030 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME3 ;
 ANTENNADIFFAREA                          1.293 LAYER ME4 ;
END DO22
PIN DI21
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 214.451 0.000 214.731 0.720 ;
  LAYER ME3 ;
  RECT 214.451 0.000 214.731 0.720 ;
  LAYER ME2 ;
  RECT 214.451 0.000 214.731 0.720 ;
  LAYER ME1 ;
  RECT 214.451 0.000 214.731 0.720 ;
 END
 ANTENNAPARTIALMETALAREA                  0.522 LAYER ME1 ;
 ANTENNAGATEAREA                          0.072 LAYER ME1 ;
 ANTENNAGATEAREA                          0.072 LAYER ME2 ;
 ANTENNAGATEAREA                          0.072 LAYER ME3 ;
 ANTENNAGATEAREA                          0.072 LAYER ME4 ;
 ANTENNADIFFAREA                          0.218 LAYER ME1 ;
 ANTENNADIFFAREA                          0.218 LAYER ME2 ;
 ANTENNADIFFAREA                          0.218 LAYER ME3 ;
 ANTENNADIFFAREA                          0.218 LAYER ME4 ;
 ANTENNAMAXAREACAR                       10.048 LAYER ME1 ;
 ANTENNAMAXAREACAR                       12.848 LAYER ME2 ;
 ANTENNAMAXAREACAR                       15.648 LAYER ME3 ;
 ANTENNAMAXAREACAR                       18.448 LAYER ME4 ;
END DI21
PIN DO21
  DIRECTION OUTPUT ;
 PORT
  LAYER ME4 ;
  RECT 212.393 0.000 212.673 0.720 ;
  LAYER ME3 ;
  RECT 212.393 0.000 212.673 0.720 ;
  LAYER ME2 ;
  RECT 212.393 0.000 212.673 0.720 ;
  LAYER ME1 ;
  RECT 212.393 0.000 212.673 0.720 ;
 END
 ANTENNAPARTIALMETALAREA                  2.030 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME3 ;
 ANTENNADIFFAREA                          1.293 LAYER ME4 ;
END DO21
PIN WEB3
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 212.873 0.000 213.153 0.720 ;
  LAYER ME3 ;
  RECT 212.873 0.000 213.153 0.720 ;
  LAYER ME2 ;
  RECT 212.873 0.000 213.153 0.720 ;
  LAYER ME1 ;
  RECT 212.873 0.000 213.153 0.720 ;
 END
 ANTENNAPARTIALMETALAREA                  0.436 LAYER ME2 ;
 ANTENNAGATEAREA                          0.288 LAYER ME2 ;
 ANTENNAGATEAREA                          0.288 LAYER ME3 ;
 ANTENNAGATEAREA                          0.288 LAYER ME4 ;
 ANTENNADIFFAREA                          0.218 LAYER ME2 ;
 ANTENNADIFFAREA                          0.218 LAYER ME3 ;
 ANTENNADIFFAREA                          0.218 LAYER ME4 ;
 ANTENNAMAXAREACAR                        4.602 LAYER ME2 ;
 ANTENNAMAXAREACAR                        5.302 LAYER ME3 ;
 ANTENNAMAXAREACAR                        6.002 LAYER ME4 ;
END WEB3
OBS
  LAYER ME3 ;
  RECT 0.000 0.000 379.835 68.179 ;
  LAYER ME2 ;
  RECT 0.000 0.000 379.835 68.179 ;
  LAYER ME1 ;
  RECT 0.000 0.000 379.835 68.179 ;
  LAYER ME4 ;
  RECT 0.000 0.000 183.910 68.179 ;
  LAYER ME4 ;
  RECT 185.564 0.000 186.684 68.179 ;
  LAYER ME4 ;
  RECT 188.279 0.000 188.999 68.179 ;
  LAYER ME4 ;
  RECT 189.729 0.000 190.449 68.179 ;
  LAYER ME4 ;
  RECT 192.509 0.000 193.109 68.179 ;
  LAYER ME4 ;
  RECT 195.723 0.000 197.409 68.179 ;
  LAYER ME4 ;
  RECT 198.799 0.000 199.919 68.179 ;
  LAYER ME4 ;
  RECT 201.194 0.000 201.914 68.179 ;
  LAYER ME4 ;
  RECT 202.909 0.000 203.629 68.179 ;
  LAYER ME4 ;
  RECT 204.829 0.000 379.835 68.179 ;
END
END SYKB110_128X7X6CM4
END LIBRARY





