# ________________________________________________________________________________________________
# 
# 
#             Synchronous Two-Port Register File Compiler
# 
#                 UMC 0.11um LL AE Logic Process
# 
# ________________________________________________________________________________________________
# 
#               
#         Copyright (C) 2024 Faraday Technology Corporation. All Rights Reserved.       
#                
#         This source code is an unpublished work belongs to Faraday Technology Corporation       
#         It is considered a trade secret and is not to be divulged or       
#         used by parties who have not received written authorization from       
#         Faraday Technology Corporation       
#                
#         Faraday's home page can be found at: http://www.faraday-tech.com/       
#                
# ________________________________________________________________________________________________
# 
#        IP Name            :  FSR0K_D_SZ                
#        IP Version         :  1.7.0                     
#        IP Release Status  :  Active                    
#        Word               :  256                       
#        Bit                :  9                         
#        Byte               :  8                         
#        Mux                :  2                         
#        Output Loading     :  0.01                      
#        Clock Input Slew   :  0.016                     
#        Data Input Slew    :  0.016                     
#        Ring Type          :  Ringless Model            
#        Ring Width         :  0                         
#        Bus Format         :  0                         
#        Memaker Path       :  /home/mem/Desktop/memlib  
#        GUI Version        :  m20230904                 
#        Date               :  2024/09/10 14:55:51       
# ________________________________________________________________________________________________
# 

VERSION 5.5 ;
NAMESCASESENSITIVE ON ;
MACRO SZKD110_256X9X8CM2
CLASS BLOCK ;
FOREIGN SZKD110_256X9X8CM2 0.000 0.000 ;
ORIGIN 0.000 0.000 ;
SIZE 539.250 BY 221.080 ;
SYMMETRY x y r90 ;
SITE core ;
PIN VCC
  DIRECTION INOUT ;
  USE POWER ;
 PORT
  LAYER ME4 ;
  RECT 300.870 0.000 301.290 221.080 ;
 END
 PORT
  LAYER ME4 ;
  RECT 301.770 197.090 302.370 221.080 ;
 END
 PORT
  LAYER ME4 ;
  RECT 304.170 0.000 304.590 220.280 ;
 END
 PORT
  LAYER ME4 ;
  RECT 307.470 0.000 307.890 221.080 ;
 END
 PORT
  LAYER ME4 ;
  RECT 308.370 197.090 308.970 221.080 ;
 END
 PORT
  LAYER ME4 ;
  RECT 310.770 0.000 311.190 220.280 ;
 END
 PORT
  LAYER ME4 ;
  RECT 314.070 0.000 314.490 221.080 ;
 END
 PORT
  LAYER ME4 ;
  RECT 314.970 197.090 315.570 221.080 ;
 END
 PORT
  LAYER ME4 ;
  RECT 317.370 0.000 317.790 220.280 ;
 END
 PORT
  LAYER ME4 ;
  RECT 320.670 0.000 321.090 221.080 ;
 END
 PORT
  LAYER ME4 ;
  RECT 321.570 197.090 322.170 221.080 ;
 END
 PORT
  LAYER ME4 ;
  RECT 323.970 0.000 324.390 220.280 ;
 END
 PORT
  LAYER ME4 ;
  RECT 327.270 0.000 327.690 221.080 ;
 END
 PORT
  LAYER ME4 ;
  RECT 328.170 197.090 328.770 221.080 ;
 END
 PORT
  LAYER ME4 ;
  RECT 330.570 0.000 330.990 220.280 ;
 END
 PORT
  LAYER ME4 ;
  RECT 333.870 0.000 334.290 221.080 ;
 END
 PORT
  LAYER ME4 ;
  RECT 334.770 197.090 335.370 221.080 ;
 END
 PORT
  LAYER ME4 ;
  RECT 337.170 0.000 337.590 220.280 ;
 END
 PORT
  LAYER ME4 ;
  RECT 340.470 0.000 340.890 221.080 ;
 END
 PORT
  LAYER ME4 ;
  RECT 341.370 197.090 341.970 221.080 ;
 END
 PORT
  LAYER ME4 ;
  RECT 343.770 0.000 344.190 220.280 ;
 END
 PORT
  LAYER ME4 ;
  RECT 347.070 0.000 347.490 221.080 ;
 END
 PORT
  LAYER ME4 ;
  RECT 347.970 197.090 348.570 221.080 ;
 END
 PORT
  LAYER ME4 ;
  RECT 350.370 0.000 350.790 220.280 ;
 END
 PORT
  LAYER ME4 ;
  RECT 353.670 0.000 354.090 221.080 ;
 END
 PORT
  LAYER ME4 ;
  RECT 354.570 197.090 355.170 221.080 ;
 END
 PORT
  LAYER ME4 ;
  RECT 356.970 0.000 357.390 220.280 ;
 END
 PORT
  LAYER ME4 ;
  RECT 360.270 0.000 360.690 221.080 ;
 END
 PORT
  LAYER ME4 ;
  RECT 361.170 197.090 361.770 221.080 ;
 END
 PORT
  LAYER ME4 ;
  RECT 363.570 0.000 363.990 220.280 ;
 END
 PORT
  LAYER ME4 ;
  RECT 366.870 0.000 367.290 221.080 ;
 END
 PORT
  LAYER ME4 ;
  RECT 367.770 197.090 368.370 221.080 ;
 END
 PORT
  LAYER ME4 ;
  RECT 370.170 0.000 370.590 220.280 ;
 END
 PORT
  LAYER ME4 ;
  RECT 373.470 0.000 373.890 221.080 ;
 END
 PORT
  LAYER ME4 ;
  RECT 374.370 197.090 374.970 221.080 ;
 END
 PORT
  LAYER ME4 ;
  RECT 376.770 0.000 377.190 220.280 ;
 END
 PORT
  LAYER ME4 ;
  RECT 380.070 0.000 380.490 221.080 ;
 END
 PORT
  LAYER ME4 ;
  RECT 380.970 197.090 381.570 221.080 ;
 END
 PORT
  LAYER ME4 ;
  RECT 383.370 0.000 383.790 220.280 ;
 END
 PORT
  LAYER ME4 ;
  RECT 386.670 0.000 387.090 221.080 ;
 END
 PORT
  LAYER ME4 ;
  RECT 387.570 197.090 388.170 221.080 ;
 END
 PORT
  LAYER ME4 ;
  RECT 389.970 0.000 390.390 220.280 ;
 END
 PORT
  LAYER ME4 ;
  RECT 393.270 0.000 393.690 221.080 ;
 END
 PORT
  LAYER ME4 ;
  RECT 394.170 197.090 394.770 221.080 ;
 END
 PORT
  LAYER ME4 ;
  RECT 396.570 0.000 396.990 220.280 ;
 END
 PORT
  LAYER ME4 ;
  RECT 399.870 0.000 400.290 221.080 ;
 END
 PORT
  LAYER ME4 ;
  RECT 400.770 197.090 401.370 221.080 ;
 END
 PORT
  LAYER ME4 ;
  RECT 403.170 0.000 403.590 220.280 ;
 END
 PORT
  LAYER ME4 ;
  RECT 406.470 0.000 406.890 221.080 ;
 END
 PORT
  LAYER ME4 ;
  RECT 407.370 197.090 407.970 221.080 ;
 END
 PORT
  LAYER ME4 ;
  RECT 409.770 0.000 410.190 220.280 ;
 END
 PORT
  LAYER ME4 ;
  RECT 413.070 0.000 413.490 221.080 ;
 END
 PORT
  LAYER ME4 ;
  RECT 413.970 197.090 414.570 221.080 ;
 END
 PORT
  LAYER ME4 ;
  RECT 416.370 0.000 416.790 220.280 ;
 END
 PORT
  LAYER ME4 ;
  RECT 419.670 0.000 420.090 221.080 ;
 END
 PORT
  LAYER ME4 ;
  RECT 420.570 197.090 421.170 221.080 ;
 END
 PORT
  LAYER ME4 ;
  RECT 422.970 0.000 423.390 220.280 ;
 END
 PORT
  LAYER ME4 ;
  RECT 426.270 0.000 426.690 221.080 ;
 END
 PORT
  LAYER ME4 ;
  RECT 427.170 197.090 427.770 221.080 ;
 END
 PORT
  LAYER ME4 ;
  RECT 429.570 0.000 429.990 220.280 ;
 END
 PORT
  LAYER ME4 ;
  RECT 432.870 0.000 433.290 221.080 ;
 END
 PORT
  LAYER ME4 ;
  RECT 433.770 197.090 434.370 221.080 ;
 END
 PORT
  LAYER ME4 ;
  RECT 436.170 0.000 436.590 220.280 ;
 END
 PORT
  LAYER ME4 ;
  RECT 439.470 0.000 439.890 221.080 ;
 END
 PORT
  LAYER ME4 ;
  RECT 440.370 197.090 440.970 221.080 ;
 END
 PORT
  LAYER ME4 ;
  RECT 442.770 0.000 443.190 220.280 ;
 END
 PORT
  LAYER ME4 ;
  RECT 446.070 0.000 446.490 221.080 ;
 END
 PORT
  LAYER ME4 ;
  RECT 446.970 197.090 447.570 221.080 ;
 END
 PORT
  LAYER ME4 ;
  RECT 449.370 0.000 449.790 220.280 ;
 END
 PORT
  LAYER ME4 ;
  RECT 452.670 0.000 453.090 221.080 ;
 END
 PORT
  LAYER ME4 ;
  RECT 453.570 197.090 454.170 221.080 ;
 END
 PORT
  LAYER ME4 ;
  RECT 455.970 0.000 456.390 220.280 ;
 END
 PORT
  LAYER ME4 ;
  RECT 459.270 0.000 459.690 221.080 ;
 END
 PORT
  LAYER ME4 ;
  RECT 460.170 197.090 460.770 221.080 ;
 END
 PORT
  LAYER ME4 ;
  RECT 462.570 0.000 462.990 220.280 ;
 END
 PORT
  LAYER ME4 ;
  RECT 465.870 0.000 466.290 221.080 ;
 END
 PORT
  LAYER ME4 ;
  RECT 466.770 197.090 467.370 221.080 ;
 END
 PORT
  LAYER ME4 ;
  RECT 469.170 0.000 469.590 220.280 ;
 END
 PORT
  LAYER ME4 ;
  RECT 472.470 0.000 472.890 221.080 ;
 END
 PORT
  LAYER ME4 ;
  RECT 473.370 197.090 473.970 221.080 ;
 END
 PORT
  LAYER ME4 ;
  RECT 475.770 0.000 476.190 220.280 ;
 END
 PORT
  LAYER ME4 ;
  RECT 479.070 0.000 479.490 221.080 ;
 END
 PORT
  LAYER ME4 ;
  RECT 479.970 197.090 480.570 221.080 ;
 END
 PORT
  LAYER ME4 ;
  RECT 482.370 0.000 482.790 220.280 ;
 END
 PORT
  LAYER ME4 ;
  RECT 485.670 0.000 486.090 221.080 ;
 END
 PORT
  LAYER ME4 ;
  RECT 486.570 197.090 487.170 221.080 ;
 END
 PORT
  LAYER ME4 ;
  RECT 488.970 0.000 489.390 220.280 ;
 END
 PORT
  LAYER ME4 ;
  RECT 492.270 0.000 492.690 221.080 ;
 END
 PORT
  LAYER ME4 ;
  RECT 493.170 197.090 493.770 221.080 ;
 END
 PORT
  LAYER ME4 ;
  RECT 495.570 0.000 495.990 220.280 ;
 END
 PORT
  LAYER ME4 ;
  RECT 498.870 0.000 499.290 221.080 ;
 END
 PORT
  LAYER ME4 ;
  RECT 499.770 197.090 500.370 221.080 ;
 END
 PORT
  LAYER ME4 ;
  RECT 502.170 0.000 502.590 220.280 ;
 END
 PORT
  LAYER ME4 ;
  RECT 505.470 0.000 505.890 221.080 ;
 END
 PORT
  LAYER ME4 ;
  RECT 506.370 197.090 506.970 221.080 ;
 END
 PORT
  LAYER ME4 ;
  RECT 508.770 0.000 509.190 220.280 ;
 END
 PORT
  LAYER ME4 ;
  RECT 512.070 0.000 512.490 221.080 ;
 END
 PORT
  LAYER ME4 ;
  RECT 512.970 197.090 513.570 221.080 ;
 END
 PORT
  LAYER ME4 ;
  RECT 515.370 0.000 515.790 220.280 ;
 END
 PORT
  LAYER ME4 ;
  RECT 518.670 0.000 519.090 221.080 ;
 END
 PORT
  LAYER ME4 ;
  RECT 519.570 197.090 520.170 221.080 ;
 END
 PORT
  LAYER ME4 ;
  RECT 521.970 0.000 522.390 220.280 ;
 END
 PORT
  LAYER ME4 ;
  RECT 525.270 0.000 525.690 221.080 ;
 END
 PORT
  LAYER ME4 ;
  RECT 526.170 197.090 526.770 221.080 ;
 END
 PORT
  LAYER ME4 ;
  RECT 528.570 0.000 528.990 220.280 ;
 END
 PORT
  LAYER ME4 ;
  RECT 531.870 0.000 532.290 221.080 ;
 END
 PORT
  LAYER ME4 ;
  RECT 532.770 197.090 533.370 221.080 ;
 END
 PORT
  LAYER ME4 ;
  RECT 535.170 0.000 535.590 220.280 ;
 END
 PORT
  LAYER ME4 ;
  RECT 538.480 192.316 538.880 221.080 ;
 END
 PORT
  LAYER ME4 ;
  RECT 297.570 0.000 297.990 221.080 ;
 END
 PORT
  LAYER ME4 ;
  RECT 294.270 0.800 294.690 220.250 ;
 END
 PORT
  LAYER ME4 ;
  RECT 290.980 0.000 291.380 221.080 ;
 END
 PORT
  LAYER ME4 ;
  RECT 538.480 24.565 538.880 192.315 ;
 END
 PORT
  LAYER ME4 ;
  RECT 538.480 0.000 538.880 24.564 ;
 END
 PORT
  LAYER ME4 ;
  RECT 303.090 0.000 303.690 20.650 ;
 END
 PORT
  LAYER ME4 ;
  RECT 309.690 0.000 310.290 20.650 ;
 END
 PORT
  LAYER ME4 ;
  RECT 316.290 0.000 316.890 20.650 ;
 END
 PORT
  LAYER ME4 ;
  RECT 322.890 0.000 323.490 20.650 ;
 END
 PORT
  LAYER ME4 ;
  RECT 329.490 0.000 330.090 20.650 ;
 END
 PORT
  LAYER ME4 ;
  RECT 336.090 0.000 336.690 20.650 ;
 END
 PORT
  LAYER ME4 ;
  RECT 342.690 0.000 343.290 20.650 ;
 END
 PORT
  LAYER ME4 ;
  RECT 349.290 0.000 349.890 20.650 ;
 END
 PORT
  LAYER ME4 ;
  RECT 355.890 0.000 356.490 20.650 ;
 END
 PORT
  LAYER ME4 ;
  RECT 362.490 0.000 363.090 20.650 ;
 END
 PORT
  LAYER ME4 ;
  RECT 369.090 0.000 369.690 20.650 ;
 END
 PORT
  LAYER ME4 ;
  RECT 375.690 0.000 376.290 20.650 ;
 END
 PORT
  LAYER ME4 ;
  RECT 382.290 0.000 382.890 20.650 ;
 END
 PORT
  LAYER ME4 ;
  RECT 388.890 0.000 389.490 20.650 ;
 END
 PORT
  LAYER ME4 ;
  RECT 395.490 0.000 396.090 20.650 ;
 END
 PORT
  LAYER ME4 ;
  RECT 402.090 0.000 402.690 20.650 ;
 END
 PORT
  LAYER ME4 ;
  RECT 408.690 0.000 409.290 20.650 ;
 END
 PORT
  LAYER ME4 ;
  RECT 415.290 0.000 415.890 20.650 ;
 END
 PORT
  LAYER ME4 ;
  RECT 421.890 0.000 422.490 20.650 ;
 END
 PORT
  LAYER ME4 ;
  RECT 428.490 0.000 429.090 20.650 ;
 END
 PORT
  LAYER ME4 ;
  RECT 435.090 0.000 435.690 20.650 ;
 END
 PORT
  LAYER ME4 ;
  RECT 441.690 0.000 442.290 20.650 ;
 END
 PORT
  LAYER ME4 ;
  RECT 448.290 0.000 448.890 20.650 ;
 END
 PORT
  LAYER ME4 ;
  RECT 454.890 0.000 455.490 20.650 ;
 END
 PORT
  LAYER ME4 ;
  RECT 461.490 0.000 462.090 20.650 ;
 END
 PORT
  LAYER ME4 ;
  RECT 468.090 0.000 468.690 20.650 ;
 END
 PORT
  LAYER ME4 ;
  RECT 474.690 0.000 475.290 20.650 ;
 END
 PORT
  LAYER ME4 ;
  RECT 481.290 0.000 481.890 20.650 ;
 END
 PORT
  LAYER ME4 ;
  RECT 487.890 0.000 488.490 20.650 ;
 END
 PORT
  LAYER ME4 ;
  RECT 494.490 0.000 495.090 20.650 ;
 END
 PORT
  LAYER ME4 ;
  RECT 501.090 0.000 501.690 20.650 ;
 END
 PORT
  LAYER ME4 ;
  RECT 507.690 0.000 508.290 20.650 ;
 END
 PORT
  LAYER ME4 ;
  RECT 514.290 0.000 514.890 20.650 ;
 END
 PORT
  LAYER ME4 ;
  RECT 520.890 0.000 521.490 20.650 ;
 END
 PORT
  LAYER ME4 ;
  RECT 527.490 0.000 528.090 20.650 ;
 END
 PORT
  LAYER ME4 ;
  RECT 534.090 0.000 534.690 20.650 ;
 END
 PORT
  LAYER ME4 ;
  RECT 0.370 0.000 0.770 221.080 ;
 END
 PORT
  LAYER ME4 ;
  RECT 3.660 0.000 4.080 221.080 ;
 END
 PORT
  LAYER ME4 ;
  RECT 4.560 197.090 5.160 221.080 ;
 END
 PORT
  LAYER ME4 ;
  RECT 6.960 0.000 7.380 220.280 ;
 END
 PORT
  LAYER ME4 ;
  RECT 10.260 0.000 10.680 221.080 ;
 END
 PORT
  LAYER ME4 ;
  RECT 11.160 197.090 11.760 221.080 ;
 END
 PORT
  LAYER ME4 ;
  RECT 13.560 0.000 13.980 220.280 ;
 END
 PORT
  LAYER ME4 ;
  RECT 16.860 0.000 17.280 221.080 ;
 END
 PORT
  LAYER ME4 ;
  RECT 17.760 197.090 18.360 221.080 ;
 END
 PORT
  LAYER ME4 ;
  RECT 20.160 0.000 20.580 220.280 ;
 END
 PORT
  LAYER ME4 ;
  RECT 23.460 0.000 23.880 221.080 ;
 END
 PORT
  LAYER ME4 ;
  RECT 24.360 197.090 24.960 221.080 ;
 END
 PORT
  LAYER ME4 ;
  RECT 26.760 0.000 27.180 220.280 ;
 END
 PORT
  LAYER ME4 ;
  RECT 30.060 0.000 30.480 221.080 ;
 END
 PORT
  LAYER ME4 ;
  RECT 30.960 197.090 31.560 221.080 ;
 END
 PORT
  LAYER ME4 ;
  RECT 33.360 0.000 33.780 220.280 ;
 END
 PORT
  LAYER ME4 ;
  RECT 36.660 0.000 37.080 221.080 ;
 END
 PORT
  LAYER ME4 ;
  RECT 37.560 197.090 38.160 221.080 ;
 END
 PORT
  LAYER ME4 ;
  RECT 39.960 0.000 40.380 220.280 ;
 END
 PORT
  LAYER ME4 ;
  RECT 43.260 0.000 43.680 221.080 ;
 END
 PORT
  LAYER ME4 ;
  RECT 44.160 197.090 44.760 221.080 ;
 END
 PORT
  LAYER ME4 ;
  RECT 46.560 0.000 46.980 220.280 ;
 END
 PORT
  LAYER ME4 ;
  RECT 49.860 0.000 50.280 221.080 ;
 END
 PORT
  LAYER ME4 ;
  RECT 50.760 197.090 51.360 221.080 ;
 END
 PORT
  LAYER ME4 ;
  RECT 53.160 0.000 53.580 220.280 ;
 END
 PORT
  LAYER ME4 ;
  RECT 56.460 0.000 56.880 221.080 ;
 END
 PORT
  LAYER ME4 ;
  RECT 57.360 197.090 57.960 221.080 ;
 END
 PORT
  LAYER ME4 ;
  RECT 59.760 0.000 60.180 220.280 ;
 END
 PORT
  LAYER ME4 ;
  RECT 63.060 0.000 63.480 221.080 ;
 END
 PORT
  LAYER ME4 ;
  RECT 63.960 197.090 64.560 221.080 ;
 END
 PORT
  LAYER ME4 ;
  RECT 66.360 0.000 66.780 220.280 ;
 END
 PORT
  LAYER ME4 ;
  RECT 69.660 0.000 70.080 221.080 ;
 END
 PORT
  LAYER ME4 ;
  RECT 70.560 197.090 71.160 221.080 ;
 END
 PORT
  LAYER ME4 ;
  RECT 72.960 0.000 73.380 220.280 ;
 END
 PORT
  LAYER ME4 ;
  RECT 76.260 0.000 76.680 221.080 ;
 END
 PORT
  LAYER ME4 ;
  RECT 77.160 197.090 77.760 221.080 ;
 END
 PORT
  LAYER ME4 ;
  RECT 79.560 0.000 79.980 220.280 ;
 END
 PORT
  LAYER ME4 ;
  RECT 82.860 0.000 83.280 221.080 ;
 END
 PORT
  LAYER ME4 ;
  RECT 83.760 197.090 84.360 221.080 ;
 END
 PORT
  LAYER ME4 ;
  RECT 86.160 0.000 86.580 220.280 ;
 END
 PORT
  LAYER ME4 ;
  RECT 89.460 0.000 89.880 221.080 ;
 END
 PORT
  LAYER ME4 ;
  RECT 90.360 197.090 90.960 221.080 ;
 END
 PORT
  LAYER ME4 ;
  RECT 92.760 0.000 93.180 220.280 ;
 END
 PORT
  LAYER ME4 ;
  RECT 96.060 0.000 96.480 221.080 ;
 END
 PORT
  LAYER ME4 ;
  RECT 96.960 197.090 97.560 221.080 ;
 END
 PORT
  LAYER ME4 ;
  RECT 99.360 0.000 99.780 220.280 ;
 END
 PORT
  LAYER ME4 ;
  RECT 102.660 0.000 103.080 221.080 ;
 END
 PORT
  LAYER ME4 ;
  RECT 103.560 197.090 104.160 221.080 ;
 END
 PORT
  LAYER ME4 ;
  RECT 105.960 0.000 106.380 220.280 ;
 END
 PORT
  LAYER ME4 ;
  RECT 109.260 0.000 109.680 221.080 ;
 END
 PORT
  LAYER ME4 ;
  RECT 110.160 197.090 110.760 221.080 ;
 END
 PORT
  LAYER ME4 ;
  RECT 112.560 0.000 112.980 220.280 ;
 END
 PORT
  LAYER ME4 ;
  RECT 115.860 0.000 116.280 221.080 ;
 END
 PORT
  LAYER ME4 ;
  RECT 116.760 197.090 117.360 221.080 ;
 END
 PORT
  LAYER ME4 ;
  RECT 119.160 0.000 119.580 220.280 ;
 END
 PORT
  LAYER ME4 ;
  RECT 122.460 0.000 122.880 221.080 ;
 END
 PORT
  LAYER ME4 ;
  RECT 123.360 197.090 123.960 221.080 ;
 END
 PORT
  LAYER ME4 ;
  RECT 125.760 0.000 126.180 220.280 ;
 END
 PORT
  LAYER ME4 ;
  RECT 129.060 0.000 129.480 221.080 ;
 END
 PORT
  LAYER ME4 ;
  RECT 129.960 197.090 130.560 221.080 ;
 END
 PORT
  LAYER ME4 ;
  RECT 132.360 0.000 132.780 220.280 ;
 END
 PORT
  LAYER ME4 ;
  RECT 135.660 0.000 136.080 221.080 ;
 END
 PORT
  LAYER ME4 ;
  RECT 136.560 197.090 137.160 221.080 ;
 END
 PORT
  LAYER ME4 ;
  RECT 138.960 0.000 139.380 220.280 ;
 END
 PORT
  LAYER ME4 ;
  RECT 142.260 0.000 142.680 221.080 ;
 END
 PORT
  LAYER ME4 ;
  RECT 143.160 197.090 143.760 221.080 ;
 END
 PORT
  LAYER ME4 ;
  RECT 145.560 0.000 145.980 220.280 ;
 END
 PORT
  LAYER ME4 ;
  RECT 148.860 0.000 149.280 221.080 ;
 END
 PORT
  LAYER ME4 ;
  RECT 149.760 197.090 150.360 221.080 ;
 END
 PORT
  LAYER ME4 ;
  RECT 152.160 0.000 152.580 220.280 ;
 END
 PORT
  LAYER ME4 ;
  RECT 155.460 0.000 155.880 221.080 ;
 END
 PORT
  LAYER ME4 ;
  RECT 156.360 197.090 156.960 221.080 ;
 END
 PORT
  LAYER ME4 ;
  RECT 158.760 0.000 159.180 220.280 ;
 END
 PORT
  LAYER ME4 ;
  RECT 162.060 0.000 162.480 221.080 ;
 END
 PORT
  LAYER ME4 ;
  RECT 162.960 197.090 163.560 221.080 ;
 END
 PORT
  LAYER ME4 ;
  RECT 165.360 0.000 165.780 220.280 ;
 END
 PORT
  LAYER ME4 ;
  RECT 168.660 0.000 169.080 221.080 ;
 END
 PORT
  LAYER ME4 ;
  RECT 169.560 197.090 170.160 221.080 ;
 END
 PORT
  LAYER ME4 ;
  RECT 171.960 0.000 172.380 220.280 ;
 END
 PORT
  LAYER ME4 ;
  RECT 175.260 0.000 175.680 221.080 ;
 END
 PORT
  LAYER ME4 ;
  RECT 176.160 197.090 176.760 221.080 ;
 END
 PORT
  LAYER ME4 ;
  RECT 178.560 0.000 178.980 220.280 ;
 END
 PORT
  LAYER ME4 ;
  RECT 181.860 0.000 182.280 221.080 ;
 END
 PORT
  LAYER ME4 ;
  RECT 182.760 197.090 183.360 221.080 ;
 END
 PORT
  LAYER ME4 ;
  RECT 185.160 0.000 185.580 220.280 ;
 END
 PORT
  LAYER ME4 ;
  RECT 188.460 0.000 188.880 221.080 ;
 END
 PORT
  LAYER ME4 ;
  RECT 189.360 197.090 189.960 221.080 ;
 END
 PORT
  LAYER ME4 ;
  RECT 191.760 0.000 192.180 220.280 ;
 END
 PORT
  LAYER ME4 ;
  RECT 195.060 0.000 195.480 221.080 ;
 END
 PORT
  LAYER ME4 ;
  RECT 195.960 197.090 196.560 221.080 ;
 END
 PORT
  LAYER ME4 ;
  RECT 198.360 0.000 198.780 220.280 ;
 END
 PORT
  LAYER ME4 ;
  RECT 201.660 0.000 202.080 221.080 ;
 END
 PORT
  LAYER ME4 ;
  RECT 202.560 197.090 203.160 221.080 ;
 END
 PORT
  LAYER ME4 ;
  RECT 204.960 0.000 205.380 220.280 ;
 END
 PORT
  LAYER ME4 ;
  RECT 208.260 0.000 208.680 221.080 ;
 END
 PORT
  LAYER ME4 ;
  RECT 209.160 197.090 209.760 221.080 ;
 END
 PORT
  LAYER ME4 ;
  RECT 211.560 0.000 211.980 220.280 ;
 END
 PORT
  LAYER ME4 ;
  RECT 214.860 0.000 215.280 221.080 ;
 END
 PORT
  LAYER ME4 ;
  RECT 215.760 197.090 216.360 221.080 ;
 END
 PORT
  LAYER ME4 ;
  RECT 218.160 0.000 218.580 220.280 ;
 END
 PORT
  LAYER ME4 ;
  RECT 221.460 0.000 221.880 221.080 ;
 END
 PORT
  LAYER ME4 ;
  RECT 222.360 197.090 222.960 221.080 ;
 END
 PORT
  LAYER ME4 ;
  RECT 224.760 0.000 225.180 220.280 ;
 END
 PORT
  LAYER ME4 ;
  RECT 228.060 0.000 228.480 221.080 ;
 END
 PORT
  LAYER ME4 ;
  RECT 228.960 197.090 229.560 221.080 ;
 END
 PORT
  LAYER ME4 ;
  RECT 231.360 0.000 231.780 220.280 ;
 END
 PORT
  LAYER ME4 ;
  RECT 234.660 0.000 235.080 221.080 ;
 END
 PORT
  LAYER ME4 ;
  RECT 235.560 197.090 236.160 221.080 ;
 END
 PORT
  LAYER ME4 ;
  RECT 237.960 0.000 238.380 220.280 ;
 END
 PORT
  LAYER ME4 ;
  RECT 241.270 0.000 241.670 221.080 ;
 END
 PORT
  LAYER ME4 ;
  RECT 5.880 0.000 6.480 20.650 ;
 END
 PORT
  LAYER ME4 ;
  RECT 12.480 0.000 13.080 20.650 ;
 END
 PORT
  LAYER ME4 ;
  RECT 19.080 0.000 19.680 20.650 ;
 END
 PORT
  LAYER ME4 ;
  RECT 25.680 0.000 26.280 20.650 ;
 END
 PORT
  LAYER ME4 ;
  RECT 32.280 0.000 32.880 20.650 ;
 END
 PORT
  LAYER ME4 ;
  RECT 38.880 0.000 39.480 20.650 ;
 END
 PORT
  LAYER ME4 ;
  RECT 45.480 0.000 46.080 20.650 ;
 END
 PORT
  LAYER ME4 ;
  RECT 52.080 0.000 52.680 20.650 ;
 END
 PORT
  LAYER ME4 ;
  RECT 58.680 0.000 59.280 20.650 ;
 END
 PORT
  LAYER ME4 ;
  RECT 65.280 0.000 65.880 20.650 ;
 END
 PORT
  LAYER ME4 ;
  RECT 71.880 0.000 72.480 20.650 ;
 END
 PORT
  LAYER ME4 ;
  RECT 78.480 0.000 79.080 20.650 ;
 END
 PORT
  LAYER ME4 ;
  RECT 85.080 0.000 85.680 20.650 ;
 END
 PORT
  LAYER ME4 ;
  RECT 91.680 0.000 92.280 20.650 ;
 END
 PORT
  LAYER ME4 ;
  RECT 98.280 0.000 98.880 20.650 ;
 END
 PORT
  LAYER ME4 ;
  RECT 104.880 0.000 105.480 20.650 ;
 END
 PORT
  LAYER ME4 ;
  RECT 111.480 0.000 112.080 20.650 ;
 END
 PORT
  LAYER ME4 ;
  RECT 118.080 0.000 118.680 20.650 ;
 END
 PORT
  LAYER ME4 ;
  RECT 124.680 0.000 125.280 20.650 ;
 END
 PORT
  LAYER ME4 ;
  RECT 131.280 0.000 131.880 20.650 ;
 END
 PORT
  LAYER ME4 ;
  RECT 137.880 0.000 138.480 20.650 ;
 END
 PORT
  LAYER ME4 ;
  RECT 144.480 0.000 145.080 20.650 ;
 END
 PORT
  LAYER ME4 ;
  RECT 151.080 0.000 151.680 20.650 ;
 END
 PORT
  LAYER ME4 ;
  RECT 157.680 0.000 158.280 20.650 ;
 END
 PORT
  LAYER ME4 ;
  RECT 164.280 0.000 164.880 20.650 ;
 END
 PORT
  LAYER ME4 ;
  RECT 170.880 0.000 171.480 20.650 ;
 END
 PORT
  LAYER ME4 ;
  RECT 177.480 0.000 178.080 20.650 ;
 END
 PORT
  LAYER ME4 ;
  RECT 184.080 0.000 184.680 20.650 ;
 END
 PORT
  LAYER ME4 ;
  RECT 190.680 0.000 191.280 20.650 ;
 END
 PORT
  LAYER ME4 ;
  RECT 197.280 0.000 197.880 20.650 ;
 END
 PORT
  LAYER ME4 ;
  RECT 203.880 0.000 204.480 20.650 ;
 END
 PORT
  LAYER ME4 ;
  RECT 210.480 0.000 211.080 20.650 ;
 END
 PORT
  LAYER ME4 ;
  RECT 217.080 0.000 217.680 20.650 ;
 END
 PORT
  LAYER ME4 ;
  RECT 223.680 0.000 224.280 20.650 ;
 END
 PORT
  LAYER ME4 ;
  RECT 230.280 0.000 230.880 20.650 ;
 END
 PORT
  LAYER ME4 ;
  RECT 236.880 0.000 237.480 20.650 ;
 END
 PORT
  LAYER ME4 ;
  RECT 268.320 0.000 268.920 221.080 ;
 END
 PORT
  LAYER ME4 ;
  RECT 270.520 0.800 271.120 220.250 ;
 END
 PORT
  LAYER ME4 ;
  RECT 272.720 0.800 273.320 220.250 ;
 END
 PORT
  LAYER ME4 ;
  RECT 274.920 0.000 275.520 221.080 ;
 END
 PORT
  LAYER ME4 ;
  RECT 277.120 0.000 277.720 221.080 ;
 END
 PORT
  LAYER ME4 ;
  RECT 279.320 0.000 279.920 221.080 ;
 END
 PORT
  LAYER ME4 ;
  RECT 281.970 0.800 282.570 221.080 ;
 END
 PORT
  LAYER ME4 ;
  RECT 284.170 0.000 284.770 221.080 ;
 END
 PORT
  LAYER ME4 ;
  RECT 286.370 0.000 286.970 221.080 ;
 END
 PORT
  LAYER ME4 ;
  RECT 287.470 0.000 288.070 221.080 ;
 END
 PORT
  LAYER ME4 ;
  RECT 295.170 197.090 295.770 221.080 ;
 END
 PORT
  LAYER ME4 ;
  RECT 261.470 0.000 262.070 221.080 ;
 END
 PORT
  LAYER ME4 ;
  RECT 263.670 0.000 264.270 221.080 ;
 END
 PORT
  LAYER ME4 ;
  RECT 265.870 197.090 266.470 221.080 ;
 END
 PORT
  LAYER ME4 ;
  RECT 254.870 197.090 255.470 221.080 ;
 END
 PORT
  LAYER ME4 ;
  RECT 257.070 197.090 257.670 220.250 ;
 END
 PORT
  LAYER ME4 ;
  RECT 259.270 197.090 259.870 221.080 ;
 END
 PORT
  LAYER ME4 ;
  RECT 248.510 197.090 249.110 221.080 ;
 END
 PORT
  LAYER ME4 ;
  RECT 250.710 197.090 251.310 220.250 ;
 END
 PORT
  LAYER ME4 ;
  RECT 252.910 197.090 253.510 221.080 ;
 END
 PORT
  LAYER ME4 ;
  RECT 242.150 197.090 242.750 221.080 ;
 END
 PORT
  LAYER ME4 ;
  RECT 244.350 197.090 244.950 220.250 ;
 END
 PORT
  LAYER ME4 ;
  RECT 246.550 197.090 247.150 221.080 ;
 END
 PORT
  LAYER ME4 ;
  RECT 296.490 0.000 297.090 20.650 ;
 END
 PORT
  LAYER ME4 ;
  RECT 265.870 0.000 266.470 20.650 ;
 END
 PORT
  LAYER ME4 ;
  RECT 254.870 0.000 255.470 20.650 ;
 END
 PORT
  LAYER ME4 ;
  RECT 257.070 0.800 257.670 20.650 ;
 END
 PORT
  LAYER ME4 ;
  RECT 259.270 0.000 259.870 20.650 ;
 END
 PORT
  LAYER ME4 ;
  RECT 248.510 0.000 249.110 20.650 ;
 END
 PORT
  LAYER ME4 ;
  RECT 250.710 0.800 251.310 20.650 ;
 END
 PORT
  LAYER ME4 ;
  RECT 252.910 0.000 253.510 20.650 ;
 END
 PORT
  LAYER ME4 ;
  RECT 242.150 0.000 242.750 20.650 ;
 END
 PORT
  LAYER ME4 ;
  RECT 244.350 0.800 244.950 20.650 ;
 END
 PORT
  LAYER ME4 ;
  RECT 246.550 0.000 247.150 20.650 ;
 END
END VCC
PIN GND
  DIRECTION INOUT ;
  USE GROUND ;
 PORT
  LAYER ME4 ;
  RECT 300.070 0.940 300.390 221.080 ;
 END
 PORT
  LAYER ME4 ;
  RECT 299.270 0.000 299.590 221.080 ;
 END
 PORT
  LAYER ME4 ;
  RECT 302.570 0.000 302.890 221.080 ;
 END
 PORT
  LAYER ME4 ;
  RECT 305.070 0.940 305.390 221.080 ;
 END
 PORT
  LAYER ME4 ;
  RECT 305.870 0.000 306.190 221.080 ;
 END
 PORT
  LAYER ME4 ;
  RECT 303.370 21.610 303.690 221.080 ;
 END
 PORT
  LAYER ME4 ;
  RECT 306.670 0.000 306.990 221.080 ;
 END
 PORT
  LAYER ME4 ;
  RECT 309.170 0.000 309.490 221.080 ;
 END
 PORT
  LAYER ME4 ;
  RECT 311.670 0.810 311.990 221.080 ;
 END
 PORT
  LAYER ME4 ;
  RECT 312.470 0.000 312.790 221.080 ;
 END
 PORT
  LAYER ME4 ;
  RECT 309.970 21.610 310.290 221.080 ;
 END
 PORT
  LAYER ME4 ;
  RECT 313.270 0.000 313.590 221.080 ;
 END
 PORT
  LAYER ME4 ;
  RECT 315.770 0.000 316.090 221.080 ;
 END
 PORT
  LAYER ME4 ;
  RECT 318.270 0.810 318.590 221.080 ;
 END
 PORT
  LAYER ME4 ;
  RECT 319.070 0.000 319.390 221.080 ;
 END
 PORT
  LAYER ME4 ;
  RECT 316.570 21.610 316.890 221.080 ;
 END
 PORT
  LAYER ME4 ;
  RECT 319.870 0.000 320.190 221.080 ;
 END
 PORT
  LAYER ME4 ;
  RECT 322.370 0.000 322.690 221.080 ;
 END
 PORT
  LAYER ME4 ;
  RECT 324.870 0.810 325.190 221.080 ;
 END
 PORT
  LAYER ME4 ;
  RECT 325.670 0.000 325.990 221.080 ;
 END
 PORT
  LAYER ME4 ;
  RECT 323.170 21.610 323.490 221.080 ;
 END
 PORT
  LAYER ME4 ;
  RECT 326.470 0.000 326.790 221.080 ;
 END
 PORT
  LAYER ME4 ;
  RECT 328.970 0.000 329.290 221.080 ;
 END
 PORT
  LAYER ME4 ;
  RECT 331.470 0.810 331.790 221.080 ;
 END
 PORT
  LAYER ME4 ;
  RECT 332.270 0.000 332.590 221.080 ;
 END
 PORT
  LAYER ME4 ;
  RECT 329.770 21.610 330.090 221.080 ;
 END
 PORT
  LAYER ME4 ;
  RECT 333.070 0.000 333.390 221.080 ;
 END
 PORT
  LAYER ME4 ;
  RECT 335.570 0.000 335.890 221.080 ;
 END
 PORT
  LAYER ME4 ;
  RECT 338.070 0.810 338.390 221.080 ;
 END
 PORT
  LAYER ME4 ;
  RECT 338.870 0.000 339.190 221.080 ;
 END
 PORT
  LAYER ME4 ;
  RECT 336.370 21.610 336.690 221.080 ;
 END
 PORT
  LAYER ME4 ;
  RECT 339.670 0.000 339.990 221.080 ;
 END
 PORT
  LAYER ME4 ;
  RECT 342.170 0.000 342.490 221.080 ;
 END
 PORT
  LAYER ME4 ;
  RECT 344.670 0.810 344.990 221.080 ;
 END
 PORT
  LAYER ME4 ;
  RECT 345.470 0.000 345.790 221.080 ;
 END
 PORT
  LAYER ME4 ;
  RECT 342.970 21.610 343.290 221.080 ;
 END
 PORT
  LAYER ME4 ;
  RECT 346.270 0.000 346.590 221.080 ;
 END
 PORT
  LAYER ME4 ;
  RECT 348.770 0.000 349.090 221.080 ;
 END
 PORT
  LAYER ME4 ;
  RECT 351.270 0.810 351.590 221.080 ;
 END
 PORT
  LAYER ME4 ;
  RECT 352.070 0.000 352.390 221.080 ;
 END
 PORT
  LAYER ME4 ;
  RECT 349.570 21.610 349.890 221.080 ;
 END
 PORT
  LAYER ME4 ;
  RECT 352.870 0.000 353.190 221.080 ;
 END
 PORT
  LAYER ME4 ;
  RECT 355.370 0.000 355.690 221.080 ;
 END
 PORT
  LAYER ME4 ;
  RECT 357.870 0.810 358.190 221.080 ;
 END
 PORT
  LAYER ME4 ;
  RECT 358.670 0.000 358.990 221.080 ;
 END
 PORT
  LAYER ME4 ;
  RECT 356.170 21.610 356.490 221.080 ;
 END
 PORT
  LAYER ME4 ;
  RECT 359.470 0.940 359.790 221.080 ;
 END
 PORT
  LAYER ME4 ;
  RECT 361.970 0.000 362.290 221.080 ;
 END
 PORT
  LAYER ME4 ;
  RECT 364.470 0.940 364.790 221.080 ;
 END
 PORT
  LAYER ME4 ;
  RECT 365.270 0.000 365.590 221.080 ;
 END
 PORT
  LAYER ME4 ;
  RECT 362.770 21.610 363.090 221.080 ;
 END
 PORT
  LAYER ME4 ;
  RECT 366.070 0.000 366.390 221.080 ;
 END
 PORT
  LAYER ME4 ;
  RECT 368.570 0.000 368.890 221.080 ;
 END
 PORT
  LAYER ME4 ;
  RECT 371.070 0.810 371.390 221.080 ;
 END
 PORT
  LAYER ME4 ;
  RECT 371.870 0.000 372.190 221.080 ;
 END
 PORT
  LAYER ME4 ;
  RECT 369.370 21.610 369.690 221.080 ;
 END
 PORT
  LAYER ME4 ;
  RECT 372.670 0.000 372.990 221.080 ;
 END
 PORT
  LAYER ME4 ;
  RECT 375.170 0.000 375.490 221.080 ;
 END
 PORT
  LAYER ME4 ;
  RECT 377.670 0.810 377.990 221.080 ;
 END
 PORT
  LAYER ME4 ;
  RECT 378.470 0.000 378.790 221.080 ;
 END
 PORT
  LAYER ME4 ;
  RECT 375.970 21.610 376.290 221.080 ;
 END
 PORT
  LAYER ME4 ;
  RECT 379.270 0.000 379.590 221.080 ;
 END
 PORT
  LAYER ME4 ;
  RECT 381.770 0.000 382.090 221.080 ;
 END
 PORT
  LAYER ME4 ;
  RECT 384.270 0.810 384.590 221.080 ;
 END
 PORT
  LAYER ME4 ;
  RECT 385.070 0.000 385.390 221.080 ;
 END
 PORT
  LAYER ME4 ;
  RECT 382.570 21.610 382.890 221.080 ;
 END
 PORT
  LAYER ME4 ;
  RECT 385.870 0.000 386.190 221.080 ;
 END
 PORT
  LAYER ME4 ;
  RECT 388.370 0.000 388.690 221.080 ;
 END
 PORT
  LAYER ME4 ;
  RECT 390.870 0.810 391.190 221.080 ;
 END
 PORT
  LAYER ME4 ;
  RECT 391.670 0.000 391.990 221.080 ;
 END
 PORT
  LAYER ME4 ;
  RECT 389.170 21.610 389.490 221.080 ;
 END
 PORT
  LAYER ME4 ;
  RECT 392.470 0.000 392.790 221.080 ;
 END
 PORT
  LAYER ME4 ;
  RECT 394.970 0.000 395.290 221.080 ;
 END
 PORT
  LAYER ME4 ;
  RECT 397.470 0.810 397.790 221.080 ;
 END
 PORT
  LAYER ME4 ;
  RECT 398.270 0.000 398.590 221.080 ;
 END
 PORT
  LAYER ME4 ;
  RECT 395.770 21.610 396.090 221.080 ;
 END
 PORT
  LAYER ME4 ;
  RECT 399.070 0.000 399.390 221.080 ;
 END
 PORT
  LAYER ME4 ;
  RECT 401.570 0.000 401.890 221.080 ;
 END
 PORT
  LAYER ME4 ;
  RECT 404.070 0.810 404.390 221.080 ;
 END
 PORT
  LAYER ME4 ;
  RECT 404.870 0.000 405.190 221.080 ;
 END
 PORT
  LAYER ME4 ;
  RECT 402.370 21.610 402.690 221.080 ;
 END
 PORT
  LAYER ME4 ;
  RECT 405.670 0.000 405.990 221.080 ;
 END
 PORT
  LAYER ME4 ;
  RECT 408.170 0.000 408.490 221.080 ;
 END
 PORT
  LAYER ME4 ;
  RECT 410.670 0.810 410.990 221.080 ;
 END
 PORT
  LAYER ME4 ;
  RECT 411.470 0.000 411.790 221.080 ;
 END
 PORT
  LAYER ME4 ;
  RECT 408.970 21.610 409.290 221.080 ;
 END
 PORT
  LAYER ME4 ;
  RECT 412.270 0.000 412.590 221.080 ;
 END
 PORT
  LAYER ME4 ;
  RECT 414.770 0.000 415.090 221.080 ;
 END
 PORT
  LAYER ME4 ;
  RECT 417.270 0.810 417.590 221.080 ;
 END
 PORT
  LAYER ME4 ;
  RECT 418.070 0.000 418.390 221.080 ;
 END
 PORT
  LAYER ME4 ;
  RECT 415.570 21.610 415.890 221.080 ;
 END
 PORT
  LAYER ME4 ;
  RECT 418.870 0.940 419.190 221.080 ;
 END
 PORT
  LAYER ME4 ;
  RECT 421.370 0.000 421.690 221.080 ;
 END
 PORT
  LAYER ME4 ;
  RECT 423.870 0.940 424.190 221.080 ;
 END
 PORT
  LAYER ME4 ;
  RECT 424.670 0.000 424.990 221.080 ;
 END
 PORT
  LAYER ME4 ;
  RECT 422.170 21.610 422.490 221.080 ;
 END
 PORT
  LAYER ME4 ;
  RECT 425.470 0.000 425.790 221.080 ;
 END
 PORT
  LAYER ME4 ;
  RECT 427.970 0.000 428.290 221.080 ;
 END
 PORT
  LAYER ME4 ;
  RECT 430.470 0.810 430.790 221.080 ;
 END
 PORT
  LAYER ME4 ;
  RECT 431.270 0.000 431.590 221.080 ;
 END
 PORT
  LAYER ME4 ;
  RECT 428.770 21.610 429.090 221.080 ;
 END
 PORT
  LAYER ME4 ;
  RECT 432.070 0.000 432.390 221.080 ;
 END
 PORT
  LAYER ME4 ;
  RECT 434.570 0.000 434.890 221.080 ;
 END
 PORT
  LAYER ME4 ;
  RECT 437.070 0.810 437.390 221.080 ;
 END
 PORT
  LAYER ME4 ;
  RECT 437.870 0.000 438.190 221.080 ;
 END
 PORT
  LAYER ME4 ;
  RECT 435.370 21.610 435.690 221.080 ;
 END
 PORT
  LAYER ME4 ;
  RECT 438.670 0.000 438.990 221.080 ;
 END
 PORT
  LAYER ME4 ;
  RECT 441.170 0.000 441.490 221.080 ;
 END
 PORT
  LAYER ME4 ;
  RECT 443.670 0.810 443.990 221.080 ;
 END
 PORT
  LAYER ME4 ;
  RECT 444.470 0.000 444.790 221.080 ;
 END
 PORT
  LAYER ME4 ;
  RECT 441.970 21.610 442.290 221.080 ;
 END
 PORT
  LAYER ME4 ;
  RECT 445.270 0.000 445.590 221.080 ;
 END
 PORT
  LAYER ME4 ;
  RECT 447.770 0.000 448.090 221.080 ;
 END
 PORT
  LAYER ME4 ;
  RECT 450.270 0.810 450.590 221.080 ;
 END
 PORT
  LAYER ME4 ;
  RECT 451.070 0.000 451.390 221.080 ;
 END
 PORT
  LAYER ME4 ;
  RECT 448.570 21.610 448.890 221.080 ;
 END
 PORT
  LAYER ME4 ;
  RECT 451.870 0.000 452.190 221.080 ;
 END
 PORT
  LAYER ME4 ;
  RECT 454.370 0.000 454.690 221.080 ;
 END
 PORT
  LAYER ME4 ;
  RECT 456.870 0.810 457.190 221.080 ;
 END
 PORT
  LAYER ME4 ;
  RECT 457.670 0.000 457.990 221.080 ;
 END
 PORT
  LAYER ME4 ;
  RECT 455.170 21.610 455.490 221.080 ;
 END
 PORT
  LAYER ME4 ;
  RECT 458.470 0.000 458.790 221.080 ;
 END
 PORT
  LAYER ME4 ;
  RECT 460.970 0.000 461.290 221.080 ;
 END
 PORT
  LAYER ME4 ;
  RECT 463.470 0.810 463.790 221.080 ;
 END
 PORT
  LAYER ME4 ;
  RECT 464.270 0.000 464.590 221.080 ;
 END
 PORT
  LAYER ME4 ;
  RECT 461.770 21.610 462.090 221.080 ;
 END
 PORT
  LAYER ME4 ;
  RECT 465.070 0.000 465.390 221.080 ;
 END
 PORT
  LAYER ME4 ;
  RECT 467.570 0.000 467.890 221.080 ;
 END
 PORT
  LAYER ME4 ;
  RECT 470.070 0.810 470.390 221.080 ;
 END
 PORT
  LAYER ME4 ;
  RECT 470.870 0.000 471.190 221.080 ;
 END
 PORT
  LAYER ME4 ;
  RECT 468.370 21.610 468.690 221.080 ;
 END
 PORT
  LAYER ME4 ;
  RECT 471.670 0.000 471.990 221.080 ;
 END
 PORT
  LAYER ME4 ;
  RECT 474.170 0.000 474.490 221.080 ;
 END
 PORT
  LAYER ME4 ;
  RECT 476.670 0.810 476.990 221.080 ;
 END
 PORT
  LAYER ME4 ;
  RECT 477.470 0.000 477.790 221.080 ;
 END
 PORT
  LAYER ME4 ;
  RECT 474.970 21.610 475.290 221.080 ;
 END
 PORT
  LAYER ME4 ;
  RECT 478.270 0.940 478.590 221.080 ;
 END
 PORT
  LAYER ME4 ;
  RECT 480.770 0.000 481.090 221.080 ;
 END
 PORT
  LAYER ME4 ;
  RECT 483.270 0.940 483.590 221.080 ;
 END
 PORT
  LAYER ME4 ;
  RECT 484.070 0.000 484.390 221.080 ;
 END
 PORT
  LAYER ME4 ;
  RECT 481.570 21.610 481.890 221.080 ;
 END
 PORT
  LAYER ME4 ;
  RECT 484.870 0.000 485.190 221.080 ;
 END
 PORT
  LAYER ME4 ;
  RECT 487.370 0.000 487.690 221.080 ;
 END
 PORT
  LAYER ME4 ;
  RECT 489.870 0.810 490.190 221.080 ;
 END
 PORT
  LAYER ME4 ;
  RECT 490.670 0.000 490.990 221.080 ;
 END
 PORT
  LAYER ME4 ;
  RECT 488.170 21.610 488.490 221.080 ;
 END
 PORT
  LAYER ME4 ;
  RECT 491.470 0.000 491.790 221.080 ;
 END
 PORT
  LAYER ME4 ;
  RECT 493.970 0.000 494.290 221.080 ;
 END
 PORT
  LAYER ME4 ;
  RECT 496.470 0.810 496.790 221.080 ;
 END
 PORT
  LAYER ME4 ;
  RECT 497.270 0.000 497.590 221.080 ;
 END
 PORT
  LAYER ME4 ;
  RECT 494.770 21.610 495.090 221.080 ;
 END
 PORT
  LAYER ME4 ;
  RECT 498.070 0.000 498.390 221.080 ;
 END
 PORT
  LAYER ME4 ;
  RECT 500.570 0.000 500.890 221.080 ;
 END
 PORT
  LAYER ME4 ;
  RECT 503.070 0.810 503.390 221.080 ;
 END
 PORT
  LAYER ME4 ;
  RECT 503.870 0.000 504.190 221.080 ;
 END
 PORT
  LAYER ME4 ;
  RECT 501.370 21.610 501.690 221.080 ;
 END
 PORT
  LAYER ME4 ;
  RECT 504.670 0.000 504.990 221.080 ;
 END
 PORT
  LAYER ME4 ;
  RECT 507.170 0.000 507.490 221.080 ;
 END
 PORT
  LAYER ME4 ;
  RECT 509.670 0.810 509.990 221.080 ;
 END
 PORT
  LAYER ME4 ;
  RECT 510.470 0.000 510.790 221.080 ;
 END
 PORT
  LAYER ME4 ;
  RECT 507.970 21.610 508.290 221.080 ;
 END
 PORT
  LAYER ME4 ;
  RECT 511.270 0.000 511.590 221.080 ;
 END
 PORT
  LAYER ME4 ;
  RECT 513.770 0.000 514.090 221.080 ;
 END
 PORT
  LAYER ME4 ;
  RECT 516.270 0.810 516.590 221.080 ;
 END
 PORT
  LAYER ME4 ;
  RECT 517.070 0.000 517.390 221.080 ;
 END
 PORT
  LAYER ME4 ;
  RECT 514.570 21.610 514.890 221.080 ;
 END
 PORT
  LAYER ME4 ;
  RECT 517.870 0.000 518.190 221.080 ;
 END
 PORT
  LAYER ME4 ;
  RECT 520.370 0.000 520.690 221.080 ;
 END
 PORT
  LAYER ME4 ;
  RECT 522.870 0.810 523.190 221.080 ;
 END
 PORT
  LAYER ME4 ;
  RECT 523.670 0.000 523.990 221.080 ;
 END
 PORT
  LAYER ME4 ;
  RECT 521.170 21.610 521.490 221.080 ;
 END
 PORT
  LAYER ME4 ;
  RECT 524.470 0.000 524.790 221.080 ;
 END
 PORT
  LAYER ME4 ;
  RECT 526.970 0.000 527.290 221.080 ;
 END
 PORT
  LAYER ME4 ;
  RECT 529.470 0.810 529.790 221.080 ;
 END
 PORT
  LAYER ME4 ;
  RECT 530.270 0.000 530.590 221.080 ;
 END
 PORT
  LAYER ME4 ;
  RECT 527.770 21.610 528.090 221.080 ;
 END
 PORT
  LAYER ME4 ;
  RECT 531.070 0.000 531.390 221.080 ;
 END
 PORT
  LAYER ME4 ;
  RECT 533.570 0.000 533.890 221.080 ;
 END
 PORT
  LAYER ME4 ;
  RECT 536.070 0.810 536.390 221.080 ;
 END
 PORT
  LAYER ME4 ;
  RECT 536.870 0.000 537.190 221.080 ;
 END
 PORT
  LAYER ME4 ;
  RECT 534.370 21.610 534.690 221.080 ;
 END
 PORT
  LAYER ME4 ;
  RECT 537.670 192.316 538.000 221.080 ;
 END
 PORT
  LAYER ME4 ;
  RECT 298.470 0.800 298.790 221.080 ;
 END
 PORT
  LAYER ME4 ;
  RECT 295.970 0.800 296.290 221.080 ;
 END
 PORT
  LAYER ME4 ;
  RECT 295.170 0.800 295.490 195.270 ;
 END
 PORT
  LAYER ME4 ;
  RECT 291.860 0.000 292.190 221.080 ;
 END
 PORT
  LAYER ME4 ;
  RECT 293.470 0.800 293.790 221.080 ;
 END
 PORT
  LAYER ME4 ;
  RECT 292.670 0.000 292.990 221.080 ;
 END
 PORT
  LAYER ME4 ;
  RECT 296.770 21.610 297.090 221.080 ;
 END
 PORT
  LAYER ME4 ;
  RECT 301.770 0.000 302.090 195.270 ;
 END
 PORT
  LAYER ME4 ;
  RECT 308.370 0.000 308.690 195.270 ;
 END
 PORT
  LAYER ME4 ;
  RECT 314.970 0.000 315.290 195.270 ;
 END
 PORT
  LAYER ME4 ;
  RECT 321.570 0.000 321.890 195.270 ;
 END
 PORT
  LAYER ME4 ;
  RECT 328.170 0.000 328.490 195.270 ;
 END
 PORT
  LAYER ME4 ;
  RECT 334.770 0.000 335.090 195.270 ;
 END
 PORT
  LAYER ME4 ;
  RECT 341.370 0.000 341.690 195.270 ;
 END
 PORT
  LAYER ME4 ;
  RECT 347.970 0.000 348.290 195.270 ;
 END
 PORT
  LAYER ME4 ;
  RECT 354.570 0.000 354.890 195.270 ;
 END
 PORT
  LAYER ME4 ;
  RECT 361.170 0.000 361.490 195.270 ;
 END
 PORT
  LAYER ME4 ;
  RECT 367.770 0.000 368.090 195.270 ;
 END
 PORT
  LAYER ME4 ;
  RECT 374.370 0.000 374.690 195.270 ;
 END
 PORT
  LAYER ME4 ;
  RECT 380.970 0.000 381.290 195.270 ;
 END
 PORT
  LAYER ME4 ;
  RECT 387.570 0.000 387.890 195.270 ;
 END
 PORT
  LAYER ME4 ;
  RECT 394.170 0.000 394.490 195.270 ;
 END
 PORT
  LAYER ME4 ;
  RECT 400.770 0.000 401.090 195.270 ;
 END
 PORT
  LAYER ME4 ;
  RECT 407.370 0.000 407.690 195.270 ;
 END
 PORT
  LAYER ME4 ;
  RECT 413.970 0.000 414.290 195.270 ;
 END
 PORT
  LAYER ME4 ;
  RECT 420.570 0.000 420.890 195.270 ;
 END
 PORT
  LAYER ME4 ;
  RECT 427.170 0.000 427.490 195.270 ;
 END
 PORT
  LAYER ME4 ;
  RECT 433.770 0.000 434.090 195.270 ;
 END
 PORT
  LAYER ME4 ;
  RECT 440.370 0.000 440.690 195.270 ;
 END
 PORT
  LAYER ME4 ;
  RECT 446.970 0.000 447.290 195.270 ;
 END
 PORT
  LAYER ME4 ;
  RECT 453.570 0.000 453.890 195.270 ;
 END
 PORT
  LAYER ME4 ;
  RECT 460.170 0.000 460.490 195.270 ;
 END
 PORT
  LAYER ME4 ;
  RECT 466.770 0.000 467.090 195.270 ;
 END
 PORT
  LAYER ME4 ;
  RECT 473.370 0.000 473.690 195.270 ;
 END
 PORT
  LAYER ME4 ;
  RECT 479.970 0.000 480.290 195.270 ;
 END
 PORT
  LAYER ME4 ;
  RECT 486.570 0.000 486.890 195.270 ;
 END
 PORT
  LAYER ME4 ;
  RECT 493.170 0.000 493.490 195.270 ;
 END
 PORT
  LAYER ME4 ;
  RECT 499.770 0.000 500.090 195.270 ;
 END
 PORT
  LAYER ME4 ;
  RECT 506.370 0.000 506.690 195.270 ;
 END
 PORT
  LAYER ME4 ;
  RECT 512.970 0.000 513.290 195.270 ;
 END
 PORT
  LAYER ME4 ;
  RECT 519.570 0.000 519.890 195.270 ;
 END
 PORT
  LAYER ME4 ;
  RECT 526.170 0.000 526.490 195.270 ;
 END
 PORT
  LAYER ME4 ;
  RECT 532.770 0.000 533.090 195.270 ;
 END
 PORT
  LAYER ME4 ;
  RECT 537.670 24.565 538.000 192.315 ;
 END
 PORT
  LAYER ME4 ;
  RECT 537.670 0.000 538.000 24.564 ;
 END
 PORT
  LAYER ME4 ;
  RECT 1.250 0.000 1.580 221.080 ;
 END
 PORT
  LAYER ME4 ;
  RECT 2.860 0.940 3.180 221.080 ;
 END
 PORT
  LAYER ME4 ;
  RECT 2.060 0.000 2.380 221.080 ;
 END
 PORT
  LAYER ME4 ;
  RECT 5.360 0.000 5.680 221.080 ;
 END
 PORT
  LAYER ME4 ;
  RECT 7.860 0.940 8.180 221.080 ;
 END
 PORT
  LAYER ME4 ;
  RECT 8.660 0.000 8.980 221.080 ;
 END
 PORT
  LAYER ME4 ;
  RECT 6.160 21.610 6.480 221.080 ;
 END
 PORT
  LAYER ME4 ;
  RECT 9.460 0.000 9.780 221.080 ;
 END
 PORT
  LAYER ME4 ;
  RECT 11.960 0.000 12.280 221.080 ;
 END
 PORT
  LAYER ME4 ;
  RECT 14.460 0.810 14.780 221.080 ;
 END
 PORT
  LAYER ME4 ;
  RECT 15.260 0.000 15.580 221.080 ;
 END
 PORT
  LAYER ME4 ;
  RECT 12.760 21.610 13.080 221.080 ;
 END
 PORT
  LAYER ME4 ;
  RECT 16.060 0.000 16.380 221.080 ;
 END
 PORT
  LAYER ME4 ;
  RECT 18.560 0.000 18.880 221.080 ;
 END
 PORT
  LAYER ME4 ;
  RECT 21.060 0.810 21.380 221.080 ;
 END
 PORT
  LAYER ME4 ;
  RECT 21.860 0.000 22.180 221.080 ;
 END
 PORT
  LAYER ME4 ;
  RECT 19.360 21.610 19.680 221.080 ;
 END
 PORT
  LAYER ME4 ;
  RECT 22.660 0.000 22.980 221.080 ;
 END
 PORT
  LAYER ME4 ;
  RECT 25.160 0.000 25.480 221.080 ;
 END
 PORT
  LAYER ME4 ;
  RECT 27.660 0.810 27.980 221.080 ;
 END
 PORT
  LAYER ME4 ;
  RECT 28.460 0.000 28.780 221.080 ;
 END
 PORT
  LAYER ME4 ;
  RECT 25.960 21.610 26.280 221.080 ;
 END
 PORT
  LAYER ME4 ;
  RECT 29.260 0.000 29.580 221.080 ;
 END
 PORT
  LAYER ME4 ;
  RECT 31.760 0.000 32.080 221.080 ;
 END
 PORT
  LAYER ME4 ;
  RECT 34.260 0.810 34.580 221.080 ;
 END
 PORT
  LAYER ME4 ;
  RECT 35.060 0.000 35.380 221.080 ;
 END
 PORT
  LAYER ME4 ;
  RECT 32.560 21.610 32.880 221.080 ;
 END
 PORT
  LAYER ME4 ;
  RECT 35.860 0.000 36.180 221.080 ;
 END
 PORT
  LAYER ME4 ;
  RECT 38.360 0.000 38.680 221.080 ;
 END
 PORT
  LAYER ME4 ;
  RECT 40.860 0.810 41.180 221.080 ;
 END
 PORT
  LAYER ME4 ;
  RECT 41.660 0.000 41.980 221.080 ;
 END
 PORT
  LAYER ME4 ;
  RECT 39.160 21.610 39.480 221.080 ;
 END
 PORT
  LAYER ME4 ;
  RECT 42.460 0.000 42.780 221.080 ;
 END
 PORT
  LAYER ME4 ;
  RECT 44.960 0.000 45.280 221.080 ;
 END
 PORT
  LAYER ME4 ;
  RECT 47.460 0.810 47.780 221.080 ;
 END
 PORT
  LAYER ME4 ;
  RECT 48.260 0.000 48.580 221.080 ;
 END
 PORT
  LAYER ME4 ;
  RECT 45.760 21.610 46.080 221.080 ;
 END
 PORT
  LAYER ME4 ;
  RECT 49.060 0.000 49.380 221.080 ;
 END
 PORT
  LAYER ME4 ;
  RECT 51.560 0.000 51.880 221.080 ;
 END
 PORT
  LAYER ME4 ;
  RECT 54.060 0.810 54.380 221.080 ;
 END
 PORT
  LAYER ME4 ;
  RECT 54.860 0.000 55.180 221.080 ;
 END
 PORT
  LAYER ME4 ;
  RECT 52.360 21.610 52.680 221.080 ;
 END
 PORT
  LAYER ME4 ;
  RECT 55.660 0.000 55.980 221.080 ;
 END
 PORT
  LAYER ME4 ;
  RECT 58.160 0.000 58.480 221.080 ;
 END
 PORT
  LAYER ME4 ;
  RECT 60.660 0.810 60.980 221.080 ;
 END
 PORT
  LAYER ME4 ;
  RECT 61.460 0.000 61.780 221.080 ;
 END
 PORT
  LAYER ME4 ;
  RECT 58.960 21.610 59.280 221.080 ;
 END
 PORT
  LAYER ME4 ;
  RECT 62.260 0.940 62.580 221.080 ;
 END
 PORT
  LAYER ME4 ;
  RECT 64.760 0.000 65.080 221.080 ;
 END
 PORT
  LAYER ME4 ;
  RECT 67.260 0.940 67.580 221.080 ;
 END
 PORT
  LAYER ME4 ;
  RECT 68.060 0.000 68.380 221.080 ;
 END
 PORT
  LAYER ME4 ;
  RECT 65.560 21.610 65.880 221.080 ;
 END
 PORT
  LAYER ME4 ;
  RECT 68.860 0.000 69.180 221.080 ;
 END
 PORT
  LAYER ME4 ;
  RECT 71.360 0.000 71.680 221.080 ;
 END
 PORT
  LAYER ME4 ;
  RECT 73.860 0.810 74.180 221.080 ;
 END
 PORT
  LAYER ME4 ;
  RECT 74.660 0.000 74.980 221.080 ;
 END
 PORT
  LAYER ME4 ;
  RECT 72.160 21.610 72.480 221.080 ;
 END
 PORT
  LAYER ME4 ;
  RECT 75.460 0.000 75.780 221.080 ;
 END
 PORT
  LAYER ME4 ;
  RECT 77.960 0.000 78.280 221.080 ;
 END
 PORT
  LAYER ME4 ;
  RECT 80.460 0.810 80.780 221.080 ;
 END
 PORT
  LAYER ME4 ;
  RECT 81.260 0.000 81.580 221.080 ;
 END
 PORT
  LAYER ME4 ;
  RECT 78.760 21.610 79.080 221.080 ;
 END
 PORT
  LAYER ME4 ;
  RECT 82.060 0.000 82.380 221.080 ;
 END
 PORT
  LAYER ME4 ;
  RECT 84.560 0.000 84.880 221.080 ;
 END
 PORT
  LAYER ME4 ;
  RECT 87.060 0.810 87.380 221.080 ;
 END
 PORT
  LAYER ME4 ;
  RECT 87.860 0.000 88.180 221.080 ;
 END
 PORT
  LAYER ME4 ;
  RECT 85.360 21.610 85.680 221.080 ;
 END
 PORT
  LAYER ME4 ;
  RECT 88.660 0.000 88.980 221.080 ;
 END
 PORT
  LAYER ME4 ;
  RECT 91.160 0.000 91.480 221.080 ;
 END
 PORT
  LAYER ME4 ;
  RECT 93.660 0.810 93.980 221.080 ;
 END
 PORT
  LAYER ME4 ;
  RECT 94.460 0.000 94.780 221.080 ;
 END
 PORT
  LAYER ME4 ;
  RECT 91.960 21.610 92.280 221.080 ;
 END
 PORT
  LAYER ME4 ;
  RECT 95.260 0.000 95.580 221.080 ;
 END
 PORT
  LAYER ME4 ;
  RECT 97.760 0.000 98.080 221.080 ;
 END
 PORT
  LAYER ME4 ;
  RECT 100.260 0.810 100.580 221.080 ;
 END
 PORT
  LAYER ME4 ;
  RECT 101.060 0.000 101.380 221.080 ;
 END
 PORT
  LAYER ME4 ;
  RECT 98.560 21.610 98.880 221.080 ;
 END
 PORT
  LAYER ME4 ;
  RECT 101.860 0.000 102.180 221.080 ;
 END
 PORT
  LAYER ME4 ;
  RECT 104.360 0.000 104.680 221.080 ;
 END
 PORT
  LAYER ME4 ;
  RECT 106.860 0.810 107.180 221.080 ;
 END
 PORT
  LAYER ME4 ;
  RECT 107.660 0.000 107.980 221.080 ;
 END
 PORT
  LAYER ME4 ;
  RECT 105.160 21.610 105.480 221.080 ;
 END
 PORT
  LAYER ME4 ;
  RECT 108.460 0.000 108.780 221.080 ;
 END
 PORT
  LAYER ME4 ;
  RECT 110.960 0.000 111.280 221.080 ;
 END
 PORT
  LAYER ME4 ;
  RECT 113.460 0.810 113.780 221.080 ;
 END
 PORT
  LAYER ME4 ;
  RECT 114.260 0.000 114.580 221.080 ;
 END
 PORT
  LAYER ME4 ;
  RECT 111.760 21.610 112.080 221.080 ;
 END
 PORT
  LAYER ME4 ;
  RECT 115.060 0.000 115.380 221.080 ;
 END
 PORT
  LAYER ME4 ;
  RECT 117.560 0.000 117.880 221.080 ;
 END
 PORT
  LAYER ME4 ;
  RECT 120.060 0.810 120.380 221.080 ;
 END
 PORT
  LAYER ME4 ;
  RECT 120.860 0.000 121.180 221.080 ;
 END
 PORT
  LAYER ME4 ;
  RECT 118.360 21.610 118.680 221.080 ;
 END
 PORT
  LAYER ME4 ;
  RECT 121.660 0.940 121.980 221.080 ;
 END
 PORT
  LAYER ME4 ;
  RECT 124.160 0.000 124.480 221.080 ;
 END
 PORT
  LAYER ME4 ;
  RECT 126.660 0.940 126.980 221.080 ;
 END
 PORT
  LAYER ME4 ;
  RECT 127.460 0.000 127.780 221.080 ;
 END
 PORT
  LAYER ME4 ;
  RECT 124.960 21.610 125.280 221.080 ;
 END
 PORT
  LAYER ME4 ;
  RECT 128.260 0.000 128.580 221.080 ;
 END
 PORT
  LAYER ME4 ;
  RECT 130.760 0.000 131.080 221.080 ;
 END
 PORT
  LAYER ME4 ;
  RECT 133.260 0.810 133.580 221.080 ;
 END
 PORT
  LAYER ME4 ;
  RECT 134.060 0.000 134.380 221.080 ;
 END
 PORT
  LAYER ME4 ;
  RECT 131.560 21.610 131.880 221.080 ;
 END
 PORT
  LAYER ME4 ;
  RECT 134.860 0.000 135.180 221.080 ;
 END
 PORT
  LAYER ME4 ;
  RECT 137.360 0.000 137.680 221.080 ;
 END
 PORT
  LAYER ME4 ;
  RECT 139.860 0.810 140.180 221.080 ;
 END
 PORT
  LAYER ME4 ;
  RECT 140.660 0.000 140.980 221.080 ;
 END
 PORT
  LAYER ME4 ;
  RECT 138.160 21.610 138.480 221.080 ;
 END
 PORT
  LAYER ME4 ;
  RECT 141.460 0.000 141.780 221.080 ;
 END
 PORT
  LAYER ME4 ;
  RECT 143.960 0.000 144.280 221.080 ;
 END
 PORT
  LAYER ME4 ;
  RECT 146.460 0.810 146.780 221.080 ;
 END
 PORT
  LAYER ME4 ;
  RECT 147.260 0.000 147.580 221.080 ;
 END
 PORT
  LAYER ME4 ;
  RECT 144.760 21.610 145.080 221.080 ;
 END
 PORT
  LAYER ME4 ;
  RECT 148.060 0.000 148.380 221.080 ;
 END
 PORT
  LAYER ME4 ;
  RECT 150.560 0.000 150.880 221.080 ;
 END
 PORT
  LAYER ME4 ;
  RECT 153.060 0.810 153.380 221.080 ;
 END
 PORT
  LAYER ME4 ;
  RECT 153.860 0.000 154.180 221.080 ;
 END
 PORT
  LAYER ME4 ;
  RECT 151.360 21.610 151.680 221.080 ;
 END
 PORT
  LAYER ME4 ;
  RECT 154.660 0.000 154.980 221.080 ;
 END
 PORT
  LAYER ME4 ;
  RECT 157.160 0.000 157.480 221.080 ;
 END
 PORT
  LAYER ME4 ;
  RECT 159.660 0.810 159.980 221.080 ;
 END
 PORT
  LAYER ME4 ;
  RECT 160.460 0.000 160.780 221.080 ;
 END
 PORT
  LAYER ME4 ;
  RECT 157.960 21.610 158.280 221.080 ;
 END
 PORT
  LAYER ME4 ;
  RECT 161.260 0.000 161.580 221.080 ;
 END
 PORT
  LAYER ME4 ;
  RECT 163.760 0.000 164.080 221.080 ;
 END
 PORT
  LAYER ME4 ;
  RECT 166.260 0.810 166.580 221.080 ;
 END
 PORT
  LAYER ME4 ;
  RECT 167.060 0.000 167.380 221.080 ;
 END
 PORT
  LAYER ME4 ;
  RECT 164.560 21.610 164.880 221.080 ;
 END
 PORT
  LAYER ME4 ;
  RECT 167.860 0.000 168.180 221.080 ;
 END
 PORT
  LAYER ME4 ;
  RECT 170.360 0.000 170.680 221.080 ;
 END
 PORT
  LAYER ME4 ;
  RECT 172.860 0.810 173.180 221.080 ;
 END
 PORT
  LAYER ME4 ;
  RECT 173.660 0.000 173.980 221.080 ;
 END
 PORT
  LAYER ME4 ;
  RECT 171.160 21.610 171.480 221.080 ;
 END
 PORT
  LAYER ME4 ;
  RECT 174.460 0.000 174.780 221.080 ;
 END
 PORT
  LAYER ME4 ;
  RECT 176.960 0.000 177.280 221.080 ;
 END
 PORT
  LAYER ME4 ;
  RECT 179.460 0.810 179.780 221.080 ;
 END
 PORT
  LAYER ME4 ;
  RECT 180.260 0.000 180.580 221.080 ;
 END
 PORT
  LAYER ME4 ;
  RECT 177.760 21.610 178.080 221.080 ;
 END
 PORT
  LAYER ME4 ;
  RECT 181.060 0.940 181.380 221.080 ;
 END
 PORT
  LAYER ME4 ;
  RECT 183.560 0.000 183.880 221.080 ;
 END
 PORT
  LAYER ME4 ;
  RECT 186.060 0.940 186.380 221.080 ;
 END
 PORT
  LAYER ME4 ;
  RECT 186.860 0.000 187.180 221.080 ;
 END
 PORT
  LAYER ME4 ;
  RECT 184.360 21.610 184.680 221.080 ;
 END
 PORT
  LAYER ME4 ;
  RECT 187.660 0.000 187.980 221.080 ;
 END
 PORT
  LAYER ME4 ;
  RECT 190.160 0.000 190.480 221.080 ;
 END
 PORT
  LAYER ME4 ;
  RECT 192.660 0.810 192.980 221.080 ;
 END
 PORT
  LAYER ME4 ;
  RECT 193.460 0.000 193.780 221.080 ;
 END
 PORT
  LAYER ME4 ;
  RECT 190.960 21.610 191.280 221.080 ;
 END
 PORT
  LAYER ME4 ;
  RECT 194.260 0.000 194.580 221.080 ;
 END
 PORT
  LAYER ME4 ;
  RECT 196.760 0.000 197.080 221.080 ;
 END
 PORT
  LAYER ME4 ;
  RECT 199.260 0.810 199.580 221.080 ;
 END
 PORT
  LAYER ME4 ;
  RECT 200.060 0.000 200.380 221.080 ;
 END
 PORT
  LAYER ME4 ;
  RECT 197.560 21.610 197.880 221.080 ;
 END
 PORT
  LAYER ME4 ;
  RECT 200.860 0.000 201.180 221.080 ;
 END
 PORT
  LAYER ME4 ;
  RECT 203.360 0.000 203.680 221.080 ;
 END
 PORT
  LAYER ME4 ;
  RECT 205.860 0.810 206.180 221.080 ;
 END
 PORT
  LAYER ME4 ;
  RECT 206.660 0.000 206.980 221.080 ;
 END
 PORT
  LAYER ME4 ;
  RECT 204.160 21.610 204.480 221.080 ;
 END
 PORT
  LAYER ME4 ;
  RECT 207.460 0.000 207.780 221.080 ;
 END
 PORT
  LAYER ME4 ;
  RECT 209.960 0.000 210.280 221.080 ;
 END
 PORT
  LAYER ME4 ;
  RECT 212.460 0.810 212.780 221.080 ;
 END
 PORT
  LAYER ME4 ;
  RECT 213.260 0.000 213.580 221.080 ;
 END
 PORT
  LAYER ME4 ;
  RECT 210.760 21.610 211.080 221.080 ;
 END
 PORT
  LAYER ME4 ;
  RECT 214.060 0.000 214.380 221.080 ;
 END
 PORT
  LAYER ME4 ;
  RECT 216.560 0.000 216.880 221.080 ;
 END
 PORT
  LAYER ME4 ;
  RECT 219.060 0.810 219.380 221.080 ;
 END
 PORT
  LAYER ME4 ;
  RECT 219.860 0.000 220.180 221.080 ;
 END
 PORT
  LAYER ME4 ;
  RECT 217.360 21.610 217.680 221.080 ;
 END
 PORT
  LAYER ME4 ;
  RECT 220.660 0.000 220.980 221.080 ;
 END
 PORT
  LAYER ME4 ;
  RECT 223.160 0.000 223.480 221.080 ;
 END
 PORT
  LAYER ME4 ;
  RECT 225.660 0.810 225.980 221.080 ;
 END
 PORT
  LAYER ME4 ;
  RECT 226.460 0.000 226.780 221.080 ;
 END
 PORT
  LAYER ME4 ;
  RECT 223.960 21.610 224.280 221.080 ;
 END
 PORT
  LAYER ME4 ;
  RECT 227.260 0.000 227.580 221.080 ;
 END
 PORT
  LAYER ME4 ;
  RECT 229.760 0.000 230.080 221.080 ;
 END
 PORT
  LAYER ME4 ;
  RECT 232.260 0.810 232.580 221.080 ;
 END
 PORT
  LAYER ME4 ;
  RECT 233.060 0.000 233.380 221.080 ;
 END
 PORT
  LAYER ME4 ;
  RECT 230.560 21.610 230.880 221.080 ;
 END
 PORT
  LAYER ME4 ;
  RECT 233.860 0.000 234.180 221.080 ;
 END
 PORT
  LAYER ME4 ;
  RECT 236.360 0.000 236.680 221.080 ;
 END
 PORT
  LAYER ME4 ;
  RECT 238.860 0.810 239.180 221.080 ;
 END
 PORT
  LAYER ME4 ;
  RECT 239.660 0.000 239.980 221.080 ;
 END
 PORT
  LAYER ME4 ;
  RECT 237.160 21.610 237.480 221.080 ;
 END
 PORT
  LAYER ME4 ;
  RECT 240.460 0.000 240.790 221.080 ;
 END
 PORT
  LAYER ME4 ;
  RECT 4.560 0.000 4.880 195.270 ;
 END
 PORT
  LAYER ME4 ;
  RECT 11.160 0.000 11.480 195.270 ;
 END
 PORT
  LAYER ME4 ;
  RECT 17.760 0.000 18.080 195.270 ;
 END
 PORT
  LAYER ME4 ;
  RECT 24.360 0.000 24.680 195.270 ;
 END
 PORT
  LAYER ME4 ;
  RECT 30.960 0.000 31.280 195.270 ;
 END
 PORT
  LAYER ME4 ;
  RECT 37.560 0.000 37.880 195.270 ;
 END
 PORT
  LAYER ME4 ;
  RECT 44.160 0.000 44.480 195.270 ;
 END
 PORT
  LAYER ME4 ;
  RECT 50.760 0.000 51.080 195.270 ;
 END
 PORT
  LAYER ME4 ;
  RECT 57.360 0.000 57.680 195.270 ;
 END
 PORT
  LAYER ME4 ;
  RECT 63.960 0.000 64.280 195.270 ;
 END
 PORT
  LAYER ME4 ;
  RECT 70.560 0.000 70.880 195.270 ;
 END
 PORT
  LAYER ME4 ;
  RECT 77.160 0.000 77.480 195.270 ;
 END
 PORT
  LAYER ME4 ;
  RECT 83.760 0.000 84.080 195.270 ;
 END
 PORT
  LAYER ME4 ;
  RECT 90.360 0.000 90.680 195.270 ;
 END
 PORT
  LAYER ME4 ;
  RECT 96.960 0.000 97.280 195.270 ;
 END
 PORT
  LAYER ME4 ;
  RECT 103.560 0.000 103.880 195.270 ;
 END
 PORT
  LAYER ME4 ;
  RECT 110.160 0.000 110.480 195.270 ;
 END
 PORT
  LAYER ME4 ;
  RECT 116.760 0.000 117.080 195.270 ;
 END
 PORT
  LAYER ME4 ;
  RECT 123.360 0.000 123.680 195.270 ;
 END
 PORT
  LAYER ME4 ;
  RECT 129.960 0.000 130.280 195.270 ;
 END
 PORT
  LAYER ME4 ;
  RECT 136.560 0.000 136.880 195.270 ;
 END
 PORT
  LAYER ME4 ;
  RECT 143.160 0.000 143.480 195.270 ;
 END
 PORT
  LAYER ME4 ;
  RECT 149.760 0.000 150.080 195.270 ;
 END
 PORT
  LAYER ME4 ;
  RECT 156.360 0.000 156.680 195.270 ;
 END
 PORT
  LAYER ME4 ;
  RECT 162.960 0.000 163.280 195.270 ;
 END
 PORT
  LAYER ME4 ;
  RECT 169.560 0.000 169.880 195.270 ;
 END
 PORT
  LAYER ME4 ;
  RECT 176.160 0.000 176.480 195.270 ;
 END
 PORT
  LAYER ME4 ;
  RECT 182.760 0.000 183.080 195.270 ;
 END
 PORT
  LAYER ME4 ;
  RECT 189.360 0.000 189.680 195.270 ;
 END
 PORT
  LAYER ME4 ;
  RECT 195.960 0.000 196.280 195.270 ;
 END
 PORT
  LAYER ME4 ;
  RECT 202.560 0.000 202.880 195.270 ;
 END
 PORT
  LAYER ME4 ;
  RECT 209.160 0.000 209.480 195.270 ;
 END
 PORT
  LAYER ME4 ;
  RECT 215.760 0.000 216.080 195.270 ;
 END
 PORT
  LAYER ME4 ;
  RECT 222.360 0.000 222.680 195.270 ;
 END
 PORT
  LAYER ME4 ;
  RECT 228.960 0.000 229.280 195.270 ;
 END
 PORT
  LAYER ME4 ;
  RECT 235.560 0.000 235.880 195.270 ;
 END
 PORT
  LAYER ME4 ;
  RECT 267.220 195.270 267.820 221.080 ;
 END
 PORT
  LAYER ME4 ;
  RECT 269.420 0.000 270.020 221.080 ;
 END
 PORT
  LAYER ME4 ;
  RECT 271.620 0.000 272.220 221.080 ;
 END
 PORT
  LAYER ME4 ;
  RECT 273.820 0.000 274.420 221.080 ;
 END
 PORT
  LAYER ME4 ;
  RECT 276.020 0.000 276.620 220.250 ;
 END
 PORT
  LAYER ME4 ;
  RECT 278.220 0.000 278.820 221.080 ;
 END
 PORT
  LAYER ME4 ;
  RECT 280.645 197.080 281.245 221.080 ;
 END
 PORT
  LAYER ME4 ;
  RECT 283.070 0.000 283.670 221.080 ;
 END
 PORT
  LAYER ME4 ;
  RECT 285.270 0.000 285.870 221.080 ;
 END
 PORT
  LAYER ME4 ;
  RECT 288.570 0.000 289.170 221.080 ;
 END
 PORT
  LAYER ME4 ;
  RECT 289.670 0.000 290.270 221.080 ;
 END
 PORT
  LAYER ME4 ;
  RECT 262.570 0.000 263.170 221.080 ;
 END
 PORT
  LAYER ME4 ;
  RECT 264.770 195.270 265.370 221.080 ;
 END
 PORT
  LAYER ME4 ;
  RECT 258.170 195.270 258.770 221.080 ;
 END
 PORT
  LAYER ME4 ;
  RECT 255.970 195.270 256.570 221.080 ;
 END
 PORT
  LAYER ME4 ;
  RECT 260.370 0.800 260.970 220.250 ;
 END
 PORT
  LAYER ME4 ;
  RECT 251.810 195.270 252.410 221.080 ;
 END
 PORT
  LAYER ME4 ;
  RECT 249.610 195.270 250.210 221.080 ;
 END
 PORT
  LAYER ME4 ;
  RECT 254.010 195.270 254.610 220.250 ;
 END
 PORT
  LAYER ME4 ;
  RECT 245.450 195.270 246.050 221.080 ;
 END
 PORT
  LAYER ME4 ;
  RECT 243.250 195.270 243.850 221.080 ;
 END
 PORT
  LAYER ME4 ;
  RECT 247.650 195.270 248.250 220.250 ;
 END
 PORT
  LAYER ME4 ;
  RECT 267.220 0.000 267.820 21.610 ;
 END
 PORT
  LAYER ME4 ;
  RECT 280.870 0.000 281.470 21.610 ;
 END
 PORT
  LAYER ME4 ;
  RECT 264.770 0.000 265.370 21.700 ;
 END
 PORT
  LAYER ME4 ;
  RECT 255.970 0.000 256.570 21.700 ;
 END
 PORT
  LAYER ME4 ;
  RECT 258.170 0.000 258.770 21.700 ;
 END
 PORT
  LAYER ME4 ;
  RECT 249.610 0.000 250.210 21.700 ;
 END
 PORT
  LAYER ME4 ;
  RECT 251.810 0.000 252.410 21.700 ;
 END
 PORT
  LAYER ME4 ;
  RECT 254.010 0.800 254.610 21.700 ;
 END
 PORT
  LAYER ME4 ;
  RECT 243.250 0.000 243.850 21.700 ;
 END
 PORT
  LAYER ME4 ;
  RECT 245.450 0.000 246.050 21.700 ;
 END
 PORT
  LAYER ME4 ;
  RECT 247.650 0.800 248.250 21.700 ;
 END
END GND
PIN A7
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 244.050 220.480 244.370 221.080 ;
  LAYER ME3 ;
  RECT 244.050 220.480 244.370 221.080 ;
  LAYER ME2 ;
  RECT 244.050 220.480 244.370 221.080 ;
  LAYER ME1 ;
  RECT 244.050 220.480 244.370 221.080 ;
 END
 ANTENNAPARTIALMETALAREA                  2.030 LAYER ME2 ;
 ANTENNAGATEAREA                          0.216 LAYER ME2 ;
 ANTENNAGATEAREA                          0.216 LAYER ME3 ;
 ANTENNAGATEAREA                          0.216 LAYER ME4 ;
 ANTENNADIFFAREA                          0.160 LAYER ME2 ;
 ANTENNADIFFAREA                          0.160 LAYER ME3 ;
 ANTENNADIFFAREA                          0.160 LAYER ME4 ;
 ANTENNAMAXAREACAR                       11.826 LAYER ME2 ;
 ANTENNAMAXAREACAR                       12.715 LAYER ME3 ;
 ANTENNAMAXAREACAR                       13.604 LAYER ME4 ;
END A7
PIN A6
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 247.350 220.480 247.670 221.080 ;
  LAYER ME3 ;
  RECT 247.350 220.480 247.670 221.080 ;
  LAYER ME2 ;
  RECT 247.350 220.480 247.670 221.080 ;
  LAYER ME1 ;
  RECT 247.350 220.480 247.670 221.080 ;
 END
 ANTENNAPARTIALMETALAREA                  1.478 LAYER ME2 ;
 ANTENNAGATEAREA                          0.216 LAYER ME2 ;
 ANTENNAGATEAREA                          0.216 LAYER ME3 ;
 ANTENNAGATEAREA                          0.216 LAYER ME4 ;
 ANTENNADIFFAREA                          0.160 LAYER ME2 ;
 ANTENNADIFFAREA                          0.160 LAYER ME3 ;
 ANTENNADIFFAREA                          0.160 LAYER ME4 ;
 ANTENNAMAXAREACAR                        9.307 LAYER ME2 ;
 ANTENNAMAXAREACAR                       10.196 LAYER ME3 ;
 ANTENNAMAXAREACAR                       11.085 LAYER ME4 ;
END A6
PIN A5
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 250.410 220.480 250.730 221.080 ;
  LAYER ME3 ;
  RECT 250.410 220.480 250.730 221.080 ;
  LAYER ME2 ;
  RECT 250.410 220.480 250.730 221.080 ;
  LAYER ME1 ;
  RECT 250.410 220.480 250.730 221.080 ;
 END
 ANTENNAPARTIALMETALAREA                  2.030 LAYER ME2 ;
 ANTENNAGATEAREA                          0.216 LAYER ME2 ;
 ANTENNAGATEAREA                          0.216 LAYER ME3 ;
 ANTENNAGATEAREA                          0.216 LAYER ME4 ;
 ANTENNADIFFAREA                          0.160 LAYER ME2 ;
 ANTENNADIFFAREA                          0.160 LAYER ME3 ;
 ANTENNADIFFAREA                          0.160 LAYER ME4 ;
 ANTENNAMAXAREACAR                       11.826 LAYER ME2 ;
 ANTENNAMAXAREACAR                       12.715 LAYER ME3 ;
 ANTENNAMAXAREACAR                       13.604 LAYER ME4 ;
END A5
PIN A4
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 253.710 220.480 254.030 221.080 ;
  LAYER ME3 ;
  RECT 253.710 220.480 254.030 221.080 ;
  LAYER ME2 ;
  RECT 253.710 220.480 254.030 221.080 ;
  LAYER ME1 ;
  RECT 253.710 220.480 254.030 221.080 ;
 END
 ANTENNAPARTIALMETALAREA                  1.478 LAYER ME2 ;
 ANTENNAGATEAREA                          0.216 LAYER ME2 ;
 ANTENNAGATEAREA                          0.216 LAYER ME3 ;
 ANTENNAGATEAREA                          0.216 LAYER ME4 ;
 ANTENNADIFFAREA                          0.160 LAYER ME2 ;
 ANTENNADIFFAREA                          0.160 LAYER ME3 ;
 ANTENNADIFFAREA                          0.160 LAYER ME4 ;
 ANTENNAMAXAREACAR                        9.307 LAYER ME2 ;
 ANTENNAMAXAREACAR                       10.196 LAYER ME3 ;
 ANTENNAMAXAREACAR                       11.085 LAYER ME4 ;
END A4
PIN A3
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 256.770 220.480 257.090 221.080 ;
  LAYER ME3 ;
  RECT 256.770 220.480 257.090 221.080 ;
  LAYER ME2 ;
  RECT 256.770 220.480 257.090 221.080 ;
  LAYER ME1 ;
  RECT 256.770 220.480 257.090 221.080 ;
 END
 ANTENNAPARTIALMETALAREA                  2.030 LAYER ME2 ;
 ANTENNAGATEAREA                          0.216 LAYER ME2 ;
 ANTENNAGATEAREA                          0.216 LAYER ME3 ;
 ANTENNAGATEAREA                          0.216 LAYER ME4 ;
 ANTENNADIFFAREA                          0.160 LAYER ME2 ;
 ANTENNADIFFAREA                          0.160 LAYER ME3 ;
 ANTENNADIFFAREA                          0.160 LAYER ME4 ;
 ANTENNAMAXAREACAR                       11.826 LAYER ME2 ;
 ANTENNAMAXAREACAR                       12.715 LAYER ME3 ;
 ANTENNAMAXAREACAR                       13.604 LAYER ME4 ;
END A3
PIN A2
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 260.070 220.480 260.390 221.080 ;
  LAYER ME3 ;
  RECT 260.070 220.480 260.390 221.080 ;
  LAYER ME2 ;
  RECT 260.070 220.480 260.390 221.080 ;
  LAYER ME1 ;
  RECT 260.070 220.480 260.390 221.080 ;
 END
 ANTENNAPARTIALMETALAREA                  1.478 LAYER ME2 ;
 ANTENNAGATEAREA                          0.216 LAYER ME2 ;
 ANTENNAGATEAREA                          0.216 LAYER ME3 ;
 ANTENNAGATEAREA                          0.216 LAYER ME4 ;
 ANTENNADIFFAREA                          0.160 LAYER ME2 ;
 ANTENNADIFFAREA                          0.160 LAYER ME3 ;
 ANTENNADIFFAREA                          0.160 LAYER ME4 ;
 ANTENNAMAXAREACAR                        9.307 LAYER ME2 ;
 ANTENNAMAXAREACAR                       10.196 LAYER ME3 ;
 ANTENNAMAXAREACAR                       11.085 LAYER ME4 ;
END A2
PIN A1
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 270.220 220.480 270.540 221.080 ;
  LAYER ME3 ;
  RECT 270.220 220.480 270.540 221.080 ;
  LAYER ME2 ;
  RECT 270.220 220.480 270.540 221.080 ;
  LAYER ME1 ;
  RECT 270.220 220.480 270.540 221.080 ;
 END
 ANTENNAPARTIALMETALAREA                  1.366 LAYER ME2 ;
 ANTENNAGATEAREA                          0.216 LAYER ME2 ;
 ANTENNAGATEAREA                          0.216 LAYER ME3 ;
 ANTENNAGATEAREA                          0.216 LAYER ME4 ;
 ANTENNADIFFAREA                          0.160 LAYER ME2 ;
 ANTENNADIFFAREA                          0.160 LAYER ME3 ;
 ANTENNADIFFAREA                          0.160 LAYER ME4 ;
 ANTENNAMAXAREACAR                        9.176 LAYER ME2 ;
 ANTENNAMAXAREACAR                       10.065 LAYER ME3 ;
 ANTENNAMAXAREACAR                       10.954 LAYER ME4 ;
END A1
PIN A0
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 280.125 220.480 280.445 221.080 ;
  LAYER ME3 ;
  RECT 280.125 220.480 280.445 221.080 ;
  LAYER ME2 ;
  RECT 280.125 220.480 280.445 221.080 ;
  LAYER ME1 ;
  RECT 280.125 220.480 280.445 221.080 ;
 END
 ANTENNAPARTIALMETALAREA                  1.503 LAYER ME2 ;
 ANTENNAGATEAREA                          0.216 LAYER ME2 ;
 ANTENNAGATEAREA                          0.216 LAYER ME3 ;
 ANTENNAGATEAREA                          0.216 LAYER ME4 ;
 ANTENNADIFFAREA                          0.160 LAYER ME2 ;
 ANTENNADIFFAREA                          0.160 LAYER ME3 ;
 ANTENNADIFFAREA                          0.160 LAYER ME4 ;
 ANTENNAMAXAREACAR                        9.610 LAYER ME2 ;
 ANTENNAMAXAREACAR                       10.499 LAYER ME3 ;
 ANTENNAMAXAREACAR                       11.388 LAYER ME4 ;
END A0
PIN CSAN
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 275.720 220.480 276.040 221.080 ;
  LAYER ME3 ;
  RECT 275.720 220.480 276.040 221.080 ;
  LAYER ME2 ;
  RECT 275.720 220.480 276.040 221.080 ;
  LAYER ME1 ;
  RECT 275.720 220.480 276.040 221.080 ;
 END
 ANTENNAPARTIALMETALAREA                  2.236 LAYER ME2 ;
 ANTENNAPARTIALMETALAREA                  8.466 LAYER ME3 ;
 ANTENNAGATEAREA                          0.278 LAYER ME2 ;
 ANTENNAGATEAREA                          1.526 LAYER ME3 ;
 ANTENNAGATEAREA                          1.526 LAYER ME4 ;
 ANTENNADIFFAREA                          0.160 LAYER ME2 ;
 ANTENNADIFFAREA                          0.160 LAYER ME3 ;
 ANTENNADIFFAREA                          0.160 LAYER ME4 ;
 ANTENNAMAXAREACAR                        9.239 LAYER ME2 ;
 ANTENNAMAXAREACAR                       68.973 LAYER ME3 ;
 ANTENNAMAXAREACAR                       70.402 LAYER ME4 ;
END CSAN
PIN CKA
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 272.420 220.480 272.740 221.080 ;
  LAYER ME3 ;
  RECT 272.420 220.480 272.740 221.080 ;
  LAYER ME2 ;
  RECT 272.420 220.480 272.740 221.080 ;
  LAYER ME1 ;
  RECT 272.420 220.480 272.740 221.080 ;
 END
 ANTENNAPARTIALMETALAREA                  1.870 LAYER ME2 ;
 ANTENNAPARTIALMETALAREA                  8.466 LAYER ME3 ;
 ANTENNAGATEAREA                          1.632 LAYER ME3 ;
 ANTENNAGATEAREA                          1.632 LAYER ME4 ;
 ANTENNADIFFAREA                          0.160 LAYER ME2 ;
 ANTENNADIFFAREA                          0.160 LAYER ME3 ;
 ANTENNADIFFAREA                          0.160 LAYER ME4 ;
 ANTENNAMAXAREACAR                       38.858 LAYER ME3 ;
 ANTENNAMAXAREACAR                       39.658 LAYER ME4 ;
END CKA
PIN DO35
  DIRECTION OUTPUT ;
 PORT
  LAYER ME4 ;
  RECT 237.680 220.480 238.000 221.080 ;
  LAYER ME3 ;
  RECT 237.680 220.480 238.000 221.080 ;
  LAYER ME2 ;
  RECT 237.680 220.480 238.000 221.080 ;
  LAYER ME1 ;
  RECT 237.680 220.480 238.000 221.080 ;
 END
 ANTENNAPARTIALMETALAREA                  0.802 LAYER ME2 ;
 ANTENNADIFFAREA                          2.912 LAYER ME2 ;
 ANTENNADIFFAREA                          2.912 LAYER ME3 ;
 ANTENNADIFFAREA                          2.912 LAYER ME4 ;
END DO35
PIN DO34
  DIRECTION OUTPUT ;
 PORT
  LAYER ME4 ;
  RECT 231.080 220.480 231.400 221.080 ;
  LAYER ME3 ;
  RECT 231.080 220.480 231.400 221.080 ;
  LAYER ME2 ;
  RECT 231.080 220.480 231.400 221.080 ;
  LAYER ME1 ;
  RECT 231.080 220.480 231.400 221.080 ;
 END
 ANTENNAPARTIALMETALAREA                  0.802 LAYER ME2 ;
 ANTENNADIFFAREA                          2.912 LAYER ME2 ;
 ANTENNADIFFAREA                          2.912 LAYER ME3 ;
 ANTENNADIFFAREA                          2.912 LAYER ME4 ;
END DO34
PIN DO33
  DIRECTION OUTPUT ;
 PORT
  LAYER ME4 ;
  RECT 224.480 220.480 224.800 221.080 ;
  LAYER ME3 ;
  RECT 224.480 220.480 224.800 221.080 ;
  LAYER ME2 ;
  RECT 224.480 220.480 224.800 221.080 ;
  LAYER ME1 ;
  RECT 224.480 220.480 224.800 221.080 ;
 END
 ANTENNAPARTIALMETALAREA                  0.802 LAYER ME2 ;
 ANTENNADIFFAREA                          2.912 LAYER ME2 ;
 ANTENNADIFFAREA                          2.912 LAYER ME3 ;
 ANTENNADIFFAREA                          2.912 LAYER ME4 ;
END DO33
PIN DO32
  DIRECTION OUTPUT ;
 PORT
  LAYER ME4 ;
  RECT 217.880 220.480 218.200 221.080 ;
  LAYER ME3 ;
  RECT 217.880 220.480 218.200 221.080 ;
  LAYER ME2 ;
  RECT 217.880 220.480 218.200 221.080 ;
  LAYER ME1 ;
  RECT 217.880 220.480 218.200 221.080 ;
 END
 ANTENNAPARTIALMETALAREA                  0.802 LAYER ME2 ;
 ANTENNADIFFAREA                          2.912 LAYER ME2 ;
 ANTENNADIFFAREA                          2.912 LAYER ME3 ;
 ANTENNADIFFAREA                          2.912 LAYER ME4 ;
END DO32
PIN DO31
  DIRECTION OUTPUT ;
 PORT
  LAYER ME4 ;
  RECT 211.280 220.480 211.600 221.080 ;
  LAYER ME3 ;
  RECT 211.280 220.480 211.600 221.080 ;
  LAYER ME2 ;
  RECT 211.280 220.480 211.600 221.080 ;
  LAYER ME1 ;
  RECT 211.280 220.480 211.600 221.080 ;
 END
 ANTENNAPARTIALMETALAREA                  0.802 LAYER ME2 ;
 ANTENNADIFFAREA                          2.912 LAYER ME2 ;
 ANTENNADIFFAREA                          2.912 LAYER ME3 ;
 ANTENNADIFFAREA                          2.912 LAYER ME4 ;
END DO31
PIN DO30
  DIRECTION OUTPUT ;
 PORT
  LAYER ME4 ;
  RECT 204.680 220.480 205.000 221.080 ;
  LAYER ME3 ;
  RECT 204.680 220.480 205.000 221.080 ;
  LAYER ME2 ;
  RECT 204.680 220.480 205.000 221.080 ;
  LAYER ME1 ;
  RECT 204.680 220.480 205.000 221.080 ;
 END
 ANTENNAPARTIALMETALAREA                  0.802 LAYER ME2 ;
 ANTENNADIFFAREA                          2.912 LAYER ME2 ;
 ANTENNADIFFAREA                          2.912 LAYER ME3 ;
 ANTENNADIFFAREA                          2.912 LAYER ME4 ;
END DO30
PIN DO29
  DIRECTION OUTPUT ;
 PORT
  LAYER ME4 ;
  RECT 198.080 220.480 198.400 221.080 ;
  LAYER ME3 ;
  RECT 198.080 220.480 198.400 221.080 ;
  LAYER ME2 ;
  RECT 198.080 220.480 198.400 221.080 ;
  LAYER ME1 ;
  RECT 198.080 220.480 198.400 221.080 ;
 END
 ANTENNAPARTIALMETALAREA                  0.802 LAYER ME2 ;
 ANTENNADIFFAREA                          2.912 LAYER ME2 ;
 ANTENNADIFFAREA                          2.912 LAYER ME3 ;
 ANTENNADIFFAREA                          2.912 LAYER ME4 ;
END DO29
PIN DO28
  DIRECTION OUTPUT ;
 PORT
  LAYER ME4 ;
  RECT 191.480 220.480 191.800 221.080 ;
  LAYER ME3 ;
  RECT 191.480 220.480 191.800 221.080 ;
  LAYER ME2 ;
  RECT 191.480 220.480 191.800 221.080 ;
  LAYER ME1 ;
  RECT 191.480 220.480 191.800 221.080 ;
 END
 ANTENNAPARTIALMETALAREA                  0.802 LAYER ME2 ;
 ANTENNADIFFAREA                          2.912 LAYER ME2 ;
 ANTENNADIFFAREA                          2.912 LAYER ME3 ;
 ANTENNADIFFAREA                          2.912 LAYER ME4 ;
END DO28
PIN DO27
  DIRECTION OUTPUT ;
 PORT
  LAYER ME4 ;
  RECT 184.880 220.480 185.200 221.080 ;
  LAYER ME3 ;
  RECT 184.880 220.480 185.200 221.080 ;
  LAYER ME2 ;
  RECT 184.880 220.480 185.200 221.080 ;
  LAYER ME1 ;
  RECT 184.880 220.480 185.200 221.080 ;
 END
 ANTENNAPARTIALMETALAREA                  0.802 LAYER ME2 ;
 ANTENNADIFFAREA                          2.912 LAYER ME2 ;
 ANTENNADIFFAREA                          2.912 LAYER ME3 ;
 ANTENNADIFFAREA                          2.912 LAYER ME4 ;
END DO27
PIN DO26
  DIRECTION OUTPUT ;
 PORT
  LAYER ME4 ;
  RECT 178.280 220.480 178.600 221.080 ;
  LAYER ME3 ;
  RECT 178.280 220.480 178.600 221.080 ;
  LAYER ME2 ;
  RECT 178.280 220.480 178.600 221.080 ;
  LAYER ME1 ;
  RECT 178.280 220.480 178.600 221.080 ;
 END
 ANTENNAPARTIALMETALAREA                  0.802 LAYER ME2 ;
 ANTENNADIFFAREA                          2.912 LAYER ME2 ;
 ANTENNADIFFAREA                          2.912 LAYER ME3 ;
 ANTENNADIFFAREA                          2.912 LAYER ME4 ;
END DO26
PIN DO25
  DIRECTION OUTPUT ;
 PORT
  LAYER ME4 ;
  RECT 171.680 220.480 172.000 221.080 ;
  LAYER ME3 ;
  RECT 171.680 220.480 172.000 221.080 ;
  LAYER ME2 ;
  RECT 171.680 220.480 172.000 221.080 ;
  LAYER ME1 ;
  RECT 171.680 220.480 172.000 221.080 ;
 END
 ANTENNAPARTIALMETALAREA                  0.802 LAYER ME2 ;
 ANTENNADIFFAREA                          2.912 LAYER ME2 ;
 ANTENNADIFFAREA                          2.912 LAYER ME3 ;
 ANTENNADIFFAREA                          2.912 LAYER ME4 ;
END DO25
PIN DO24
  DIRECTION OUTPUT ;
 PORT
  LAYER ME4 ;
  RECT 165.080 220.480 165.400 221.080 ;
  LAYER ME3 ;
  RECT 165.080 220.480 165.400 221.080 ;
  LAYER ME2 ;
  RECT 165.080 220.480 165.400 221.080 ;
  LAYER ME1 ;
  RECT 165.080 220.480 165.400 221.080 ;
 END
 ANTENNAPARTIALMETALAREA                  0.802 LAYER ME2 ;
 ANTENNADIFFAREA                          2.912 LAYER ME2 ;
 ANTENNADIFFAREA                          2.912 LAYER ME3 ;
 ANTENNADIFFAREA                          2.912 LAYER ME4 ;
END DO24
PIN DO23
  DIRECTION OUTPUT ;
 PORT
  LAYER ME4 ;
  RECT 158.480 220.480 158.800 221.080 ;
  LAYER ME3 ;
  RECT 158.480 220.480 158.800 221.080 ;
  LAYER ME2 ;
  RECT 158.480 220.480 158.800 221.080 ;
  LAYER ME1 ;
  RECT 158.480 220.480 158.800 221.080 ;
 END
 ANTENNAPARTIALMETALAREA                  0.802 LAYER ME2 ;
 ANTENNADIFFAREA                          2.912 LAYER ME2 ;
 ANTENNADIFFAREA                          2.912 LAYER ME3 ;
 ANTENNADIFFAREA                          2.912 LAYER ME4 ;
END DO23
PIN DO22
  DIRECTION OUTPUT ;
 PORT
  LAYER ME4 ;
  RECT 151.880 220.480 152.200 221.080 ;
  LAYER ME3 ;
  RECT 151.880 220.480 152.200 221.080 ;
  LAYER ME2 ;
  RECT 151.880 220.480 152.200 221.080 ;
  LAYER ME1 ;
  RECT 151.880 220.480 152.200 221.080 ;
 END
 ANTENNAPARTIALMETALAREA                  0.802 LAYER ME2 ;
 ANTENNADIFFAREA                          2.912 LAYER ME2 ;
 ANTENNADIFFAREA                          2.912 LAYER ME3 ;
 ANTENNADIFFAREA                          2.912 LAYER ME4 ;
END DO22
PIN DO21
  DIRECTION OUTPUT ;
 PORT
  LAYER ME4 ;
  RECT 145.280 220.480 145.600 221.080 ;
  LAYER ME3 ;
  RECT 145.280 220.480 145.600 221.080 ;
  LAYER ME2 ;
  RECT 145.280 220.480 145.600 221.080 ;
  LAYER ME1 ;
  RECT 145.280 220.480 145.600 221.080 ;
 END
 ANTENNAPARTIALMETALAREA                  0.802 LAYER ME2 ;
 ANTENNADIFFAREA                          2.912 LAYER ME2 ;
 ANTENNADIFFAREA                          2.912 LAYER ME3 ;
 ANTENNADIFFAREA                          2.912 LAYER ME4 ;
END DO21
PIN DO20
  DIRECTION OUTPUT ;
 PORT
  LAYER ME4 ;
  RECT 138.680 220.480 139.000 221.080 ;
  LAYER ME3 ;
  RECT 138.680 220.480 139.000 221.080 ;
  LAYER ME2 ;
  RECT 138.680 220.480 139.000 221.080 ;
  LAYER ME1 ;
  RECT 138.680 220.480 139.000 221.080 ;
 END
 ANTENNAPARTIALMETALAREA                  0.802 LAYER ME2 ;
 ANTENNADIFFAREA                          2.912 LAYER ME2 ;
 ANTENNADIFFAREA                          2.912 LAYER ME3 ;
 ANTENNADIFFAREA                          2.912 LAYER ME4 ;
END DO20
PIN DO19
  DIRECTION OUTPUT ;
 PORT
  LAYER ME4 ;
  RECT 132.080 220.480 132.400 221.080 ;
  LAYER ME3 ;
  RECT 132.080 220.480 132.400 221.080 ;
  LAYER ME2 ;
  RECT 132.080 220.480 132.400 221.080 ;
  LAYER ME1 ;
  RECT 132.080 220.480 132.400 221.080 ;
 END
 ANTENNAPARTIALMETALAREA                  0.802 LAYER ME2 ;
 ANTENNADIFFAREA                          2.912 LAYER ME2 ;
 ANTENNADIFFAREA                          2.912 LAYER ME3 ;
 ANTENNADIFFAREA                          2.912 LAYER ME4 ;
END DO19
PIN DO18
  DIRECTION OUTPUT ;
 PORT
  LAYER ME4 ;
  RECT 125.480 220.480 125.800 221.080 ;
  LAYER ME3 ;
  RECT 125.480 220.480 125.800 221.080 ;
  LAYER ME2 ;
  RECT 125.480 220.480 125.800 221.080 ;
  LAYER ME1 ;
  RECT 125.480 220.480 125.800 221.080 ;
 END
 ANTENNAPARTIALMETALAREA                  0.802 LAYER ME2 ;
 ANTENNADIFFAREA                          2.912 LAYER ME2 ;
 ANTENNADIFFAREA                          2.912 LAYER ME3 ;
 ANTENNADIFFAREA                          2.912 LAYER ME4 ;
END DO18
PIN DO17
  DIRECTION OUTPUT ;
 PORT
  LAYER ME4 ;
  RECT 118.880 220.480 119.200 221.080 ;
  LAYER ME3 ;
  RECT 118.880 220.480 119.200 221.080 ;
  LAYER ME2 ;
  RECT 118.880 220.480 119.200 221.080 ;
  LAYER ME1 ;
  RECT 118.880 220.480 119.200 221.080 ;
 END
 ANTENNAPARTIALMETALAREA                  0.802 LAYER ME2 ;
 ANTENNADIFFAREA                          2.912 LAYER ME2 ;
 ANTENNADIFFAREA                          2.912 LAYER ME3 ;
 ANTENNADIFFAREA                          2.912 LAYER ME4 ;
END DO17
PIN DO16
  DIRECTION OUTPUT ;
 PORT
  LAYER ME4 ;
  RECT 112.280 220.480 112.600 221.080 ;
  LAYER ME3 ;
  RECT 112.280 220.480 112.600 221.080 ;
  LAYER ME2 ;
  RECT 112.280 220.480 112.600 221.080 ;
  LAYER ME1 ;
  RECT 112.280 220.480 112.600 221.080 ;
 END
 ANTENNAPARTIALMETALAREA                  0.802 LAYER ME2 ;
 ANTENNADIFFAREA                          2.912 LAYER ME2 ;
 ANTENNADIFFAREA                          2.912 LAYER ME3 ;
 ANTENNADIFFAREA                          2.912 LAYER ME4 ;
END DO16
PIN DO15
  DIRECTION OUTPUT ;
 PORT
  LAYER ME4 ;
  RECT 105.680 220.480 106.000 221.080 ;
  LAYER ME3 ;
  RECT 105.680 220.480 106.000 221.080 ;
  LAYER ME2 ;
  RECT 105.680 220.480 106.000 221.080 ;
  LAYER ME1 ;
  RECT 105.680 220.480 106.000 221.080 ;
 END
 ANTENNAPARTIALMETALAREA                  0.802 LAYER ME2 ;
 ANTENNADIFFAREA                          2.912 LAYER ME2 ;
 ANTENNADIFFAREA                          2.912 LAYER ME3 ;
 ANTENNADIFFAREA                          2.912 LAYER ME4 ;
END DO15
PIN DO14
  DIRECTION OUTPUT ;
 PORT
  LAYER ME4 ;
  RECT 99.080 220.480 99.400 221.080 ;
  LAYER ME3 ;
  RECT 99.080 220.480 99.400 221.080 ;
  LAYER ME2 ;
  RECT 99.080 220.480 99.400 221.080 ;
  LAYER ME1 ;
  RECT 99.080 220.480 99.400 221.080 ;
 END
 ANTENNAPARTIALMETALAREA                  0.802 LAYER ME2 ;
 ANTENNADIFFAREA                          2.912 LAYER ME2 ;
 ANTENNADIFFAREA                          2.912 LAYER ME3 ;
 ANTENNADIFFAREA                          2.912 LAYER ME4 ;
END DO14
PIN DO13
  DIRECTION OUTPUT ;
 PORT
  LAYER ME4 ;
  RECT 92.480 220.480 92.800 221.080 ;
  LAYER ME3 ;
  RECT 92.480 220.480 92.800 221.080 ;
  LAYER ME2 ;
  RECT 92.480 220.480 92.800 221.080 ;
  LAYER ME1 ;
  RECT 92.480 220.480 92.800 221.080 ;
 END
 ANTENNAPARTIALMETALAREA                  0.802 LAYER ME2 ;
 ANTENNADIFFAREA                          2.912 LAYER ME2 ;
 ANTENNADIFFAREA                          2.912 LAYER ME3 ;
 ANTENNADIFFAREA                          2.912 LAYER ME4 ;
END DO13
PIN DO12
  DIRECTION OUTPUT ;
 PORT
  LAYER ME4 ;
  RECT 85.880 220.480 86.200 221.080 ;
  LAYER ME3 ;
  RECT 85.880 220.480 86.200 221.080 ;
  LAYER ME2 ;
  RECT 85.880 220.480 86.200 221.080 ;
  LAYER ME1 ;
  RECT 85.880 220.480 86.200 221.080 ;
 END
 ANTENNAPARTIALMETALAREA                  0.802 LAYER ME2 ;
 ANTENNADIFFAREA                          2.912 LAYER ME2 ;
 ANTENNADIFFAREA                          2.912 LAYER ME3 ;
 ANTENNADIFFAREA                          2.912 LAYER ME4 ;
END DO12
PIN DO11
  DIRECTION OUTPUT ;
 PORT
  LAYER ME4 ;
  RECT 79.280 220.480 79.600 221.080 ;
  LAYER ME3 ;
  RECT 79.280 220.480 79.600 221.080 ;
  LAYER ME2 ;
  RECT 79.280 220.480 79.600 221.080 ;
  LAYER ME1 ;
  RECT 79.280 220.480 79.600 221.080 ;
 END
 ANTENNAPARTIALMETALAREA                  0.802 LAYER ME2 ;
 ANTENNADIFFAREA                          2.912 LAYER ME2 ;
 ANTENNADIFFAREA                          2.912 LAYER ME3 ;
 ANTENNADIFFAREA                          2.912 LAYER ME4 ;
END DO11
PIN DO10
  DIRECTION OUTPUT ;
 PORT
  LAYER ME4 ;
  RECT 72.680 220.480 73.000 221.080 ;
  LAYER ME3 ;
  RECT 72.680 220.480 73.000 221.080 ;
  LAYER ME2 ;
  RECT 72.680 220.480 73.000 221.080 ;
  LAYER ME1 ;
  RECT 72.680 220.480 73.000 221.080 ;
 END
 ANTENNAPARTIALMETALAREA                  0.802 LAYER ME2 ;
 ANTENNADIFFAREA                          2.912 LAYER ME2 ;
 ANTENNADIFFAREA                          2.912 LAYER ME3 ;
 ANTENNADIFFAREA                          2.912 LAYER ME4 ;
END DO10
PIN DO9
  DIRECTION OUTPUT ;
 PORT
  LAYER ME4 ;
  RECT 66.080 220.480 66.400 221.080 ;
  LAYER ME3 ;
  RECT 66.080 220.480 66.400 221.080 ;
  LAYER ME2 ;
  RECT 66.080 220.480 66.400 221.080 ;
  LAYER ME1 ;
  RECT 66.080 220.480 66.400 221.080 ;
 END
 ANTENNAPARTIALMETALAREA                  0.802 LAYER ME2 ;
 ANTENNADIFFAREA                          2.912 LAYER ME2 ;
 ANTENNADIFFAREA                          2.912 LAYER ME3 ;
 ANTENNADIFFAREA                          2.912 LAYER ME4 ;
END DO9
PIN DO8
  DIRECTION OUTPUT ;
 PORT
  LAYER ME4 ;
  RECT 59.480 220.480 59.800 221.080 ;
  LAYER ME3 ;
  RECT 59.480 220.480 59.800 221.080 ;
  LAYER ME2 ;
  RECT 59.480 220.480 59.800 221.080 ;
  LAYER ME1 ;
  RECT 59.480 220.480 59.800 221.080 ;
 END
 ANTENNAPARTIALMETALAREA                  0.802 LAYER ME2 ;
 ANTENNADIFFAREA                          2.912 LAYER ME2 ;
 ANTENNADIFFAREA                          2.912 LAYER ME3 ;
 ANTENNADIFFAREA                          2.912 LAYER ME4 ;
END DO8
PIN DO7
  DIRECTION OUTPUT ;
 PORT
  LAYER ME4 ;
  RECT 52.880 220.480 53.200 221.080 ;
  LAYER ME3 ;
  RECT 52.880 220.480 53.200 221.080 ;
  LAYER ME2 ;
  RECT 52.880 220.480 53.200 221.080 ;
  LAYER ME1 ;
  RECT 52.880 220.480 53.200 221.080 ;
 END
 ANTENNAPARTIALMETALAREA                  0.802 LAYER ME2 ;
 ANTENNADIFFAREA                          2.912 LAYER ME2 ;
 ANTENNADIFFAREA                          2.912 LAYER ME3 ;
 ANTENNADIFFAREA                          2.912 LAYER ME4 ;
END DO7
PIN DO6
  DIRECTION OUTPUT ;
 PORT
  LAYER ME4 ;
  RECT 46.280 220.480 46.600 221.080 ;
  LAYER ME3 ;
  RECT 46.280 220.480 46.600 221.080 ;
  LAYER ME2 ;
  RECT 46.280 220.480 46.600 221.080 ;
  LAYER ME1 ;
  RECT 46.280 220.480 46.600 221.080 ;
 END
 ANTENNAPARTIALMETALAREA                  0.802 LAYER ME2 ;
 ANTENNADIFFAREA                          2.912 LAYER ME2 ;
 ANTENNADIFFAREA                          2.912 LAYER ME3 ;
 ANTENNADIFFAREA                          2.912 LAYER ME4 ;
END DO6
PIN DO5
  DIRECTION OUTPUT ;
 PORT
  LAYER ME4 ;
  RECT 39.680 220.480 40.000 221.080 ;
  LAYER ME3 ;
  RECT 39.680 220.480 40.000 221.080 ;
  LAYER ME2 ;
  RECT 39.680 220.480 40.000 221.080 ;
  LAYER ME1 ;
  RECT 39.680 220.480 40.000 221.080 ;
 END
 ANTENNAPARTIALMETALAREA                  0.802 LAYER ME2 ;
 ANTENNADIFFAREA                          2.912 LAYER ME2 ;
 ANTENNADIFFAREA                          2.912 LAYER ME3 ;
 ANTENNADIFFAREA                          2.912 LAYER ME4 ;
END DO5
PIN DO4
  DIRECTION OUTPUT ;
 PORT
  LAYER ME4 ;
  RECT 33.080 220.480 33.400 221.080 ;
  LAYER ME3 ;
  RECT 33.080 220.480 33.400 221.080 ;
  LAYER ME2 ;
  RECT 33.080 220.480 33.400 221.080 ;
  LAYER ME1 ;
  RECT 33.080 220.480 33.400 221.080 ;
 END
 ANTENNAPARTIALMETALAREA                  0.802 LAYER ME2 ;
 ANTENNADIFFAREA                          2.912 LAYER ME2 ;
 ANTENNADIFFAREA                          2.912 LAYER ME3 ;
 ANTENNADIFFAREA                          2.912 LAYER ME4 ;
END DO4
PIN DO3
  DIRECTION OUTPUT ;
 PORT
  LAYER ME4 ;
  RECT 26.480 220.480 26.800 221.080 ;
  LAYER ME3 ;
  RECT 26.480 220.480 26.800 221.080 ;
  LAYER ME2 ;
  RECT 26.480 220.480 26.800 221.080 ;
  LAYER ME1 ;
  RECT 26.480 220.480 26.800 221.080 ;
 END
 ANTENNAPARTIALMETALAREA                  0.802 LAYER ME2 ;
 ANTENNADIFFAREA                          2.912 LAYER ME2 ;
 ANTENNADIFFAREA                          2.912 LAYER ME3 ;
 ANTENNADIFFAREA                          2.912 LAYER ME4 ;
END DO3
PIN DO2
  DIRECTION OUTPUT ;
 PORT
  LAYER ME4 ;
  RECT 19.880 220.480 20.200 221.080 ;
  LAYER ME3 ;
  RECT 19.880 220.480 20.200 221.080 ;
  LAYER ME2 ;
  RECT 19.880 220.480 20.200 221.080 ;
  LAYER ME1 ;
  RECT 19.880 220.480 20.200 221.080 ;
 END
 ANTENNAPARTIALMETALAREA                  0.802 LAYER ME2 ;
 ANTENNADIFFAREA                          2.912 LAYER ME2 ;
 ANTENNADIFFAREA                          2.912 LAYER ME3 ;
 ANTENNADIFFAREA                          2.912 LAYER ME4 ;
END DO2
PIN DO1
  DIRECTION OUTPUT ;
 PORT
  LAYER ME4 ;
  RECT 13.280 220.480 13.600 221.080 ;
  LAYER ME3 ;
  RECT 13.280 220.480 13.600 221.080 ;
  LAYER ME2 ;
  RECT 13.280 220.480 13.600 221.080 ;
  LAYER ME1 ;
  RECT 13.280 220.480 13.600 221.080 ;
 END
 ANTENNAPARTIALMETALAREA                  0.802 LAYER ME2 ;
 ANTENNADIFFAREA                          2.912 LAYER ME2 ;
 ANTENNADIFFAREA                          2.912 LAYER ME3 ;
 ANTENNADIFFAREA                          2.912 LAYER ME4 ;
END DO1
PIN DO0
  DIRECTION OUTPUT ;
 PORT
  LAYER ME4 ;
  RECT 6.680 220.480 7.000 221.080 ;
  LAYER ME3 ;
  RECT 6.680 220.480 7.000 221.080 ;
  LAYER ME2 ;
  RECT 6.680 220.480 7.000 221.080 ;
  LAYER ME1 ;
  RECT 6.680 220.480 7.000 221.080 ;
 END
 ANTENNAPARTIALMETALAREA                  0.802 LAYER ME2 ;
 ANTENNADIFFAREA                          2.912 LAYER ME2 ;
 ANTENNADIFFAREA                          2.912 LAYER ME3 ;
 ANTENNADIFFAREA                          2.912 LAYER ME4 ;
END DO0
PIN DO71
  DIRECTION OUTPUT ;
 PORT
  LAYER ME4 ;
  RECT 534.890 220.480 535.210 221.080 ;
  LAYER ME3 ;
  RECT 534.890 220.480 535.210 221.080 ;
  LAYER ME2 ;
  RECT 534.890 220.480 535.210 221.080 ;
  LAYER ME1 ;
  RECT 534.890 220.480 535.210 221.080 ;
 END
 ANTENNAPARTIALMETALAREA                  0.802 LAYER ME2 ;
 ANTENNADIFFAREA                          2.912 LAYER ME2 ;
 ANTENNADIFFAREA                          2.912 LAYER ME3 ;
 ANTENNADIFFAREA                          2.912 LAYER ME4 ;
END DO71
PIN DO70
  DIRECTION OUTPUT ;
 PORT
  LAYER ME4 ;
  RECT 528.290 220.480 528.610 221.080 ;
  LAYER ME3 ;
  RECT 528.290 220.480 528.610 221.080 ;
  LAYER ME2 ;
  RECT 528.290 220.480 528.610 221.080 ;
  LAYER ME1 ;
  RECT 528.290 220.480 528.610 221.080 ;
 END
 ANTENNAPARTIALMETALAREA                  0.802 LAYER ME2 ;
 ANTENNADIFFAREA                          2.912 LAYER ME2 ;
 ANTENNADIFFAREA                          2.912 LAYER ME3 ;
 ANTENNADIFFAREA                          2.912 LAYER ME4 ;
END DO70
PIN DO69
  DIRECTION OUTPUT ;
 PORT
  LAYER ME4 ;
  RECT 521.690 220.480 522.010 221.080 ;
  LAYER ME3 ;
  RECT 521.690 220.480 522.010 221.080 ;
  LAYER ME2 ;
  RECT 521.690 220.480 522.010 221.080 ;
  LAYER ME1 ;
  RECT 521.690 220.480 522.010 221.080 ;
 END
 ANTENNAPARTIALMETALAREA                  0.802 LAYER ME2 ;
 ANTENNADIFFAREA                          2.912 LAYER ME2 ;
 ANTENNADIFFAREA                          2.912 LAYER ME3 ;
 ANTENNADIFFAREA                          2.912 LAYER ME4 ;
END DO69
PIN DO68
  DIRECTION OUTPUT ;
 PORT
  LAYER ME4 ;
  RECT 515.090 220.480 515.410 221.080 ;
  LAYER ME3 ;
  RECT 515.090 220.480 515.410 221.080 ;
  LAYER ME2 ;
  RECT 515.090 220.480 515.410 221.080 ;
  LAYER ME1 ;
  RECT 515.090 220.480 515.410 221.080 ;
 END
 ANTENNAPARTIALMETALAREA                  0.802 LAYER ME2 ;
 ANTENNADIFFAREA                          2.912 LAYER ME2 ;
 ANTENNADIFFAREA                          2.912 LAYER ME3 ;
 ANTENNADIFFAREA                          2.912 LAYER ME4 ;
END DO68
PIN DO67
  DIRECTION OUTPUT ;
 PORT
  LAYER ME4 ;
  RECT 508.490 220.480 508.810 221.080 ;
  LAYER ME3 ;
  RECT 508.490 220.480 508.810 221.080 ;
  LAYER ME2 ;
  RECT 508.490 220.480 508.810 221.080 ;
  LAYER ME1 ;
  RECT 508.490 220.480 508.810 221.080 ;
 END
 ANTENNAPARTIALMETALAREA                  0.802 LAYER ME2 ;
 ANTENNADIFFAREA                          2.912 LAYER ME2 ;
 ANTENNADIFFAREA                          2.912 LAYER ME3 ;
 ANTENNADIFFAREA                          2.912 LAYER ME4 ;
END DO67
PIN DO66
  DIRECTION OUTPUT ;
 PORT
  LAYER ME4 ;
  RECT 501.890 220.480 502.210 221.080 ;
  LAYER ME3 ;
  RECT 501.890 220.480 502.210 221.080 ;
  LAYER ME2 ;
  RECT 501.890 220.480 502.210 221.080 ;
  LAYER ME1 ;
  RECT 501.890 220.480 502.210 221.080 ;
 END
 ANTENNAPARTIALMETALAREA                  0.802 LAYER ME2 ;
 ANTENNADIFFAREA                          2.912 LAYER ME2 ;
 ANTENNADIFFAREA                          2.912 LAYER ME3 ;
 ANTENNADIFFAREA                          2.912 LAYER ME4 ;
END DO66
PIN DO65
  DIRECTION OUTPUT ;
 PORT
  LAYER ME4 ;
  RECT 495.290 220.480 495.610 221.080 ;
  LAYER ME3 ;
  RECT 495.290 220.480 495.610 221.080 ;
  LAYER ME2 ;
  RECT 495.290 220.480 495.610 221.080 ;
  LAYER ME1 ;
  RECT 495.290 220.480 495.610 221.080 ;
 END
 ANTENNAPARTIALMETALAREA                  0.802 LAYER ME2 ;
 ANTENNADIFFAREA                          2.912 LAYER ME2 ;
 ANTENNADIFFAREA                          2.912 LAYER ME3 ;
 ANTENNADIFFAREA                          2.912 LAYER ME4 ;
END DO65
PIN DO64
  DIRECTION OUTPUT ;
 PORT
  LAYER ME4 ;
  RECT 488.690 220.480 489.010 221.080 ;
  LAYER ME3 ;
  RECT 488.690 220.480 489.010 221.080 ;
  LAYER ME2 ;
  RECT 488.690 220.480 489.010 221.080 ;
  LAYER ME1 ;
  RECT 488.690 220.480 489.010 221.080 ;
 END
 ANTENNAPARTIALMETALAREA                  0.802 LAYER ME2 ;
 ANTENNADIFFAREA                          2.912 LAYER ME2 ;
 ANTENNADIFFAREA                          2.912 LAYER ME3 ;
 ANTENNADIFFAREA                          2.912 LAYER ME4 ;
END DO64
PIN DO63
  DIRECTION OUTPUT ;
 PORT
  LAYER ME4 ;
  RECT 482.090 220.480 482.410 221.080 ;
  LAYER ME3 ;
  RECT 482.090 220.480 482.410 221.080 ;
  LAYER ME2 ;
  RECT 482.090 220.480 482.410 221.080 ;
  LAYER ME1 ;
  RECT 482.090 220.480 482.410 221.080 ;
 END
 ANTENNAPARTIALMETALAREA                  0.802 LAYER ME2 ;
 ANTENNADIFFAREA                          2.912 LAYER ME2 ;
 ANTENNADIFFAREA                          2.912 LAYER ME3 ;
 ANTENNADIFFAREA                          2.912 LAYER ME4 ;
END DO63
PIN DO62
  DIRECTION OUTPUT ;
 PORT
  LAYER ME4 ;
  RECT 475.490 220.480 475.810 221.080 ;
  LAYER ME3 ;
  RECT 475.490 220.480 475.810 221.080 ;
  LAYER ME2 ;
  RECT 475.490 220.480 475.810 221.080 ;
  LAYER ME1 ;
  RECT 475.490 220.480 475.810 221.080 ;
 END
 ANTENNAPARTIALMETALAREA                  0.802 LAYER ME2 ;
 ANTENNADIFFAREA                          2.912 LAYER ME2 ;
 ANTENNADIFFAREA                          2.912 LAYER ME3 ;
 ANTENNADIFFAREA                          2.912 LAYER ME4 ;
END DO62
PIN DO61
  DIRECTION OUTPUT ;
 PORT
  LAYER ME4 ;
  RECT 468.890 220.480 469.210 221.080 ;
  LAYER ME3 ;
  RECT 468.890 220.480 469.210 221.080 ;
  LAYER ME2 ;
  RECT 468.890 220.480 469.210 221.080 ;
  LAYER ME1 ;
  RECT 468.890 220.480 469.210 221.080 ;
 END
 ANTENNAPARTIALMETALAREA                  0.802 LAYER ME2 ;
 ANTENNADIFFAREA                          2.912 LAYER ME2 ;
 ANTENNADIFFAREA                          2.912 LAYER ME3 ;
 ANTENNADIFFAREA                          2.912 LAYER ME4 ;
END DO61
PIN DO60
  DIRECTION OUTPUT ;
 PORT
  LAYER ME4 ;
  RECT 462.290 220.480 462.610 221.080 ;
  LAYER ME3 ;
  RECT 462.290 220.480 462.610 221.080 ;
  LAYER ME2 ;
  RECT 462.290 220.480 462.610 221.080 ;
  LAYER ME1 ;
  RECT 462.290 220.480 462.610 221.080 ;
 END
 ANTENNAPARTIALMETALAREA                  0.802 LAYER ME2 ;
 ANTENNADIFFAREA                          2.912 LAYER ME2 ;
 ANTENNADIFFAREA                          2.912 LAYER ME3 ;
 ANTENNADIFFAREA                          2.912 LAYER ME4 ;
END DO60
PIN DO59
  DIRECTION OUTPUT ;
 PORT
  LAYER ME4 ;
  RECT 455.690 220.480 456.010 221.080 ;
  LAYER ME3 ;
  RECT 455.690 220.480 456.010 221.080 ;
  LAYER ME2 ;
  RECT 455.690 220.480 456.010 221.080 ;
  LAYER ME1 ;
  RECT 455.690 220.480 456.010 221.080 ;
 END
 ANTENNAPARTIALMETALAREA                  0.802 LAYER ME2 ;
 ANTENNADIFFAREA                          2.912 LAYER ME2 ;
 ANTENNADIFFAREA                          2.912 LAYER ME3 ;
 ANTENNADIFFAREA                          2.912 LAYER ME4 ;
END DO59
PIN DO58
  DIRECTION OUTPUT ;
 PORT
  LAYER ME4 ;
  RECT 449.090 220.480 449.410 221.080 ;
  LAYER ME3 ;
  RECT 449.090 220.480 449.410 221.080 ;
  LAYER ME2 ;
  RECT 449.090 220.480 449.410 221.080 ;
  LAYER ME1 ;
  RECT 449.090 220.480 449.410 221.080 ;
 END
 ANTENNAPARTIALMETALAREA                  0.802 LAYER ME2 ;
 ANTENNADIFFAREA                          2.912 LAYER ME2 ;
 ANTENNADIFFAREA                          2.912 LAYER ME3 ;
 ANTENNADIFFAREA                          2.912 LAYER ME4 ;
END DO58
PIN DO57
  DIRECTION OUTPUT ;
 PORT
  LAYER ME4 ;
  RECT 442.490 220.480 442.810 221.080 ;
  LAYER ME3 ;
  RECT 442.490 220.480 442.810 221.080 ;
  LAYER ME2 ;
  RECT 442.490 220.480 442.810 221.080 ;
  LAYER ME1 ;
  RECT 442.490 220.480 442.810 221.080 ;
 END
 ANTENNAPARTIALMETALAREA                  0.802 LAYER ME2 ;
 ANTENNADIFFAREA                          2.912 LAYER ME2 ;
 ANTENNADIFFAREA                          2.912 LAYER ME3 ;
 ANTENNADIFFAREA                          2.912 LAYER ME4 ;
END DO57
PIN DO56
  DIRECTION OUTPUT ;
 PORT
  LAYER ME4 ;
  RECT 435.890 220.480 436.210 221.080 ;
  LAYER ME3 ;
  RECT 435.890 220.480 436.210 221.080 ;
  LAYER ME2 ;
  RECT 435.890 220.480 436.210 221.080 ;
  LAYER ME1 ;
  RECT 435.890 220.480 436.210 221.080 ;
 END
 ANTENNAPARTIALMETALAREA                  0.802 LAYER ME2 ;
 ANTENNADIFFAREA                          2.912 LAYER ME2 ;
 ANTENNADIFFAREA                          2.912 LAYER ME3 ;
 ANTENNADIFFAREA                          2.912 LAYER ME4 ;
END DO56
PIN DO55
  DIRECTION OUTPUT ;
 PORT
  LAYER ME4 ;
  RECT 429.290 220.480 429.610 221.080 ;
  LAYER ME3 ;
  RECT 429.290 220.480 429.610 221.080 ;
  LAYER ME2 ;
  RECT 429.290 220.480 429.610 221.080 ;
  LAYER ME1 ;
  RECT 429.290 220.480 429.610 221.080 ;
 END
 ANTENNAPARTIALMETALAREA                  0.802 LAYER ME2 ;
 ANTENNADIFFAREA                          2.912 LAYER ME2 ;
 ANTENNADIFFAREA                          2.912 LAYER ME3 ;
 ANTENNADIFFAREA                          2.912 LAYER ME4 ;
END DO55
PIN DO54
  DIRECTION OUTPUT ;
 PORT
  LAYER ME4 ;
  RECT 422.690 220.480 423.010 221.080 ;
  LAYER ME3 ;
  RECT 422.690 220.480 423.010 221.080 ;
  LAYER ME2 ;
  RECT 422.690 220.480 423.010 221.080 ;
  LAYER ME1 ;
  RECT 422.690 220.480 423.010 221.080 ;
 END
 ANTENNAPARTIALMETALAREA                  0.802 LAYER ME2 ;
 ANTENNADIFFAREA                          2.912 LAYER ME2 ;
 ANTENNADIFFAREA                          2.912 LAYER ME3 ;
 ANTENNADIFFAREA                          2.912 LAYER ME4 ;
END DO54
PIN DO53
  DIRECTION OUTPUT ;
 PORT
  LAYER ME4 ;
  RECT 416.090 220.480 416.410 221.080 ;
  LAYER ME3 ;
  RECT 416.090 220.480 416.410 221.080 ;
  LAYER ME2 ;
  RECT 416.090 220.480 416.410 221.080 ;
  LAYER ME1 ;
  RECT 416.090 220.480 416.410 221.080 ;
 END
 ANTENNAPARTIALMETALAREA                  0.802 LAYER ME2 ;
 ANTENNADIFFAREA                          2.912 LAYER ME2 ;
 ANTENNADIFFAREA                          2.912 LAYER ME3 ;
 ANTENNADIFFAREA                          2.912 LAYER ME4 ;
END DO53
PIN DO52
  DIRECTION OUTPUT ;
 PORT
  LAYER ME4 ;
  RECT 409.490 220.480 409.810 221.080 ;
  LAYER ME3 ;
  RECT 409.490 220.480 409.810 221.080 ;
  LAYER ME2 ;
  RECT 409.490 220.480 409.810 221.080 ;
  LAYER ME1 ;
  RECT 409.490 220.480 409.810 221.080 ;
 END
 ANTENNAPARTIALMETALAREA                  0.802 LAYER ME2 ;
 ANTENNADIFFAREA                          2.912 LAYER ME2 ;
 ANTENNADIFFAREA                          2.912 LAYER ME3 ;
 ANTENNADIFFAREA                          2.912 LAYER ME4 ;
END DO52
PIN DO51
  DIRECTION OUTPUT ;
 PORT
  LAYER ME4 ;
  RECT 402.890 220.480 403.210 221.080 ;
  LAYER ME3 ;
  RECT 402.890 220.480 403.210 221.080 ;
  LAYER ME2 ;
  RECT 402.890 220.480 403.210 221.080 ;
  LAYER ME1 ;
  RECT 402.890 220.480 403.210 221.080 ;
 END
 ANTENNAPARTIALMETALAREA                  0.802 LAYER ME2 ;
 ANTENNADIFFAREA                          2.912 LAYER ME2 ;
 ANTENNADIFFAREA                          2.912 LAYER ME3 ;
 ANTENNADIFFAREA                          2.912 LAYER ME4 ;
END DO51
PIN DO50
  DIRECTION OUTPUT ;
 PORT
  LAYER ME4 ;
  RECT 396.290 220.480 396.610 221.080 ;
  LAYER ME3 ;
  RECT 396.290 220.480 396.610 221.080 ;
  LAYER ME2 ;
  RECT 396.290 220.480 396.610 221.080 ;
  LAYER ME1 ;
  RECT 396.290 220.480 396.610 221.080 ;
 END
 ANTENNAPARTIALMETALAREA                  0.802 LAYER ME2 ;
 ANTENNADIFFAREA                          2.912 LAYER ME2 ;
 ANTENNADIFFAREA                          2.912 LAYER ME3 ;
 ANTENNADIFFAREA                          2.912 LAYER ME4 ;
END DO50
PIN DO49
  DIRECTION OUTPUT ;
 PORT
  LAYER ME4 ;
  RECT 389.690 220.480 390.010 221.080 ;
  LAYER ME3 ;
  RECT 389.690 220.480 390.010 221.080 ;
  LAYER ME2 ;
  RECT 389.690 220.480 390.010 221.080 ;
  LAYER ME1 ;
  RECT 389.690 220.480 390.010 221.080 ;
 END
 ANTENNAPARTIALMETALAREA                  0.802 LAYER ME2 ;
 ANTENNADIFFAREA                          2.912 LAYER ME2 ;
 ANTENNADIFFAREA                          2.912 LAYER ME3 ;
 ANTENNADIFFAREA                          2.912 LAYER ME4 ;
END DO49
PIN DO48
  DIRECTION OUTPUT ;
 PORT
  LAYER ME4 ;
  RECT 383.090 220.480 383.410 221.080 ;
  LAYER ME3 ;
  RECT 383.090 220.480 383.410 221.080 ;
  LAYER ME2 ;
  RECT 383.090 220.480 383.410 221.080 ;
  LAYER ME1 ;
  RECT 383.090 220.480 383.410 221.080 ;
 END
 ANTENNAPARTIALMETALAREA                  0.802 LAYER ME2 ;
 ANTENNADIFFAREA                          2.912 LAYER ME2 ;
 ANTENNADIFFAREA                          2.912 LAYER ME3 ;
 ANTENNADIFFAREA                          2.912 LAYER ME4 ;
END DO48
PIN DO47
  DIRECTION OUTPUT ;
 PORT
  LAYER ME4 ;
  RECT 376.490 220.480 376.810 221.080 ;
  LAYER ME3 ;
  RECT 376.490 220.480 376.810 221.080 ;
  LAYER ME2 ;
  RECT 376.490 220.480 376.810 221.080 ;
  LAYER ME1 ;
  RECT 376.490 220.480 376.810 221.080 ;
 END
 ANTENNAPARTIALMETALAREA                  0.802 LAYER ME2 ;
 ANTENNADIFFAREA                          2.912 LAYER ME2 ;
 ANTENNADIFFAREA                          2.912 LAYER ME3 ;
 ANTENNADIFFAREA                          2.912 LAYER ME4 ;
END DO47
PIN DO46
  DIRECTION OUTPUT ;
 PORT
  LAYER ME4 ;
  RECT 369.890 220.480 370.210 221.080 ;
  LAYER ME3 ;
  RECT 369.890 220.480 370.210 221.080 ;
  LAYER ME2 ;
  RECT 369.890 220.480 370.210 221.080 ;
  LAYER ME1 ;
  RECT 369.890 220.480 370.210 221.080 ;
 END
 ANTENNAPARTIALMETALAREA                  0.802 LAYER ME2 ;
 ANTENNADIFFAREA                          2.912 LAYER ME2 ;
 ANTENNADIFFAREA                          2.912 LAYER ME3 ;
 ANTENNADIFFAREA                          2.912 LAYER ME4 ;
END DO46
PIN DO45
  DIRECTION OUTPUT ;
 PORT
  LAYER ME4 ;
  RECT 363.290 220.480 363.610 221.080 ;
  LAYER ME3 ;
  RECT 363.290 220.480 363.610 221.080 ;
  LAYER ME2 ;
  RECT 363.290 220.480 363.610 221.080 ;
  LAYER ME1 ;
  RECT 363.290 220.480 363.610 221.080 ;
 END
 ANTENNAPARTIALMETALAREA                  0.802 LAYER ME2 ;
 ANTENNADIFFAREA                          2.912 LAYER ME2 ;
 ANTENNADIFFAREA                          2.912 LAYER ME3 ;
 ANTENNADIFFAREA                          2.912 LAYER ME4 ;
END DO45
PIN DO44
  DIRECTION OUTPUT ;
 PORT
  LAYER ME4 ;
  RECT 356.690 220.480 357.010 221.080 ;
  LAYER ME3 ;
  RECT 356.690 220.480 357.010 221.080 ;
  LAYER ME2 ;
  RECT 356.690 220.480 357.010 221.080 ;
  LAYER ME1 ;
  RECT 356.690 220.480 357.010 221.080 ;
 END
 ANTENNAPARTIALMETALAREA                  0.802 LAYER ME2 ;
 ANTENNADIFFAREA                          2.912 LAYER ME2 ;
 ANTENNADIFFAREA                          2.912 LAYER ME3 ;
 ANTENNADIFFAREA                          2.912 LAYER ME4 ;
END DO44
PIN DO43
  DIRECTION OUTPUT ;
 PORT
  LAYER ME4 ;
  RECT 350.090 220.480 350.410 221.080 ;
  LAYER ME3 ;
  RECT 350.090 220.480 350.410 221.080 ;
  LAYER ME2 ;
  RECT 350.090 220.480 350.410 221.080 ;
  LAYER ME1 ;
  RECT 350.090 220.480 350.410 221.080 ;
 END
 ANTENNAPARTIALMETALAREA                  0.802 LAYER ME2 ;
 ANTENNADIFFAREA                          2.912 LAYER ME2 ;
 ANTENNADIFFAREA                          2.912 LAYER ME3 ;
 ANTENNADIFFAREA                          2.912 LAYER ME4 ;
END DO43
PIN DO42
  DIRECTION OUTPUT ;
 PORT
  LAYER ME4 ;
  RECT 343.490 220.480 343.810 221.080 ;
  LAYER ME3 ;
  RECT 343.490 220.480 343.810 221.080 ;
  LAYER ME2 ;
  RECT 343.490 220.480 343.810 221.080 ;
  LAYER ME1 ;
  RECT 343.490 220.480 343.810 221.080 ;
 END
 ANTENNAPARTIALMETALAREA                  0.802 LAYER ME2 ;
 ANTENNADIFFAREA                          2.912 LAYER ME2 ;
 ANTENNADIFFAREA                          2.912 LAYER ME3 ;
 ANTENNADIFFAREA                          2.912 LAYER ME4 ;
END DO42
PIN DO41
  DIRECTION OUTPUT ;
 PORT
  LAYER ME4 ;
  RECT 336.890 220.480 337.210 221.080 ;
  LAYER ME3 ;
  RECT 336.890 220.480 337.210 221.080 ;
  LAYER ME2 ;
  RECT 336.890 220.480 337.210 221.080 ;
  LAYER ME1 ;
  RECT 336.890 220.480 337.210 221.080 ;
 END
 ANTENNAPARTIALMETALAREA                  0.802 LAYER ME2 ;
 ANTENNADIFFAREA                          2.912 LAYER ME2 ;
 ANTENNADIFFAREA                          2.912 LAYER ME3 ;
 ANTENNADIFFAREA                          2.912 LAYER ME4 ;
END DO41
PIN DO40
  DIRECTION OUTPUT ;
 PORT
  LAYER ME4 ;
  RECT 330.290 220.480 330.610 221.080 ;
  LAYER ME3 ;
  RECT 330.290 220.480 330.610 221.080 ;
  LAYER ME2 ;
  RECT 330.290 220.480 330.610 221.080 ;
  LAYER ME1 ;
  RECT 330.290 220.480 330.610 221.080 ;
 END
 ANTENNAPARTIALMETALAREA                  0.802 LAYER ME2 ;
 ANTENNADIFFAREA                          2.912 LAYER ME2 ;
 ANTENNADIFFAREA                          2.912 LAYER ME3 ;
 ANTENNADIFFAREA                          2.912 LAYER ME4 ;
END DO40
PIN DO39
  DIRECTION OUTPUT ;
 PORT
  LAYER ME4 ;
  RECT 323.690 220.480 324.010 221.080 ;
  LAYER ME3 ;
  RECT 323.690 220.480 324.010 221.080 ;
  LAYER ME2 ;
  RECT 323.690 220.480 324.010 221.080 ;
  LAYER ME1 ;
  RECT 323.690 220.480 324.010 221.080 ;
 END
 ANTENNAPARTIALMETALAREA                  0.802 LAYER ME2 ;
 ANTENNADIFFAREA                          2.912 LAYER ME2 ;
 ANTENNADIFFAREA                          2.912 LAYER ME3 ;
 ANTENNADIFFAREA                          2.912 LAYER ME4 ;
END DO39
PIN DO38
  DIRECTION OUTPUT ;
 PORT
  LAYER ME4 ;
  RECT 317.090 220.480 317.410 221.080 ;
  LAYER ME3 ;
  RECT 317.090 220.480 317.410 221.080 ;
  LAYER ME2 ;
  RECT 317.090 220.480 317.410 221.080 ;
  LAYER ME1 ;
  RECT 317.090 220.480 317.410 221.080 ;
 END
 ANTENNAPARTIALMETALAREA                  0.802 LAYER ME2 ;
 ANTENNADIFFAREA                          2.912 LAYER ME2 ;
 ANTENNADIFFAREA                          2.912 LAYER ME3 ;
 ANTENNADIFFAREA                          2.912 LAYER ME4 ;
END DO38
PIN DO37
  DIRECTION OUTPUT ;
 PORT
  LAYER ME4 ;
  RECT 310.490 220.480 310.810 221.080 ;
  LAYER ME3 ;
  RECT 310.490 220.480 310.810 221.080 ;
  LAYER ME2 ;
  RECT 310.490 220.480 310.810 221.080 ;
  LAYER ME1 ;
  RECT 310.490 220.480 310.810 221.080 ;
 END
 ANTENNAPARTIALMETALAREA                  0.802 LAYER ME2 ;
 ANTENNADIFFAREA                          2.912 LAYER ME2 ;
 ANTENNADIFFAREA                          2.912 LAYER ME3 ;
 ANTENNADIFFAREA                          2.912 LAYER ME4 ;
END DO37
PIN DO36
  DIRECTION OUTPUT ;
 PORT
  LAYER ME4 ;
  RECT 303.890 220.480 304.210 221.080 ;
  LAYER ME3 ;
  RECT 303.890 220.480 304.210 221.080 ;
  LAYER ME2 ;
  RECT 303.890 220.480 304.210 221.080 ;
  LAYER ME1 ;
  RECT 303.890 220.480 304.210 221.080 ;
 END
 ANTENNAPARTIALMETALAREA                  0.802 LAYER ME2 ;
 ANTENNADIFFAREA                          2.912 LAYER ME2 ;
 ANTENNADIFFAREA                          2.912 LAYER ME3 ;
 ANTENNADIFFAREA                          2.912 LAYER ME4 ;
END DO36
PIN B7
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 244.060 0.000 244.380 0.600 ;
  LAYER ME3 ;
  RECT 244.060 0.000 244.380 0.600 ;
  LAYER ME2 ;
  RECT 244.060 0.000 244.380 0.600 ;
  LAYER ME1 ;
  RECT 244.060 0.000 244.380 0.600 ;
 END
 ANTENNAPARTIALMETALAREA                  0.984 LAYER ME2 ;
 ANTENNAPARTIALMETALAREA                  0.768 LAYER ME3 ;
 ANTENNAGATEAREA                          0.216 LAYER ME2 ;
 ANTENNAGATEAREA                          0.216 LAYER ME3 ;
 ANTENNAGATEAREA                          0.216 LAYER ME4 ;
 ANTENNADIFFAREA                          0.160 LAYER ME2 ;
 ANTENNADIFFAREA                          0.160 LAYER ME3 ;
 ANTENNADIFFAREA                          0.160 LAYER ME4 ;
 ANTENNAMAXAREACAR                        6.983 LAYER ME2 ;
 ANTENNAMAXAREACAR                       11.428 LAYER ME3 ;
 ANTENNAMAXAREACAR                       12.317 LAYER ME4 ;
END B7
PIN B6
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 247.580 0.000 247.900 0.600 ;
  LAYER ME3 ;
  RECT 247.580 0.000 247.900 0.600 ;
  LAYER ME2 ;
  RECT 247.580 0.000 247.900 0.600 ;
  LAYER ME1 ;
  RECT 247.580 0.000 247.900 0.600 ;
 END
 ANTENNAPARTIALMETALAREA                  0.906 LAYER ME2 ;
 ANTENNAGATEAREA                          0.216 LAYER ME2 ;
 ANTENNAGATEAREA                          0.216 LAYER ME3 ;
 ANTENNAGATEAREA                          0.216 LAYER ME4 ;
 ANTENNADIFFAREA                          0.160 LAYER ME2 ;
 ANTENNADIFFAREA                          0.160 LAYER ME3 ;
 ANTENNADIFFAREA                          0.160 LAYER ME4 ;
 ANTENNAMAXAREACAR                        7.863 LAYER ME2 ;
 ANTENNAMAXAREACAR                        8.752 LAYER ME3 ;
 ANTENNAMAXAREACAR                        9.641 LAYER ME4 ;
END B6
PIN B5
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 250.420 0.000 250.740 0.600 ;
  LAYER ME3 ;
  RECT 250.420 0.000 250.740 0.600 ;
  LAYER ME2 ;
  RECT 250.420 0.000 250.740 0.600 ;
  LAYER ME1 ;
  RECT 250.420 0.000 250.740 0.600 ;
 END
 ANTENNAPARTIALMETALAREA                  0.984 LAYER ME2 ;
 ANTENNAPARTIALMETALAREA                  0.768 LAYER ME3 ;
 ANTENNAGATEAREA                          0.216 LAYER ME2 ;
 ANTENNAGATEAREA                          0.216 LAYER ME3 ;
 ANTENNAGATEAREA                          0.216 LAYER ME4 ;
 ANTENNADIFFAREA                          0.160 LAYER ME2 ;
 ANTENNADIFFAREA                          0.160 LAYER ME3 ;
 ANTENNADIFFAREA                          0.160 LAYER ME4 ;
 ANTENNAMAXAREACAR                        6.983 LAYER ME2 ;
 ANTENNAMAXAREACAR                       11.428 LAYER ME3 ;
 ANTENNAMAXAREACAR                       12.317 LAYER ME4 ;
END B5
PIN B4
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 253.940 0.000 254.260 0.600 ;
  LAYER ME3 ;
  RECT 253.940 0.000 254.260 0.600 ;
  LAYER ME2 ;
  RECT 253.940 0.000 254.260 0.600 ;
  LAYER ME1 ;
  RECT 253.940 0.000 254.260 0.600 ;
 END
 ANTENNAPARTIALMETALAREA                  0.906 LAYER ME2 ;
 ANTENNAGATEAREA                          0.216 LAYER ME2 ;
 ANTENNAGATEAREA                          0.216 LAYER ME3 ;
 ANTENNAGATEAREA                          0.216 LAYER ME4 ;
 ANTENNADIFFAREA                          0.160 LAYER ME2 ;
 ANTENNADIFFAREA                          0.160 LAYER ME3 ;
 ANTENNADIFFAREA                          0.160 LAYER ME4 ;
 ANTENNAMAXAREACAR                        7.863 LAYER ME2 ;
 ANTENNAMAXAREACAR                        8.752 LAYER ME3 ;
 ANTENNAMAXAREACAR                        9.641 LAYER ME4 ;
END B4
PIN B3
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 256.780 0.000 257.100 0.600 ;
  LAYER ME3 ;
  RECT 256.780 0.000 257.100 0.600 ;
  LAYER ME2 ;
  RECT 256.780 0.000 257.100 0.600 ;
  LAYER ME1 ;
  RECT 256.780 0.000 257.100 0.600 ;
 END
 ANTENNAPARTIALMETALAREA                  0.984 LAYER ME2 ;
 ANTENNAPARTIALMETALAREA                  0.768 LAYER ME3 ;
 ANTENNAGATEAREA                          0.216 LAYER ME2 ;
 ANTENNAGATEAREA                          0.216 LAYER ME3 ;
 ANTENNAGATEAREA                          0.216 LAYER ME4 ;
 ANTENNADIFFAREA                          0.160 LAYER ME2 ;
 ANTENNADIFFAREA                          0.160 LAYER ME3 ;
 ANTENNADIFFAREA                          0.160 LAYER ME4 ;
 ANTENNAMAXAREACAR                        6.983 LAYER ME2 ;
 ANTENNAMAXAREACAR                       11.428 LAYER ME3 ;
 ANTENNAMAXAREACAR                       12.317 LAYER ME4 ;
END B3
PIN B2
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 260.300 0.000 260.620 0.600 ;
  LAYER ME3 ;
  RECT 260.300 0.000 260.620 0.600 ;
  LAYER ME2 ;
  RECT 260.300 0.000 260.620 0.600 ;
  LAYER ME1 ;
  RECT 260.300 0.000 260.620 0.600 ;
 END
 ANTENNAPARTIALMETALAREA                  0.906 LAYER ME2 ;
 ANTENNAGATEAREA                          0.216 LAYER ME2 ;
 ANTENNAGATEAREA                          0.216 LAYER ME3 ;
 ANTENNAGATEAREA                          0.216 LAYER ME4 ;
 ANTENNADIFFAREA                          0.160 LAYER ME2 ;
 ANTENNADIFFAREA                          0.160 LAYER ME3 ;
 ANTENNADIFFAREA                          0.160 LAYER ME4 ;
 ANTENNAMAXAREACAR                        7.863 LAYER ME2 ;
 ANTENNAMAXAREACAR                        8.752 LAYER ME3 ;
 ANTENNAMAXAREACAR                        9.641 LAYER ME4 ;
END B2
PIN B1
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 270.220 0.000 270.540 0.600 ;
  LAYER ME3 ;
  RECT 270.220 0.000 270.540 0.600 ;
  LAYER ME2 ;
  RECT 270.220 0.000 270.540 0.600 ;
  LAYER ME1 ;
  RECT 270.220 0.000 270.540 0.600 ;
 END
 ANTENNAPARTIALMETALAREA                  0.982 LAYER ME2 ;
 ANTENNAGATEAREA                          0.216 LAYER ME2 ;
 ANTENNAGATEAREA                          0.216 LAYER ME3 ;
 ANTENNAGATEAREA                          0.216 LAYER ME4 ;
 ANTENNADIFFAREA                          0.160 LAYER ME2 ;
 ANTENNADIFFAREA                          0.160 LAYER ME3 ;
 ANTENNADIFFAREA                          0.160 LAYER ME4 ;
 ANTENNAMAXAREACAR                        7.372 LAYER ME2 ;
 ANTENNAMAXAREACAR                        8.261 LAYER ME3 ;
 ANTENNAMAXAREACAR                        9.150 LAYER ME4 ;
END B1
PIN B0
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 281.670 0.000 281.990 0.600 ;
  LAYER ME3 ;
  RECT 281.670 0.000 281.990 0.600 ;
  LAYER ME2 ;
  RECT 281.670 0.000 281.990 0.600 ;
  LAYER ME1 ;
  RECT 281.670 0.000 281.990 0.600 ;
 END
 ANTENNAPARTIALMETALAREA                  1.002 LAYER ME2 ;
 ANTENNAGATEAREA                          0.216 LAYER ME2 ;
 ANTENNAGATEAREA                          0.216 LAYER ME3 ;
 ANTENNAGATEAREA                          0.216 LAYER ME4 ;
 ANTENNADIFFAREA                          0.160 LAYER ME2 ;
 ANTENNADIFFAREA                          0.160 LAYER ME3 ;
 ANTENNADIFFAREA                          0.160 LAYER ME4 ;
 ANTENNAMAXAREACAR                        7.465 LAYER ME2 ;
 ANTENNAMAXAREACAR                        8.354 LAYER ME3 ;
 ANTENNAMAXAREACAR                        9.243 LAYER ME4 ;
END B0
PIN CSBN
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 272.420 0.000 272.740 0.600 ;
  LAYER ME3 ;
  RECT 272.420 0.000 272.740 0.600 ;
  LAYER ME2 ;
  RECT 272.420 0.000 272.740 0.600 ;
  LAYER ME1 ;
  RECT 272.420 0.000 272.740 0.600 ;
 END
 ANTENNAPARTIALMETALAREA                  1.272 LAYER ME2 ;
 ANTENNAPARTIALMETALAREA                  9.794 LAYER ME3 ;
 ANTENNAGATEAREA                          1.896 LAYER ME3 ;
 ANTENNAGATEAREA                          1.896 LAYER ME4 ;
 ANTENNADIFFAREA                          0.160 LAYER ME2 ;
 ANTENNADIFFAREA                          0.160 LAYER ME3 ;
 ANTENNADIFFAREA                          0.160 LAYER ME4 ;
 ANTENNAMAXAREACAR                       37.277 LAYER ME3 ;
 ANTENNAMAXAREACAR                       37.967 LAYER ME4 ;
END CSBN
PIN CKB
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 272.940 0.000 273.260 0.600 ;
  LAYER ME3 ;
  RECT 272.940 0.000 273.260 0.600 ;
  LAYER ME2 ;
  RECT 272.940 0.000 273.260 0.600 ;
  LAYER ME1 ;
  RECT 272.940 0.000 273.260 0.600 ;
 END
 ANTENNAPARTIALMETALAREA                  1.216 LAYER ME2 ;
 ANTENNAPARTIALMETALAREA                 10.394 LAYER ME3 ;
 ANTENNAGATEAREA                          1.632 LAYER ME3 ;
 ANTENNAGATEAREA                          1.632 LAYER ME4 ;
 ANTENNADIFFAREA                          0.160 LAYER ME2 ;
 ANTENNADIFFAREA                          0.160 LAYER ME3 ;
 ANTENNADIFFAREA                          0.160 LAYER ME4 ;
 ANTENNAMAXAREACAR                       46.935 LAYER ME3 ;
 ANTENNAMAXAREACAR                       47.735 LAYER ME4 ;
END CKB
PIN DI35
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 239.140 0.000 239.460 0.600 ;
  LAYER ME3 ;
  RECT 239.140 0.000 239.460 0.600 ;
  LAYER ME2 ;
  RECT 239.140 0.000 239.460 0.600 ;
  LAYER ME1 ;
  RECT 239.140 0.000 239.460 0.600 ;
 END
 ANTENNAPARTIALMETALAREA                  1.918 LAYER ME2 ;
 ANTENNAGATEAREA                          0.101 LAYER ME2 ;
 ANTENNAGATEAREA                          0.101 LAYER ME3 ;
 ANTENNAGATEAREA                          0.101 LAYER ME4 ;
 ANTENNADIFFAREA                          0.160 LAYER ME2 ;
 ANTENNADIFFAREA                          0.160 LAYER ME3 ;
 ANTENNADIFFAREA                          0.160 LAYER ME4 ;
 ANTENNAMAXAREACAR                       22.361 LAYER ME2 ;
 ANTENNAMAXAREACAR                       24.266 LAYER ME3 ;
 ANTENNAMAXAREACAR                       26.171 LAYER ME4 ;
END DI35
PIN DI34
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 232.540 0.000 232.860 0.600 ;
  LAYER ME3 ;
  RECT 232.540 0.000 232.860 0.600 ;
  LAYER ME2 ;
  RECT 232.540 0.000 232.860 0.600 ;
  LAYER ME1 ;
  RECT 232.540 0.000 232.860 0.600 ;
 END
 ANTENNAPARTIALMETALAREA                  1.918 LAYER ME2 ;
 ANTENNAGATEAREA                          0.101 LAYER ME2 ;
 ANTENNAGATEAREA                          0.101 LAYER ME3 ;
 ANTENNAGATEAREA                          0.101 LAYER ME4 ;
 ANTENNADIFFAREA                          0.160 LAYER ME2 ;
 ANTENNADIFFAREA                          0.160 LAYER ME3 ;
 ANTENNADIFFAREA                          0.160 LAYER ME4 ;
 ANTENNAMAXAREACAR                       22.361 LAYER ME2 ;
 ANTENNAMAXAREACAR                       24.266 LAYER ME3 ;
 ANTENNAMAXAREACAR                       26.171 LAYER ME4 ;
END DI34
PIN DI33
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 225.940 0.000 226.260 0.600 ;
  LAYER ME3 ;
  RECT 225.940 0.000 226.260 0.600 ;
  LAYER ME2 ;
  RECT 225.940 0.000 226.260 0.600 ;
  LAYER ME1 ;
  RECT 225.940 0.000 226.260 0.600 ;
 END
 ANTENNAPARTIALMETALAREA                  1.918 LAYER ME2 ;
 ANTENNAGATEAREA                          0.101 LAYER ME2 ;
 ANTENNAGATEAREA                          0.101 LAYER ME3 ;
 ANTENNAGATEAREA                          0.101 LAYER ME4 ;
 ANTENNADIFFAREA                          0.160 LAYER ME2 ;
 ANTENNADIFFAREA                          0.160 LAYER ME3 ;
 ANTENNADIFFAREA                          0.160 LAYER ME4 ;
 ANTENNAMAXAREACAR                       22.361 LAYER ME2 ;
 ANTENNAMAXAREACAR                       24.266 LAYER ME3 ;
 ANTENNAMAXAREACAR                       26.171 LAYER ME4 ;
END DI33
PIN DI32
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 219.340 0.000 219.660 0.600 ;
  LAYER ME3 ;
  RECT 219.340 0.000 219.660 0.600 ;
  LAYER ME2 ;
  RECT 219.340 0.000 219.660 0.600 ;
  LAYER ME1 ;
  RECT 219.340 0.000 219.660 0.600 ;
 END
 ANTENNAPARTIALMETALAREA                  1.918 LAYER ME2 ;
 ANTENNAGATEAREA                          0.101 LAYER ME2 ;
 ANTENNAGATEAREA                          0.101 LAYER ME3 ;
 ANTENNAGATEAREA                          0.101 LAYER ME4 ;
 ANTENNADIFFAREA                          0.160 LAYER ME2 ;
 ANTENNADIFFAREA                          0.160 LAYER ME3 ;
 ANTENNADIFFAREA                          0.160 LAYER ME4 ;
 ANTENNAMAXAREACAR                       22.361 LAYER ME2 ;
 ANTENNAMAXAREACAR                       24.266 LAYER ME3 ;
 ANTENNAMAXAREACAR                       26.171 LAYER ME4 ;
END DI32
PIN DI31
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 212.740 0.000 213.060 0.600 ;
  LAYER ME3 ;
  RECT 212.740 0.000 213.060 0.600 ;
  LAYER ME2 ;
  RECT 212.740 0.000 213.060 0.600 ;
  LAYER ME1 ;
  RECT 212.740 0.000 213.060 0.600 ;
 END
 ANTENNAPARTIALMETALAREA                  1.918 LAYER ME2 ;
 ANTENNAGATEAREA                          0.101 LAYER ME2 ;
 ANTENNAGATEAREA                          0.101 LAYER ME3 ;
 ANTENNAGATEAREA                          0.101 LAYER ME4 ;
 ANTENNADIFFAREA                          0.160 LAYER ME2 ;
 ANTENNADIFFAREA                          0.160 LAYER ME3 ;
 ANTENNADIFFAREA                          0.160 LAYER ME4 ;
 ANTENNAMAXAREACAR                       22.361 LAYER ME2 ;
 ANTENNAMAXAREACAR                       24.266 LAYER ME3 ;
 ANTENNAMAXAREACAR                       26.171 LAYER ME4 ;
END DI31
PIN DI30
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 206.140 0.000 206.460 0.600 ;
  LAYER ME3 ;
  RECT 206.140 0.000 206.460 0.600 ;
  LAYER ME2 ;
  RECT 206.140 0.000 206.460 0.600 ;
  LAYER ME1 ;
  RECT 206.140 0.000 206.460 0.600 ;
 END
 ANTENNAPARTIALMETALAREA                  1.918 LAYER ME2 ;
 ANTENNAGATEAREA                          0.101 LAYER ME2 ;
 ANTENNAGATEAREA                          0.101 LAYER ME3 ;
 ANTENNAGATEAREA                          0.101 LAYER ME4 ;
 ANTENNADIFFAREA                          0.160 LAYER ME2 ;
 ANTENNADIFFAREA                          0.160 LAYER ME3 ;
 ANTENNADIFFAREA                          0.160 LAYER ME4 ;
 ANTENNAMAXAREACAR                       22.361 LAYER ME2 ;
 ANTENNAMAXAREACAR                       24.266 LAYER ME3 ;
 ANTENNAMAXAREACAR                       26.171 LAYER ME4 ;
END DI30
PIN DI29
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 199.540 0.000 199.860 0.600 ;
  LAYER ME3 ;
  RECT 199.540 0.000 199.860 0.600 ;
  LAYER ME2 ;
  RECT 199.540 0.000 199.860 0.600 ;
  LAYER ME1 ;
  RECT 199.540 0.000 199.860 0.600 ;
 END
 ANTENNAPARTIALMETALAREA                  1.918 LAYER ME2 ;
 ANTENNAGATEAREA                          0.101 LAYER ME2 ;
 ANTENNAGATEAREA                          0.101 LAYER ME3 ;
 ANTENNAGATEAREA                          0.101 LAYER ME4 ;
 ANTENNADIFFAREA                          0.160 LAYER ME2 ;
 ANTENNADIFFAREA                          0.160 LAYER ME3 ;
 ANTENNADIFFAREA                          0.160 LAYER ME4 ;
 ANTENNAMAXAREACAR                       22.361 LAYER ME2 ;
 ANTENNAMAXAREACAR                       24.266 LAYER ME3 ;
 ANTENNAMAXAREACAR                       26.171 LAYER ME4 ;
END DI29
PIN DI28
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 192.940 0.000 193.260 0.600 ;
  LAYER ME3 ;
  RECT 192.940 0.000 193.260 0.600 ;
  LAYER ME2 ;
  RECT 192.940 0.000 193.260 0.600 ;
  LAYER ME1 ;
  RECT 192.940 0.000 193.260 0.600 ;
 END
 ANTENNAPARTIALMETALAREA                  1.918 LAYER ME2 ;
 ANTENNAGATEAREA                          0.101 LAYER ME2 ;
 ANTENNAGATEAREA                          0.101 LAYER ME3 ;
 ANTENNAGATEAREA                          0.101 LAYER ME4 ;
 ANTENNADIFFAREA                          0.160 LAYER ME2 ;
 ANTENNADIFFAREA                          0.160 LAYER ME3 ;
 ANTENNADIFFAREA                          0.160 LAYER ME4 ;
 ANTENNAMAXAREACAR                       22.361 LAYER ME2 ;
 ANTENNAMAXAREACAR                       24.266 LAYER ME3 ;
 ANTENNAMAXAREACAR                       26.171 LAYER ME4 ;
END DI28
PIN WEB3
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 180.970 0.000 181.290 0.600 ;
  LAYER ME3 ;
  RECT 180.970 0.000 181.290 0.600 ;
  LAYER ME2 ;
  RECT 180.970 0.000 181.290 0.600 ;
  LAYER ME1 ;
  RECT 180.970 0.000 181.290 0.600 ;
 END
 ANTENNAPARTIALMETALAREA                  0.436 LAYER ME2 ;
 ANTENNAPARTIALMETALAREA                  0.310 LAYER ME3 ;
 ANTENNAGATEAREA                          0.322 LAYER ME2 ;
 ANTENNAGATEAREA                          0.322 LAYER ME3 ;
 ANTENNAGATEAREA                          0.322 LAYER ME4 ;
 ANTENNADIFFAREA                          0.160 LAYER ME2 ;
 ANTENNADIFFAREA                          0.160 LAYER ME3 ;
 ANTENNADIFFAREA                          0.160 LAYER ME4 ;
 ANTENNAMAXAREACAR                        3.197 LAYER ME2 ;
 ANTENNAMAXAREACAR                        4.757 LAYER ME3 ;
 ANTENNAMAXAREACAR                        5.354 LAYER ME4 ;
END WEB3
PIN DI27
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 186.340 0.000 186.660 0.600 ;
  LAYER ME3 ;
  RECT 186.340 0.000 186.660 0.600 ;
  LAYER ME2 ;
  RECT 186.340 0.000 186.660 0.600 ;
  LAYER ME1 ;
  RECT 186.340 0.000 186.660 0.600 ;
 END
 ANTENNAPARTIALMETALAREA                  1.904 LAYER ME2 ;
 ANTENNAGATEAREA                          0.101 LAYER ME2 ;
 ANTENNAGATEAREA                          0.101 LAYER ME3 ;
 ANTENNAGATEAREA                          0.101 LAYER ME4 ;
 ANTENNADIFFAREA                          0.160 LAYER ME2 ;
 ANTENNADIFFAREA                          0.160 LAYER ME3 ;
 ANTENNADIFFAREA                          0.160 LAYER ME4 ;
 ANTENNAMAXAREACAR                       22.222 LAYER ME2 ;
 ANTENNAMAXAREACAR                       24.127 LAYER ME3 ;
 ANTENNAMAXAREACAR                       26.032 LAYER ME4 ;
END DI27
PIN DI26
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 179.740 0.000 180.060 0.600 ;
  LAYER ME3 ;
  RECT 179.740 0.000 180.060 0.600 ;
  LAYER ME2 ;
  RECT 179.740 0.000 180.060 0.600 ;
  LAYER ME1 ;
  RECT 179.740 0.000 180.060 0.600 ;
 END
 ANTENNAPARTIALMETALAREA                  1.918 LAYER ME2 ;
 ANTENNAGATEAREA                          0.101 LAYER ME2 ;
 ANTENNAGATEAREA                          0.101 LAYER ME3 ;
 ANTENNAGATEAREA                          0.101 LAYER ME4 ;
 ANTENNADIFFAREA                          0.160 LAYER ME2 ;
 ANTENNADIFFAREA                          0.160 LAYER ME3 ;
 ANTENNADIFFAREA                          0.160 LAYER ME4 ;
 ANTENNAMAXAREACAR                       22.361 LAYER ME2 ;
 ANTENNAMAXAREACAR                       24.266 LAYER ME3 ;
 ANTENNAMAXAREACAR                       26.171 LAYER ME4 ;
END DI26
PIN DI25
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 173.140 0.000 173.460 0.600 ;
  LAYER ME3 ;
  RECT 173.140 0.000 173.460 0.600 ;
  LAYER ME2 ;
  RECT 173.140 0.000 173.460 0.600 ;
  LAYER ME1 ;
  RECT 173.140 0.000 173.460 0.600 ;
 END
 ANTENNAPARTIALMETALAREA                  1.918 LAYER ME2 ;
 ANTENNAGATEAREA                          0.101 LAYER ME2 ;
 ANTENNAGATEAREA                          0.101 LAYER ME3 ;
 ANTENNAGATEAREA                          0.101 LAYER ME4 ;
 ANTENNADIFFAREA                          0.160 LAYER ME2 ;
 ANTENNADIFFAREA                          0.160 LAYER ME3 ;
 ANTENNADIFFAREA                          0.160 LAYER ME4 ;
 ANTENNAMAXAREACAR                       22.361 LAYER ME2 ;
 ANTENNAMAXAREACAR                       24.266 LAYER ME3 ;
 ANTENNAMAXAREACAR                       26.171 LAYER ME4 ;
END DI25
PIN DI24
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 166.540 0.000 166.860 0.600 ;
  LAYER ME3 ;
  RECT 166.540 0.000 166.860 0.600 ;
  LAYER ME2 ;
  RECT 166.540 0.000 166.860 0.600 ;
  LAYER ME1 ;
  RECT 166.540 0.000 166.860 0.600 ;
 END
 ANTENNAPARTIALMETALAREA                  1.918 LAYER ME2 ;
 ANTENNAGATEAREA                          0.101 LAYER ME2 ;
 ANTENNAGATEAREA                          0.101 LAYER ME3 ;
 ANTENNAGATEAREA                          0.101 LAYER ME4 ;
 ANTENNADIFFAREA                          0.160 LAYER ME2 ;
 ANTENNADIFFAREA                          0.160 LAYER ME3 ;
 ANTENNADIFFAREA                          0.160 LAYER ME4 ;
 ANTENNAMAXAREACAR                       22.361 LAYER ME2 ;
 ANTENNAMAXAREACAR                       24.266 LAYER ME3 ;
 ANTENNAMAXAREACAR                       26.171 LAYER ME4 ;
END DI24
PIN DI23
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 159.940 0.000 160.260 0.600 ;
  LAYER ME3 ;
  RECT 159.940 0.000 160.260 0.600 ;
  LAYER ME2 ;
  RECT 159.940 0.000 160.260 0.600 ;
  LAYER ME1 ;
  RECT 159.940 0.000 160.260 0.600 ;
 END
 ANTENNAPARTIALMETALAREA                  1.918 LAYER ME2 ;
 ANTENNAGATEAREA                          0.101 LAYER ME2 ;
 ANTENNAGATEAREA                          0.101 LAYER ME3 ;
 ANTENNAGATEAREA                          0.101 LAYER ME4 ;
 ANTENNADIFFAREA                          0.160 LAYER ME2 ;
 ANTENNADIFFAREA                          0.160 LAYER ME3 ;
 ANTENNADIFFAREA                          0.160 LAYER ME4 ;
 ANTENNAMAXAREACAR                       22.361 LAYER ME2 ;
 ANTENNAMAXAREACAR                       24.266 LAYER ME3 ;
 ANTENNAMAXAREACAR                       26.171 LAYER ME4 ;
END DI23
PIN DI22
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 153.340 0.000 153.660 0.600 ;
  LAYER ME3 ;
  RECT 153.340 0.000 153.660 0.600 ;
  LAYER ME2 ;
  RECT 153.340 0.000 153.660 0.600 ;
  LAYER ME1 ;
  RECT 153.340 0.000 153.660 0.600 ;
 END
 ANTENNAPARTIALMETALAREA                  1.918 LAYER ME2 ;
 ANTENNAGATEAREA                          0.101 LAYER ME2 ;
 ANTENNAGATEAREA                          0.101 LAYER ME3 ;
 ANTENNAGATEAREA                          0.101 LAYER ME4 ;
 ANTENNADIFFAREA                          0.160 LAYER ME2 ;
 ANTENNADIFFAREA                          0.160 LAYER ME3 ;
 ANTENNADIFFAREA                          0.160 LAYER ME4 ;
 ANTENNAMAXAREACAR                       22.361 LAYER ME2 ;
 ANTENNAMAXAREACAR                       24.266 LAYER ME3 ;
 ANTENNAMAXAREACAR                       26.171 LAYER ME4 ;
END DI22
PIN DI21
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 146.740 0.000 147.060 0.600 ;
  LAYER ME3 ;
  RECT 146.740 0.000 147.060 0.600 ;
  LAYER ME2 ;
  RECT 146.740 0.000 147.060 0.600 ;
  LAYER ME1 ;
  RECT 146.740 0.000 147.060 0.600 ;
 END
 ANTENNAPARTIALMETALAREA                  1.918 LAYER ME2 ;
 ANTENNAGATEAREA                          0.101 LAYER ME2 ;
 ANTENNAGATEAREA                          0.101 LAYER ME3 ;
 ANTENNAGATEAREA                          0.101 LAYER ME4 ;
 ANTENNADIFFAREA                          0.160 LAYER ME2 ;
 ANTENNADIFFAREA                          0.160 LAYER ME3 ;
 ANTENNADIFFAREA                          0.160 LAYER ME4 ;
 ANTENNAMAXAREACAR                       22.361 LAYER ME2 ;
 ANTENNAMAXAREACAR                       24.266 LAYER ME3 ;
 ANTENNAMAXAREACAR                       26.171 LAYER ME4 ;
END DI21
PIN DI20
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 140.140 0.000 140.460 0.600 ;
  LAYER ME3 ;
  RECT 140.140 0.000 140.460 0.600 ;
  LAYER ME2 ;
  RECT 140.140 0.000 140.460 0.600 ;
  LAYER ME1 ;
  RECT 140.140 0.000 140.460 0.600 ;
 END
 ANTENNAPARTIALMETALAREA                  1.918 LAYER ME2 ;
 ANTENNAGATEAREA                          0.101 LAYER ME2 ;
 ANTENNAGATEAREA                          0.101 LAYER ME3 ;
 ANTENNAGATEAREA                          0.101 LAYER ME4 ;
 ANTENNADIFFAREA                          0.160 LAYER ME2 ;
 ANTENNADIFFAREA                          0.160 LAYER ME3 ;
 ANTENNADIFFAREA                          0.160 LAYER ME4 ;
 ANTENNAMAXAREACAR                       22.361 LAYER ME2 ;
 ANTENNAMAXAREACAR                       24.266 LAYER ME3 ;
 ANTENNAMAXAREACAR                       26.171 LAYER ME4 ;
END DI20
PIN DI19
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 133.540 0.000 133.860 0.600 ;
  LAYER ME3 ;
  RECT 133.540 0.000 133.860 0.600 ;
  LAYER ME2 ;
  RECT 133.540 0.000 133.860 0.600 ;
  LAYER ME1 ;
  RECT 133.540 0.000 133.860 0.600 ;
 END
 ANTENNAPARTIALMETALAREA                  1.918 LAYER ME2 ;
 ANTENNAGATEAREA                          0.101 LAYER ME2 ;
 ANTENNAGATEAREA                          0.101 LAYER ME3 ;
 ANTENNAGATEAREA                          0.101 LAYER ME4 ;
 ANTENNADIFFAREA                          0.160 LAYER ME2 ;
 ANTENNADIFFAREA                          0.160 LAYER ME3 ;
 ANTENNADIFFAREA                          0.160 LAYER ME4 ;
 ANTENNAMAXAREACAR                       22.361 LAYER ME2 ;
 ANTENNAMAXAREACAR                       24.266 LAYER ME3 ;
 ANTENNAMAXAREACAR                       26.171 LAYER ME4 ;
END DI19
PIN WEB2
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 121.570 0.000 121.890 0.600 ;
  LAYER ME3 ;
  RECT 121.570 0.000 121.890 0.600 ;
  LAYER ME2 ;
  RECT 121.570 0.000 121.890 0.600 ;
  LAYER ME1 ;
  RECT 121.570 0.000 121.890 0.600 ;
 END
 ANTENNAPARTIALMETALAREA                  0.436 LAYER ME2 ;
 ANTENNAPARTIALMETALAREA                  0.310 LAYER ME3 ;
 ANTENNAGATEAREA                          0.322 LAYER ME2 ;
 ANTENNAGATEAREA                          0.322 LAYER ME3 ;
 ANTENNAGATEAREA                          0.322 LAYER ME4 ;
 ANTENNADIFFAREA                          0.160 LAYER ME2 ;
 ANTENNADIFFAREA                          0.160 LAYER ME3 ;
 ANTENNADIFFAREA                          0.160 LAYER ME4 ;
 ANTENNAMAXAREACAR                        3.197 LAYER ME2 ;
 ANTENNAMAXAREACAR                        4.757 LAYER ME3 ;
 ANTENNAMAXAREACAR                        5.354 LAYER ME4 ;
END WEB2
PIN DI18
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 126.940 0.000 127.260 0.600 ;
  LAYER ME3 ;
  RECT 126.940 0.000 127.260 0.600 ;
  LAYER ME2 ;
  RECT 126.940 0.000 127.260 0.600 ;
  LAYER ME1 ;
  RECT 126.940 0.000 127.260 0.600 ;
 END
 ANTENNAPARTIALMETALAREA                  1.904 LAYER ME2 ;
 ANTENNAGATEAREA                          0.101 LAYER ME2 ;
 ANTENNAGATEAREA                          0.101 LAYER ME3 ;
 ANTENNAGATEAREA                          0.101 LAYER ME4 ;
 ANTENNADIFFAREA                          0.160 LAYER ME2 ;
 ANTENNADIFFAREA                          0.160 LAYER ME3 ;
 ANTENNADIFFAREA                          0.160 LAYER ME4 ;
 ANTENNAMAXAREACAR                       22.222 LAYER ME2 ;
 ANTENNAMAXAREACAR                       24.127 LAYER ME3 ;
 ANTENNAMAXAREACAR                       26.032 LAYER ME4 ;
END DI18
PIN DI17
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 120.340 0.000 120.660 0.600 ;
  LAYER ME3 ;
  RECT 120.340 0.000 120.660 0.600 ;
  LAYER ME2 ;
  RECT 120.340 0.000 120.660 0.600 ;
  LAYER ME1 ;
  RECT 120.340 0.000 120.660 0.600 ;
 END
 ANTENNAPARTIALMETALAREA                  1.918 LAYER ME2 ;
 ANTENNAGATEAREA                          0.101 LAYER ME2 ;
 ANTENNAGATEAREA                          0.101 LAYER ME3 ;
 ANTENNAGATEAREA                          0.101 LAYER ME4 ;
 ANTENNADIFFAREA                          0.160 LAYER ME2 ;
 ANTENNADIFFAREA                          0.160 LAYER ME3 ;
 ANTENNADIFFAREA                          0.160 LAYER ME4 ;
 ANTENNAMAXAREACAR                       22.361 LAYER ME2 ;
 ANTENNAMAXAREACAR                       24.266 LAYER ME3 ;
 ANTENNAMAXAREACAR                       26.171 LAYER ME4 ;
END DI17
PIN DI16
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 113.740 0.000 114.060 0.600 ;
  LAYER ME3 ;
  RECT 113.740 0.000 114.060 0.600 ;
  LAYER ME2 ;
  RECT 113.740 0.000 114.060 0.600 ;
  LAYER ME1 ;
  RECT 113.740 0.000 114.060 0.600 ;
 END
 ANTENNAPARTIALMETALAREA                  1.918 LAYER ME2 ;
 ANTENNAGATEAREA                          0.101 LAYER ME2 ;
 ANTENNAGATEAREA                          0.101 LAYER ME3 ;
 ANTENNAGATEAREA                          0.101 LAYER ME4 ;
 ANTENNADIFFAREA                          0.160 LAYER ME2 ;
 ANTENNADIFFAREA                          0.160 LAYER ME3 ;
 ANTENNADIFFAREA                          0.160 LAYER ME4 ;
 ANTENNAMAXAREACAR                       22.361 LAYER ME2 ;
 ANTENNAMAXAREACAR                       24.266 LAYER ME3 ;
 ANTENNAMAXAREACAR                       26.171 LAYER ME4 ;
END DI16
PIN DI15
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 107.140 0.000 107.460 0.600 ;
  LAYER ME3 ;
  RECT 107.140 0.000 107.460 0.600 ;
  LAYER ME2 ;
  RECT 107.140 0.000 107.460 0.600 ;
  LAYER ME1 ;
  RECT 107.140 0.000 107.460 0.600 ;
 END
 ANTENNAPARTIALMETALAREA                  1.918 LAYER ME2 ;
 ANTENNAGATEAREA                          0.101 LAYER ME2 ;
 ANTENNAGATEAREA                          0.101 LAYER ME3 ;
 ANTENNAGATEAREA                          0.101 LAYER ME4 ;
 ANTENNADIFFAREA                          0.160 LAYER ME2 ;
 ANTENNADIFFAREA                          0.160 LAYER ME3 ;
 ANTENNADIFFAREA                          0.160 LAYER ME4 ;
 ANTENNAMAXAREACAR                       22.361 LAYER ME2 ;
 ANTENNAMAXAREACAR                       24.266 LAYER ME3 ;
 ANTENNAMAXAREACAR                       26.171 LAYER ME4 ;
END DI15
PIN DI14
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 100.540 0.000 100.860 0.600 ;
  LAYER ME3 ;
  RECT 100.540 0.000 100.860 0.600 ;
  LAYER ME2 ;
  RECT 100.540 0.000 100.860 0.600 ;
  LAYER ME1 ;
  RECT 100.540 0.000 100.860 0.600 ;
 END
 ANTENNAPARTIALMETALAREA                  1.918 LAYER ME2 ;
 ANTENNAGATEAREA                          0.101 LAYER ME2 ;
 ANTENNAGATEAREA                          0.101 LAYER ME3 ;
 ANTENNAGATEAREA                          0.101 LAYER ME4 ;
 ANTENNADIFFAREA                          0.160 LAYER ME2 ;
 ANTENNADIFFAREA                          0.160 LAYER ME3 ;
 ANTENNADIFFAREA                          0.160 LAYER ME4 ;
 ANTENNAMAXAREACAR                       22.361 LAYER ME2 ;
 ANTENNAMAXAREACAR                       24.266 LAYER ME3 ;
 ANTENNAMAXAREACAR                       26.171 LAYER ME4 ;
END DI14
PIN DI13
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 93.940 0.000 94.260 0.600 ;
  LAYER ME3 ;
  RECT 93.940 0.000 94.260 0.600 ;
  LAYER ME2 ;
  RECT 93.940 0.000 94.260 0.600 ;
  LAYER ME1 ;
  RECT 93.940 0.000 94.260 0.600 ;
 END
 ANTENNAPARTIALMETALAREA                  1.918 LAYER ME2 ;
 ANTENNAGATEAREA                          0.101 LAYER ME2 ;
 ANTENNAGATEAREA                          0.101 LAYER ME3 ;
 ANTENNAGATEAREA                          0.101 LAYER ME4 ;
 ANTENNADIFFAREA                          0.160 LAYER ME2 ;
 ANTENNADIFFAREA                          0.160 LAYER ME3 ;
 ANTENNADIFFAREA                          0.160 LAYER ME4 ;
 ANTENNAMAXAREACAR                       22.361 LAYER ME2 ;
 ANTENNAMAXAREACAR                       24.266 LAYER ME3 ;
 ANTENNAMAXAREACAR                       26.171 LAYER ME4 ;
END DI13
PIN DI12
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 87.340 0.000 87.660 0.600 ;
  LAYER ME3 ;
  RECT 87.340 0.000 87.660 0.600 ;
  LAYER ME2 ;
  RECT 87.340 0.000 87.660 0.600 ;
  LAYER ME1 ;
  RECT 87.340 0.000 87.660 0.600 ;
 END
 ANTENNAPARTIALMETALAREA                  1.918 LAYER ME2 ;
 ANTENNAGATEAREA                          0.101 LAYER ME2 ;
 ANTENNAGATEAREA                          0.101 LAYER ME3 ;
 ANTENNAGATEAREA                          0.101 LAYER ME4 ;
 ANTENNADIFFAREA                          0.160 LAYER ME2 ;
 ANTENNADIFFAREA                          0.160 LAYER ME3 ;
 ANTENNADIFFAREA                          0.160 LAYER ME4 ;
 ANTENNAMAXAREACAR                       22.361 LAYER ME2 ;
 ANTENNAMAXAREACAR                       24.266 LAYER ME3 ;
 ANTENNAMAXAREACAR                       26.171 LAYER ME4 ;
END DI12
PIN DI11
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 80.740 0.000 81.060 0.600 ;
  LAYER ME3 ;
  RECT 80.740 0.000 81.060 0.600 ;
  LAYER ME2 ;
  RECT 80.740 0.000 81.060 0.600 ;
  LAYER ME1 ;
  RECT 80.740 0.000 81.060 0.600 ;
 END
 ANTENNAPARTIALMETALAREA                  1.918 LAYER ME2 ;
 ANTENNAGATEAREA                          0.101 LAYER ME2 ;
 ANTENNAGATEAREA                          0.101 LAYER ME3 ;
 ANTENNAGATEAREA                          0.101 LAYER ME4 ;
 ANTENNADIFFAREA                          0.160 LAYER ME2 ;
 ANTENNADIFFAREA                          0.160 LAYER ME3 ;
 ANTENNADIFFAREA                          0.160 LAYER ME4 ;
 ANTENNAMAXAREACAR                       22.361 LAYER ME2 ;
 ANTENNAMAXAREACAR                       24.266 LAYER ME3 ;
 ANTENNAMAXAREACAR                       26.171 LAYER ME4 ;
END DI11
PIN DI10
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 74.140 0.000 74.460 0.600 ;
  LAYER ME3 ;
  RECT 74.140 0.000 74.460 0.600 ;
  LAYER ME2 ;
  RECT 74.140 0.000 74.460 0.600 ;
  LAYER ME1 ;
  RECT 74.140 0.000 74.460 0.600 ;
 END
 ANTENNAPARTIALMETALAREA                  1.918 LAYER ME2 ;
 ANTENNAGATEAREA                          0.101 LAYER ME2 ;
 ANTENNAGATEAREA                          0.101 LAYER ME3 ;
 ANTENNAGATEAREA                          0.101 LAYER ME4 ;
 ANTENNADIFFAREA                          0.160 LAYER ME2 ;
 ANTENNADIFFAREA                          0.160 LAYER ME3 ;
 ANTENNADIFFAREA                          0.160 LAYER ME4 ;
 ANTENNAMAXAREACAR                       22.361 LAYER ME2 ;
 ANTENNAMAXAREACAR                       24.266 LAYER ME3 ;
 ANTENNAMAXAREACAR                       26.171 LAYER ME4 ;
END DI10
PIN WEB1
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 62.170 0.000 62.490 0.600 ;
  LAYER ME3 ;
  RECT 62.170 0.000 62.490 0.600 ;
  LAYER ME2 ;
  RECT 62.170 0.000 62.490 0.600 ;
  LAYER ME1 ;
  RECT 62.170 0.000 62.490 0.600 ;
 END
 ANTENNAPARTIALMETALAREA                  0.436 LAYER ME2 ;
 ANTENNAPARTIALMETALAREA                  0.310 LAYER ME3 ;
 ANTENNAGATEAREA                          0.322 LAYER ME2 ;
 ANTENNAGATEAREA                          0.322 LAYER ME3 ;
 ANTENNAGATEAREA                          0.322 LAYER ME4 ;
 ANTENNADIFFAREA                          0.160 LAYER ME2 ;
 ANTENNADIFFAREA                          0.160 LAYER ME3 ;
 ANTENNADIFFAREA                          0.160 LAYER ME4 ;
 ANTENNAMAXAREACAR                        3.197 LAYER ME2 ;
 ANTENNAMAXAREACAR                        4.757 LAYER ME3 ;
 ANTENNAMAXAREACAR                        5.354 LAYER ME4 ;
END WEB1
PIN DI9
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 67.540 0.000 67.860 0.600 ;
  LAYER ME3 ;
  RECT 67.540 0.000 67.860 0.600 ;
  LAYER ME2 ;
  RECT 67.540 0.000 67.860 0.600 ;
  LAYER ME1 ;
  RECT 67.540 0.000 67.860 0.600 ;
 END
 ANTENNAPARTIALMETALAREA                  1.904 LAYER ME2 ;
 ANTENNAGATEAREA                          0.101 LAYER ME2 ;
 ANTENNAGATEAREA                          0.101 LAYER ME3 ;
 ANTENNAGATEAREA                          0.101 LAYER ME4 ;
 ANTENNADIFFAREA                          0.160 LAYER ME2 ;
 ANTENNADIFFAREA                          0.160 LAYER ME3 ;
 ANTENNADIFFAREA                          0.160 LAYER ME4 ;
 ANTENNAMAXAREACAR                       22.222 LAYER ME2 ;
 ANTENNAMAXAREACAR                       24.127 LAYER ME3 ;
 ANTENNAMAXAREACAR                       26.032 LAYER ME4 ;
END DI9
PIN DI8
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 60.940 0.000 61.260 0.600 ;
  LAYER ME3 ;
  RECT 60.940 0.000 61.260 0.600 ;
  LAYER ME2 ;
  RECT 60.940 0.000 61.260 0.600 ;
  LAYER ME1 ;
  RECT 60.940 0.000 61.260 0.600 ;
 END
 ANTENNAPARTIALMETALAREA                  1.918 LAYER ME2 ;
 ANTENNAGATEAREA                          0.101 LAYER ME2 ;
 ANTENNAGATEAREA                          0.101 LAYER ME3 ;
 ANTENNAGATEAREA                          0.101 LAYER ME4 ;
 ANTENNADIFFAREA                          0.160 LAYER ME2 ;
 ANTENNADIFFAREA                          0.160 LAYER ME3 ;
 ANTENNADIFFAREA                          0.160 LAYER ME4 ;
 ANTENNAMAXAREACAR                       22.361 LAYER ME2 ;
 ANTENNAMAXAREACAR                       24.266 LAYER ME3 ;
 ANTENNAMAXAREACAR                       26.171 LAYER ME4 ;
END DI8
PIN DI7
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 54.340 0.000 54.660 0.600 ;
  LAYER ME3 ;
  RECT 54.340 0.000 54.660 0.600 ;
  LAYER ME2 ;
  RECT 54.340 0.000 54.660 0.600 ;
  LAYER ME1 ;
  RECT 54.340 0.000 54.660 0.600 ;
 END
 ANTENNAPARTIALMETALAREA                  1.918 LAYER ME2 ;
 ANTENNAGATEAREA                          0.101 LAYER ME2 ;
 ANTENNAGATEAREA                          0.101 LAYER ME3 ;
 ANTENNAGATEAREA                          0.101 LAYER ME4 ;
 ANTENNADIFFAREA                          0.160 LAYER ME2 ;
 ANTENNADIFFAREA                          0.160 LAYER ME3 ;
 ANTENNADIFFAREA                          0.160 LAYER ME4 ;
 ANTENNAMAXAREACAR                       22.361 LAYER ME2 ;
 ANTENNAMAXAREACAR                       24.266 LAYER ME3 ;
 ANTENNAMAXAREACAR                       26.171 LAYER ME4 ;
END DI7
PIN DI6
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 47.740 0.000 48.060 0.600 ;
  LAYER ME3 ;
  RECT 47.740 0.000 48.060 0.600 ;
  LAYER ME2 ;
  RECT 47.740 0.000 48.060 0.600 ;
  LAYER ME1 ;
  RECT 47.740 0.000 48.060 0.600 ;
 END
 ANTENNAPARTIALMETALAREA                  1.918 LAYER ME2 ;
 ANTENNAGATEAREA                          0.101 LAYER ME2 ;
 ANTENNAGATEAREA                          0.101 LAYER ME3 ;
 ANTENNAGATEAREA                          0.101 LAYER ME4 ;
 ANTENNADIFFAREA                          0.160 LAYER ME2 ;
 ANTENNADIFFAREA                          0.160 LAYER ME3 ;
 ANTENNADIFFAREA                          0.160 LAYER ME4 ;
 ANTENNAMAXAREACAR                       22.361 LAYER ME2 ;
 ANTENNAMAXAREACAR                       24.266 LAYER ME3 ;
 ANTENNAMAXAREACAR                       26.171 LAYER ME4 ;
END DI6
PIN DI5
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 41.140 0.000 41.460 0.600 ;
  LAYER ME3 ;
  RECT 41.140 0.000 41.460 0.600 ;
  LAYER ME2 ;
  RECT 41.140 0.000 41.460 0.600 ;
  LAYER ME1 ;
  RECT 41.140 0.000 41.460 0.600 ;
 END
 ANTENNAPARTIALMETALAREA                  1.918 LAYER ME2 ;
 ANTENNAGATEAREA                          0.101 LAYER ME2 ;
 ANTENNAGATEAREA                          0.101 LAYER ME3 ;
 ANTENNAGATEAREA                          0.101 LAYER ME4 ;
 ANTENNADIFFAREA                          0.160 LAYER ME2 ;
 ANTENNADIFFAREA                          0.160 LAYER ME3 ;
 ANTENNADIFFAREA                          0.160 LAYER ME4 ;
 ANTENNAMAXAREACAR                       22.361 LAYER ME2 ;
 ANTENNAMAXAREACAR                       24.266 LAYER ME3 ;
 ANTENNAMAXAREACAR                       26.171 LAYER ME4 ;
END DI5
PIN DI4
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 34.540 0.000 34.860 0.600 ;
  LAYER ME3 ;
  RECT 34.540 0.000 34.860 0.600 ;
  LAYER ME2 ;
  RECT 34.540 0.000 34.860 0.600 ;
  LAYER ME1 ;
  RECT 34.540 0.000 34.860 0.600 ;
 END
 ANTENNAPARTIALMETALAREA                  1.918 LAYER ME2 ;
 ANTENNAGATEAREA                          0.101 LAYER ME2 ;
 ANTENNAGATEAREA                          0.101 LAYER ME3 ;
 ANTENNAGATEAREA                          0.101 LAYER ME4 ;
 ANTENNADIFFAREA                          0.160 LAYER ME2 ;
 ANTENNADIFFAREA                          0.160 LAYER ME3 ;
 ANTENNADIFFAREA                          0.160 LAYER ME4 ;
 ANTENNAMAXAREACAR                       22.361 LAYER ME2 ;
 ANTENNAMAXAREACAR                       24.266 LAYER ME3 ;
 ANTENNAMAXAREACAR                       26.171 LAYER ME4 ;
END DI4
PIN DI3
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 27.940 0.000 28.260 0.600 ;
  LAYER ME3 ;
  RECT 27.940 0.000 28.260 0.600 ;
  LAYER ME2 ;
  RECT 27.940 0.000 28.260 0.600 ;
  LAYER ME1 ;
  RECT 27.940 0.000 28.260 0.600 ;
 END
 ANTENNAPARTIALMETALAREA                  1.918 LAYER ME2 ;
 ANTENNAGATEAREA                          0.101 LAYER ME2 ;
 ANTENNAGATEAREA                          0.101 LAYER ME3 ;
 ANTENNAGATEAREA                          0.101 LAYER ME4 ;
 ANTENNADIFFAREA                          0.160 LAYER ME2 ;
 ANTENNADIFFAREA                          0.160 LAYER ME3 ;
 ANTENNADIFFAREA                          0.160 LAYER ME4 ;
 ANTENNAMAXAREACAR                       22.361 LAYER ME2 ;
 ANTENNAMAXAREACAR                       24.266 LAYER ME3 ;
 ANTENNAMAXAREACAR                       26.171 LAYER ME4 ;
END DI3
PIN DI2
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 21.340 0.000 21.660 0.600 ;
  LAYER ME3 ;
  RECT 21.340 0.000 21.660 0.600 ;
  LAYER ME2 ;
  RECT 21.340 0.000 21.660 0.600 ;
  LAYER ME1 ;
  RECT 21.340 0.000 21.660 0.600 ;
 END
 ANTENNAPARTIALMETALAREA                  1.918 LAYER ME2 ;
 ANTENNAGATEAREA                          0.101 LAYER ME2 ;
 ANTENNAGATEAREA                          0.101 LAYER ME3 ;
 ANTENNAGATEAREA                          0.101 LAYER ME4 ;
 ANTENNADIFFAREA                          0.160 LAYER ME2 ;
 ANTENNADIFFAREA                          0.160 LAYER ME3 ;
 ANTENNADIFFAREA                          0.160 LAYER ME4 ;
 ANTENNAMAXAREACAR                       22.361 LAYER ME2 ;
 ANTENNAMAXAREACAR                       24.266 LAYER ME3 ;
 ANTENNAMAXAREACAR                       26.171 LAYER ME4 ;
END DI2
PIN DI1
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 14.740 0.000 15.060 0.600 ;
  LAYER ME3 ;
  RECT 14.740 0.000 15.060 0.600 ;
  LAYER ME2 ;
  RECT 14.740 0.000 15.060 0.600 ;
  LAYER ME1 ;
  RECT 14.740 0.000 15.060 0.600 ;
 END
 ANTENNAPARTIALMETALAREA                  1.918 LAYER ME2 ;
 ANTENNAGATEAREA                          0.101 LAYER ME2 ;
 ANTENNAGATEAREA                          0.101 LAYER ME3 ;
 ANTENNAGATEAREA                          0.101 LAYER ME4 ;
 ANTENNADIFFAREA                          0.160 LAYER ME2 ;
 ANTENNADIFFAREA                          0.160 LAYER ME3 ;
 ANTENNADIFFAREA                          0.160 LAYER ME4 ;
 ANTENNAMAXAREACAR                       22.361 LAYER ME2 ;
 ANTENNAMAXAREACAR                       24.266 LAYER ME3 ;
 ANTENNAMAXAREACAR                       26.171 LAYER ME4 ;
END DI1
PIN WEB0
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 2.770 0.000 3.090 0.600 ;
  LAYER ME3 ;
  RECT 2.770 0.000 3.090 0.600 ;
  LAYER ME2 ;
  RECT 2.770 0.000 3.090 0.600 ;
  LAYER ME1 ;
  RECT 2.770 0.000 3.090 0.600 ;
 END
 ANTENNAPARTIALMETALAREA                  0.436 LAYER ME2 ;
 ANTENNAPARTIALMETALAREA                  0.310 LAYER ME3 ;
 ANTENNAGATEAREA                          0.322 LAYER ME2 ;
 ANTENNAGATEAREA                          0.322 LAYER ME3 ;
 ANTENNAGATEAREA                          0.322 LAYER ME4 ;
 ANTENNADIFFAREA                          0.160 LAYER ME2 ;
 ANTENNADIFFAREA                          0.160 LAYER ME3 ;
 ANTENNADIFFAREA                          0.160 LAYER ME4 ;
 ANTENNAMAXAREACAR                        3.197 LAYER ME2 ;
 ANTENNAMAXAREACAR                        4.757 LAYER ME3 ;
 ANTENNAMAXAREACAR                        5.354 LAYER ME4 ;
END WEB0
PIN DI0
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 8.140 0.000 8.460 0.600 ;
  LAYER ME3 ;
  RECT 8.140 0.000 8.460 0.600 ;
  LAYER ME2 ;
  RECT 8.140 0.000 8.460 0.600 ;
  LAYER ME1 ;
  RECT 8.140 0.000 8.460 0.600 ;
 END
 ANTENNAPARTIALMETALAREA                  1.904 LAYER ME2 ;
 ANTENNAGATEAREA                          0.101 LAYER ME2 ;
 ANTENNAGATEAREA                          0.101 LAYER ME3 ;
 ANTENNAGATEAREA                          0.101 LAYER ME4 ;
 ANTENNADIFFAREA                          0.160 LAYER ME2 ;
 ANTENNADIFFAREA                          0.160 LAYER ME3 ;
 ANTENNADIFFAREA                          0.160 LAYER ME4 ;
 ANTENNAMAXAREACAR                       22.222 LAYER ME2 ;
 ANTENNAMAXAREACAR                       24.127 LAYER ME3 ;
 ANTENNAMAXAREACAR                       26.032 LAYER ME4 ;
END DI0
PIN DI71
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 536.350 0.000 536.670 0.600 ;
  LAYER ME3 ;
  RECT 536.350 0.000 536.670 0.600 ;
  LAYER ME2 ;
  RECT 536.350 0.000 536.670 0.600 ;
  LAYER ME1 ;
  RECT 536.350 0.000 536.670 0.600 ;
 END
 ANTENNAPARTIALMETALAREA                  1.918 LAYER ME2 ;
 ANTENNAGATEAREA                          0.101 LAYER ME2 ;
 ANTENNAGATEAREA                          0.101 LAYER ME3 ;
 ANTENNAGATEAREA                          0.101 LAYER ME4 ;
 ANTENNADIFFAREA                          0.160 LAYER ME2 ;
 ANTENNADIFFAREA                          0.160 LAYER ME3 ;
 ANTENNADIFFAREA                          0.160 LAYER ME4 ;
 ANTENNAMAXAREACAR                       22.361 LAYER ME2 ;
 ANTENNAMAXAREACAR                       24.266 LAYER ME3 ;
 ANTENNAMAXAREACAR                       26.171 LAYER ME4 ;
END DI71
PIN DI70
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 529.750 0.000 530.070 0.600 ;
  LAYER ME3 ;
  RECT 529.750 0.000 530.070 0.600 ;
  LAYER ME2 ;
  RECT 529.750 0.000 530.070 0.600 ;
  LAYER ME1 ;
  RECT 529.750 0.000 530.070 0.600 ;
 END
 ANTENNAPARTIALMETALAREA                  1.918 LAYER ME2 ;
 ANTENNAGATEAREA                          0.101 LAYER ME2 ;
 ANTENNAGATEAREA                          0.101 LAYER ME3 ;
 ANTENNAGATEAREA                          0.101 LAYER ME4 ;
 ANTENNADIFFAREA                          0.160 LAYER ME2 ;
 ANTENNADIFFAREA                          0.160 LAYER ME3 ;
 ANTENNADIFFAREA                          0.160 LAYER ME4 ;
 ANTENNAMAXAREACAR                       22.361 LAYER ME2 ;
 ANTENNAMAXAREACAR                       24.266 LAYER ME3 ;
 ANTENNAMAXAREACAR                       26.171 LAYER ME4 ;
END DI70
PIN DI69
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 523.150 0.000 523.470 0.600 ;
  LAYER ME3 ;
  RECT 523.150 0.000 523.470 0.600 ;
  LAYER ME2 ;
  RECT 523.150 0.000 523.470 0.600 ;
  LAYER ME1 ;
  RECT 523.150 0.000 523.470 0.600 ;
 END
 ANTENNAPARTIALMETALAREA                  1.918 LAYER ME2 ;
 ANTENNAGATEAREA                          0.101 LAYER ME2 ;
 ANTENNAGATEAREA                          0.101 LAYER ME3 ;
 ANTENNAGATEAREA                          0.101 LAYER ME4 ;
 ANTENNADIFFAREA                          0.160 LAYER ME2 ;
 ANTENNADIFFAREA                          0.160 LAYER ME3 ;
 ANTENNADIFFAREA                          0.160 LAYER ME4 ;
 ANTENNAMAXAREACAR                       22.361 LAYER ME2 ;
 ANTENNAMAXAREACAR                       24.266 LAYER ME3 ;
 ANTENNAMAXAREACAR                       26.171 LAYER ME4 ;
END DI69
PIN DI68
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 516.550 0.000 516.870 0.600 ;
  LAYER ME3 ;
  RECT 516.550 0.000 516.870 0.600 ;
  LAYER ME2 ;
  RECT 516.550 0.000 516.870 0.600 ;
  LAYER ME1 ;
  RECT 516.550 0.000 516.870 0.600 ;
 END
 ANTENNAPARTIALMETALAREA                  1.918 LAYER ME2 ;
 ANTENNAGATEAREA                          0.101 LAYER ME2 ;
 ANTENNAGATEAREA                          0.101 LAYER ME3 ;
 ANTENNAGATEAREA                          0.101 LAYER ME4 ;
 ANTENNADIFFAREA                          0.160 LAYER ME2 ;
 ANTENNADIFFAREA                          0.160 LAYER ME3 ;
 ANTENNADIFFAREA                          0.160 LAYER ME4 ;
 ANTENNAMAXAREACAR                       22.361 LAYER ME2 ;
 ANTENNAMAXAREACAR                       24.266 LAYER ME3 ;
 ANTENNAMAXAREACAR                       26.171 LAYER ME4 ;
END DI68
PIN DI67
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 509.950 0.000 510.270 0.600 ;
  LAYER ME3 ;
  RECT 509.950 0.000 510.270 0.600 ;
  LAYER ME2 ;
  RECT 509.950 0.000 510.270 0.600 ;
  LAYER ME1 ;
  RECT 509.950 0.000 510.270 0.600 ;
 END
 ANTENNAPARTIALMETALAREA                  1.918 LAYER ME2 ;
 ANTENNAGATEAREA                          0.101 LAYER ME2 ;
 ANTENNAGATEAREA                          0.101 LAYER ME3 ;
 ANTENNAGATEAREA                          0.101 LAYER ME4 ;
 ANTENNADIFFAREA                          0.160 LAYER ME2 ;
 ANTENNADIFFAREA                          0.160 LAYER ME3 ;
 ANTENNADIFFAREA                          0.160 LAYER ME4 ;
 ANTENNAMAXAREACAR                       22.361 LAYER ME2 ;
 ANTENNAMAXAREACAR                       24.266 LAYER ME3 ;
 ANTENNAMAXAREACAR                       26.171 LAYER ME4 ;
END DI67
PIN DI66
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 503.350 0.000 503.670 0.600 ;
  LAYER ME3 ;
  RECT 503.350 0.000 503.670 0.600 ;
  LAYER ME2 ;
  RECT 503.350 0.000 503.670 0.600 ;
  LAYER ME1 ;
  RECT 503.350 0.000 503.670 0.600 ;
 END
 ANTENNAPARTIALMETALAREA                  1.918 LAYER ME2 ;
 ANTENNAGATEAREA                          0.101 LAYER ME2 ;
 ANTENNAGATEAREA                          0.101 LAYER ME3 ;
 ANTENNAGATEAREA                          0.101 LAYER ME4 ;
 ANTENNADIFFAREA                          0.160 LAYER ME2 ;
 ANTENNADIFFAREA                          0.160 LAYER ME3 ;
 ANTENNADIFFAREA                          0.160 LAYER ME4 ;
 ANTENNAMAXAREACAR                       22.361 LAYER ME2 ;
 ANTENNAMAXAREACAR                       24.266 LAYER ME3 ;
 ANTENNAMAXAREACAR                       26.171 LAYER ME4 ;
END DI66
PIN DI65
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 496.750 0.000 497.070 0.600 ;
  LAYER ME3 ;
  RECT 496.750 0.000 497.070 0.600 ;
  LAYER ME2 ;
  RECT 496.750 0.000 497.070 0.600 ;
  LAYER ME1 ;
  RECT 496.750 0.000 497.070 0.600 ;
 END
 ANTENNAPARTIALMETALAREA                  1.918 LAYER ME2 ;
 ANTENNAGATEAREA                          0.101 LAYER ME2 ;
 ANTENNAGATEAREA                          0.101 LAYER ME3 ;
 ANTENNAGATEAREA                          0.101 LAYER ME4 ;
 ANTENNADIFFAREA                          0.160 LAYER ME2 ;
 ANTENNADIFFAREA                          0.160 LAYER ME3 ;
 ANTENNADIFFAREA                          0.160 LAYER ME4 ;
 ANTENNAMAXAREACAR                       22.361 LAYER ME2 ;
 ANTENNAMAXAREACAR                       24.266 LAYER ME3 ;
 ANTENNAMAXAREACAR                       26.171 LAYER ME4 ;
END DI65
PIN DI64
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 490.150 0.000 490.470 0.600 ;
  LAYER ME3 ;
  RECT 490.150 0.000 490.470 0.600 ;
  LAYER ME2 ;
  RECT 490.150 0.000 490.470 0.600 ;
  LAYER ME1 ;
  RECT 490.150 0.000 490.470 0.600 ;
 END
 ANTENNAPARTIALMETALAREA                  1.918 LAYER ME2 ;
 ANTENNAGATEAREA                          0.101 LAYER ME2 ;
 ANTENNAGATEAREA                          0.101 LAYER ME3 ;
 ANTENNAGATEAREA                          0.101 LAYER ME4 ;
 ANTENNADIFFAREA                          0.160 LAYER ME2 ;
 ANTENNADIFFAREA                          0.160 LAYER ME3 ;
 ANTENNADIFFAREA                          0.160 LAYER ME4 ;
 ANTENNAMAXAREACAR                       22.361 LAYER ME2 ;
 ANTENNAMAXAREACAR                       24.266 LAYER ME3 ;
 ANTENNAMAXAREACAR                       26.171 LAYER ME4 ;
END DI64
PIN DI63
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 483.550 0.000 483.870 0.600 ;
  LAYER ME3 ;
  RECT 483.550 0.000 483.870 0.600 ;
  LAYER ME2 ;
  RECT 483.550 0.000 483.870 0.600 ;
  LAYER ME1 ;
  RECT 483.550 0.000 483.870 0.600 ;
 END
 ANTENNAPARTIALMETALAREA                  1.904 LAYER ME2 ;
 ANTENNAGATEAREA                          0.101 LAYER ME2 ;
 ANTENNAGATEAREA                          0.101 LAYER ME3 ;
 ANTENNAGATEAREA                          0.101 LAYER ME4 ;
 ANTENNADIFFAREA                          0.160 LAYER ME2 ;
 ANTENNADIFFAREA                          0.160 LAYER ME3 ;
 ANTENNADIFFAREA                          0.160 LAYER ME4 ;
 ANTENNAMAXAREACAR                       22.222 LAYER ME2 ;
 ANTENNAMAXAREACAR                       24.127 LAYER ME3 ;
 ANTENNAMAXAREACAR                       26.032 LAYER ME4 ;
END DI63
PIN WEB7
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 478.180 0.000 478.500 0.600 ;
  LAYER ME3 ;
  RECT 478.180 0.000 478.500 0.600 ;
  LAYER ME2 ;
  RECT 478.180 0.000 478.500 0.600 ;
  LAYER ME1 ;
  RECT 478.180 0.000 478.500 0.600 ;
 END
 ANTENNAPARTIALMETALAREA                  0.436 LAYER ME2 ;
 ANTENNAPARTIALMETALAREA                  0.310 LAYER ME3 ;
 ANTENNAGATEAREA                          0.322 LAYER ME2 ;
 ANTENNAGATEAREA                          0.322 LAYER ME3 ;
 ANTENNAGATEAREA                          0.322 LAYER ME4 ;
 ANTENNADIFFAREA                          0.160 LAYER ME2 ;
 ANTENNADIFFAREA                          0.160 LAYER ME3 ;
 ANTENNADIFFAREA                          0.160 LAYER ME4 ;
 ANTENNAMAXAREACAR                        3.197 LAYER ME2 ;
 ANTENNAMAXAREACAR                        4.757 LAYER ME3 ;
 ANTENNAMAXAREACAR                        5.354 LAYER ME4 ;
END WEB7
PIN DI62
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 476.950 0.000 477.270 0.600 ;
  LAYER ME3 ;
  RECT 476.950 0.000 477.270 0.600 ;
  LAYER ME2 ;
  RECT 476.950 0.000 477.270 0.600 ;
  LAYER ME1 ;
  RECT 476.950 0.000 477.270 0.600 ;
 END
 ANTENNAPARTIALMETALAREA                  1.918 LAYER ME2 ;
 ANTENNAGATEAREA                          0.101 LAYER ME2 ;
 ANTENNAGATEAREA                          0.101 LAYER ME3 ;
 ANTENNAGATEAREA                          0.101 LAYER ME4 ;
 ANTENNADIFFAREA                          0.160 LAYER ME2 ;
 ANTENNADIFFAREA                          0.160 LAYER ME3 ;
 ANTENNADIFFAREA                          0.160 LAYER ME4 ;
 ANTENNAMAXAREACAR                       22.361 LAYER ME2 ;
 ANTENNAMAXAREACAR                       24.266 LAYER ME3 ;
 ANTENNAMAXAREACAR                       26.171 LAYER ME4 ;
END DI62
PIN DI61
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 470.350 0.000 470.670 0.600 ;
  LAYER ME3 ;
  RECT 470.350 0.000 470.670 0.600 ;
  LAYER ME2 ;
  RECT 470.350 0.000 470.670 0.600 ;
  LAYER ME1 ;
  RECT 470.350 0.000 470.670 0.600 ;
 END
 ANTENNAPARTIALMETALAREA                  1.918 LAYER ME2 ;
 ANTENNAGATEAREA                          0.101 LAYER ME2 ;
 ANTENNAGATEAREA                          0.101 LAYER ME3 ;
 ANTENNAGATEAREA                          0.101 LAYER ME4 ;
 ANTENNADIFFAREA                          0.160 LAYER ME2 ;
 ANTENNADIFFAREA                          0.160 LAYER ME3 ;
 ANTENNADIFFAREA                          0.160 LAYER ME4 ;
 ANTENNAMAXAREACAR                       22.361 LAYER ME2 ;
 ANTENNAMAXAREACAR                       24.266 LAYER ME3 ;
 ANTENNAMAXAREACAR                       26.171 LAYER ME4 ;
END DI61
PIN DI60
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 463.750 0.000 464.070 0.600 ;
  LAYER ME3 ;
  RECT 463.750 0.000 464.070 0.600 ;
  LAYER ME2 ;
  RECT 463.750 0.000 464.070 0.600 ;
  LAYER ME1 ;
  RECT 463.750 0.000 464.070 0.600 ;
 END
 ANTENNAPARTIALMETALAREA                  1.918 LAYER ME2 ;
 ANTENNAGATEAREA                          0.101 LAYER ME2 ;
 ANTENNAGATEAREA                          0.101 LAYER ME3 ;
 ANTENNAGATEAREA                          0.101 LAYER ME4 ;
 ANTENNADIFFAREA                          0.160 LAYER ME2 ;
 ANTENNADIFFAREA                          0.160 LAYER ME3 ;
 ANTENNADIFFAREA                          0.160 LAYER ME4 ;
 ANTENNAMAXAREACAR                       22.361 LAYER ME2 ;
 ANTENNAMAXAREACAR                       24.266 LAYER ME3 ;
 ANTENNAMAXAREACAR                       26.171 LAYER ME4 ;
END DI60
PIN DI59
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 457.150 0.000 457.470 0.600 ;
  LAYER ME3 ;
  RECT 457.150 0.000 457.470 0.600 ;
  LAYER ME2 ;
  RECT 457.150 0.000 457.470 0.600 ;
  LAYER ME1 ;
  RECT 457.150 0.000 457.470 0.600 ;
 END
 ANTENNAPARTIALMETALAREA                  1.918 LAYER ME2 ;
 ANTENNAGATEAREA                          0.101 LAYER ME2 ;
 ANTENNAGATEAREA                          0.101 LAYER ME3 ;
 ANTENNAGATEAREA                          0.101 LAYER ME4 ;
 ANTENNADIFFAREA                          0.160 LAYER ME2 ;
 ANTENNADIFFAREA                          0.160 LAYER ME3 ;
 ANTENNADIFFAREA                          0.160 LAYER ME4 ;
 ANTENNAMAXAREACAR                       22.361 LAYER ME2 ;
 ANTENNAMAXAREACAR                       24.266 LAYER ME3 ;
 ANTENNAMAXAREACAR                       26.171 LAYER ME4 ;
END DI59
PIN DI58
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 450.550 0.000 450.870 0.600 ;
  LAYER ME3 ;
  RECT 450.550 0.000 450.870 0.600 ;
  LAYER ME2 ;
  RECT 450.550 0.000 450.870 0.600 ;
  LAYER ME1 ;
  RECT 450.550 0.000 450.870 0.600 ;
 END
 ANTENNAPARTIALMETALAREA                  1.918 LAYER ME2 ;
 ANTENNAGATEAREA                          0.101 LAYER ME2 ;
 ANTENNAGATEAREA                          0.101 LAYER ME3 ;
 ANTENNAGATEAREA                          0.101 LAYER ME4 ;
 ANTENNADIFFAREA                          0.160 LAYER ME2 ;
 ANTENNADIFFAREA                          0.160 LAYER ME3 ;
 ANTENNADIFFAREA                          0.160 LAYER ME4 ;
 ANTENNAMAXAREACAR                       22.361 LAYER ME2 ;
 ANTENNAMAXAREACAR                       24.266 LAYER ME3 ;
 ANTENNAMAXAREACAR                       26.171 LAYER ME4 ;
END DI58
PIN DI57
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 443.950 0.000 444.270 0.600 ;
  LAYER ME3 ;
  RECT 443.950 0.000 444.270 0.600 ;
  LAYER ME2 ;
  RECT 443.950 0.000 444.270 0.600 ;
  LAYER ME1 ;
  RECT 443.950 0.000 444.270 0.600 ;
 END
 ANTENNAPARTIALMETALAREA                  1.918 LAYER ME2 ;
 ANTENNAGATEAREA                          0.101 LAYER ME2 ;
 ANTENNAGATEAREA                          0.101 LAYER ME3 ;
 ANTENNAGATEAREA                          0.101 LAYER ME4 ;
 ANTENNADIFFAREA                          0.160 LAYER ME2 ;
 ANTENNADIFFAREA                          0.160 LAYER ME3 ;
 ANTENNADIFFAREA                          0.160 LAYER ME4 ;
 ANTENNAMAXAREACAR                       22.361 LAYER ME2 ;
 ANTENNAMAXAREACAR                       24.266 LAYER ME3 ;
 ANTENNAMAXAREACAR                       26.171 LAYER ME4 ;
END DI57
PIN DI56
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 437.350 0.000 437.670 0.600 ;
  LAYER ME3 ;
  RECT 437.350 0.000 437.670 0.600 ;
  LAYER ME2 ;
  RECT 437.350 0.000 437.670 0.600 ;
  LAYER ME1 ;
  RECT 437.350 0.000 437.670 0.600 ;
 END
 ANTENNAPARTIALMETALAREA                  1.918 LAYER ME2 ;
 ANTENNAGATEAREA                          0.101 LAYER ME2 ;
 ANTENNAGATEAREA                          0.101 LAYER ME3 ;
 ANTENNAGATEAREA                          0.101 LAYER ME4 ;
 ANTENNADIFFAREA                          0.160 LAYER ME2 ;
 ANTENNADIFFAREA                          0.160 LAYER ME3 ;
 ANTENNADIFFAREA                          0.160 LAYER ME4 ;
 ANTENNAMAXAREACAR                       22.361 LAYER ME2 ;
 ANTENNAMAXAREACAR                       24.266 LAYER ME3 ;
 ANTENNAMAXAREACAR                       26.171 LAYER ME4 ;
END DI56
PIN DI55
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 430.750 0.000 431.070 0.600 ;
  LAYER ME3 ;
  RECT 430.750 0.000 431.070 0.600 ;
  LAYER ME2 ;
  RECT 430.750 0.000 431.070 0.600 ;
  LAYER ME1 ;
  RECT 430.750 0.000 431.070 0.600 ;
 END
 ANTENNAPARTIALMETALAREA                  1.918 LAYER ME2 ;
 ANTENNAGATEAREA                          0.101 LAYER ME2 ;
 ANTENNAGATEAREA                          0.101 LAYER ME3 ;
 ANTENNAGATEAREA                          0.101 LAYER ME4 ;
 ANTENNADIFFAREA                          0.160 LAYER ME2 ;
 ANTENNADIFFAREA                          0.160 LAYER ME3 ;
 ANTENNADIFFAREA                          0.160 LAYER ME4 ;
 ANTENNAMAXAREACAR                       22.361 LAYER ME2 ;
 ANTENNAMAXAREACAR                       24.266 LAYER ME3 ;
 ANTENNAMAXAREACAR                       26.171 LAYER ME4 ;
END DI55
PIN DI54
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 424.150 0.000 424.470 0.600 ;
  LAYER ME3 ;
  RECT 424.150 0.000 424.470 0.600 ;
  LAYER ME2 ;
  RECT 424.150 0.000 424.470 0.600 ;
  LAYER ME1 ;
  RECT 424.150 0.000 424.470 0.600 ;
 END
 ANTENNAPARTIALMETALAREA                  1.904 LAYER ME2 ;
 ANTENNAGATEAREA                          0.101 LAYER ME2 ;
 ANTENNAGATEAREA                          0.101 LAYER ME3 ;
 ANTENNAGATEAREA                          0.101 LAYER ME4 ;
 ANTENNADIFFAREA                          0.160 LAYER ME2 ;
 ANTENNADIFFAREA                          0.160 LAYER ME3 ;
 ANTENNADIFFAREA                          0.160 LAYER ME4 ;
 ANTENNAMAXAREACAR                       22.222 LAYER ME2 ;
 ANTENNAMAXAREACAR                       24.127 LAYER ME3 ;
 ANTENNAMAXAREACAR                       26.032 LAYER ME4 ;
END DI54
PIN WEB6
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 418.780 0.000 419.100 0.600 ;
  LAYER ME3 ;
  RECT 418.780 0.000 419.100 0.600 ;
  LAYER ME2 ;
  RECT 418.780 0.000 419.100 0.600 ;
  LAYER ME1 ;
  RECT 418.780 0.000 419.100 0.600 ;
 END
 ANTENNAPARTIALMETALAREA                  0.436 LAYER ME2 ;
 ANTENNAPARTIALMETALAREA                  0.310 LAYER ME3 ;
 ANTENNAGATEAREA                          0.322 LAYER ME2 ;
 ANTENNAGATEAREA                          0.322 LAYER ME3 ;
 ANTENNAGATEAREA                          0.322 LAYER ME4 ;
 ANTENNADIFFAREA                          0.160 LAYER ME2 ;
 ANTENNADIFFAREA                          0.160 LAYER ME3 ;
 ANTENNADIFFAREA                          0.160 LAYER ME4 ;
 ANTENNAMAXAREACAR                        3.197 LAYER ME2 ;
 ANTENNAMAXAREACAR                        4.757 LAYER ME3 ;
 ANTENNAMAXAREACAR                        5.354 LAYER ME4 ;
END WEB6
PIN DI53
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 417.550 0.000 417.870 0.600 ;
  LAYER ME3 ;
  RECT 417.550 0.000 417.870 0.600 ;
  LAYER ME2 ;
  RECT 417.550 0.000 417.870 0.600 ;
  LAYER ME1 ;
  RECT 417.550 0.000 417.870 0.600 ;
 END
 ANTENNAPARTIALMETALAREA                  1.918 LAYER ME2 ;
 ANTENNAGATEAREA                          0.101 LAYER ME2 ;
 ANTENNAGATEAREA                          0.101 LAYER ME3 ;
 ANTENNAGATEAREA                          0.101 LAYER ME4 ;
 ANTENNADIFFAREA                          0.160 LAYER ME2 ;
 ANTENNADIFFAREA                          0.160 LAYER ME3 ;
 ANTENNADIFFAREA                          0.160 LAYER ME4 ;
 ANTENNAMAXAREACAR                       22.361 LAYER ME2 ;
 ANTENNAMAXAREACAR                       24.266 LAYER ME3 ;
 ANTENNAMAXAREACAR                       26.171 LAYER ME4 ;
END DI53
PIN DI52
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 410.950 0.000 411.270 0.600 ;
  LAYER ME3 ;
  RECT 410.950 0.000 411.270 0.600 ;
  LAYER ME2 ;
  RECT 410.950 0.000 411.270 0.600 ;
  LAYER ME1 ;
  RECT 410.950 0.000 411.270 0.600 ;
 END
 ANTENNAPARTIALMETALAREA                  1.918 LAYER ME2 ;
 ANTENNAGATEAREA                          0.101 LAYER ME2 ;
 ANTENNAGATEAREA                          0.101 LAYER ME3 ;
 ANTENNAGATEAREA                          0.101 LAYER ME4 ;
 ANTENNADIFFAREA                          0.160 LAYER ME2 ;
 ANTENNADIFFAREA                          0.160 LAYER ME3 ;
 ANTENNADIFFAREA                          0.160 LAYER ME4 ;
 ANTENNAMAXAREACAR                       22.361 LAYER ME2 ;
 ANTENNAMAXAREACAR                       24.266 LAYER ME3 ;
 ANTENNAMAXAREACAR                       26.171 LAYER ME4 ;
END DI52
PIN DI51
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 404.350 0.000 404.670 0.600 ;
  LAYER ME3 ;
  RECT 404.350 0.000 404.670 0.600 ;
  LAYER ME2 ;
  RECT 404.350 0.000 404.670 0.600 ;
  LAYER ME1 ;
  RECT 404.350 0.000 404.670 0.600 ;
 END
 ANTENNAPARTIALMETALAREA                  1.918 LAYER ME2 ;
 ANTENNAGATEAREA                          0.101 LAYER ME2 ;
 ANTENNAGATEAREA                          0.101 LAYER ME3 ;
 ANTENNAGATEAREA                          0.101 LAYER ME4 ;
 ANTENNADIFFAREA                          0.160 LAYER ME2 ;
 ANTENNADIFFAREA                          0.160 LAYER ME3 ;
 ANTENNADIFFAREA                          0.160 LAYER ME4 ;
 ANTENNAMAXAREACAR                       22.361 LAYER ME2 ;
 ANTENNAMAXAREACAR                       24.266 LAYER ME3 ;
 ANTENNAMAXAREACAR                       26.171 LAYER ME4 ;
END DI51
PIN DI50
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 397.750 0.000 398.070 0.600 ;
  LAYER ME3 ;
  RECT 397.750 0.000 398.070 0.600 ;
  LAYER ME2 ;
  RECT 397.750 0.000 398.070 0.600 ;
  LAYER ME1 ;
  RECT 397.750 0.000 398.070 0.600 ;
 END
 ANTENNAPARTIALMETALAREA                  1.918 LAYER ME2 ;
 ANTENNAGATEAREA                          0.101 LAYER ME2 ;
 ANTENNAGATEAREA                          0.101 LAYER ME3 ;
 ANTENNAGATEAREA                          0.101 LAYER ME4 ;
 ANTENNADIFFAREA                          0.160 LAYER ME2 ;
 ANTENNADIFFAREA                          0.160 LAYER ME3 ;
 ANTENNADIFFAREA                          0.160 LAYER ME4 ;
 ANTENNAMAXAREACAR                       22.361 LAYER ME2 ;
 ANTENNAMAXAREACAR                       24.266 LAYER ME3 ;
 ANTENNAMAXAREACAR                       26.171 LAYER ME4 ;
END DI50
PIN DI49
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 391.150 0.000 391.470 0.600 ;
  LAYER ME3 ;
  RECT 391.150 0.000 391.470 0.600 ;
  LAYER ME2 ;
  RECT 391.150 0.000 391.470 0.600 ;
  LAYER ME1 ;
  RECT 391.150 0.000 391.470 0.600 ;
 END
 ANTENNAPARTIALMETALAREA                  1.918 LAYER ME2 ;
 ANTENNAGATEAREA                          0.101 LAYER ME2 ;
 ANTENNAGATEAREA                          0.101 LAYER ME3 ;
 ANTENNAGATEAREA                          0.101 LAYER ME4 ;
 ANTENNADIFFAREA                          0.160 LAYER ME2 ;
 ANTENNADIFFAREA                          0.160 LAYER ME3 ;
 ANTENNADIFFAREA                          0.160 LAYER ME4 ;
 ANTENNAMAXAREACAR                       22.361 LAYER ME2 ;
 ANTENNAMAXAREACAR                       24.266 LAYER ME3 ;
 ANTENNAMAXAREACAR                       26.171 LAYER ME4 ;
END DI49
PIN DI48
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 384.550 0.000 384.870 0.600 ;
  LAYER ME3 ;
  RECT 384.550 0.000 384.870 0.600 ;
  LAYER ME2 ;
  RECT 384.550 0.000 384.870 0.600 ;
  LAYER ME1 ;
  RECT 384.550 0.000 384.870 0.600 ;
 END
 ANTENNAPARTIALMETALAREA                  1.918 LAYER ME2 ;
 ANTENNAGATEAREA                          0.101 LAYER ME2 ;
 ANTENNAGATEAREA                          0.101 LAYER ME3 ;
 ANTENNAGATEAREA                          0.101 LAYER ME4 ;
 ANTENNADIFFAREA                          0.160 LAYER ME2 ;
 ANTENNADIFFAREA                          0.160 LAYER ME3 ;
 ANTENNADIFFAREA                          0.160 LAYER ME4 ;
 ANTENNAMAXAREACAR                       22.361 LAYER ME2 ;
 ANTENNAMAXAREACAR                       24.266 LAYER ME3 ;
 ANTENNAMAXAREACAR                       26.171 LAYER ME4 ;
END DI48
PIN DI47
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 377.950 0.000 378.270 0.600 ;
  LAYER ME3 ;
  RECT 377.950 0.000 378.270 0.600 ;
  LAYER ME2 ;
  RECT 377.950 0.000 378.270 0.600 ;
  LAYER ME1 ;
  RECT 377.950 0.000 378.270 0.600 ;
 END
 ANTENNAPARTIALMETALAREA                  1.918 LAYER ME2 ;
 ANTENNAGATEAREA                          0.101 LAYER ME2 ;
 ANTENNAGATEAREA                          0.101 LAYER ME3 ;
 ANTENNAGATEAREA                          0.101 LAYER ME4 ;
 ANTENNADIFFAREA                          0.160 LAYER ME2 ;
 ANTENNADIFFAREA                          0.160 LAYER ME3 ;
 ANTENNADIFFAREA                          0.160 LAYER ME4 ;
 ANTENNAMAXAREACAR                       22.361 LAYER ME2 ;
 ANTENNAMAXAREACAR                       24.266 LAYER ME3 ;
 ANTENNAMAXAREACAR                       26.171 LAYER ME4 ;
END DI47
PIN DI46
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 371.350 0.000 371.670 0.600 ;
  LAYER ME3 ;
  RECT 371.350 0.000 371.670 0.600 ;
  LAYER ME2 ;
  RECT 371.350 0.000 371.670 0.600 ;
  LAYER ME1 ;
  RECT 371.350 0.000 371.670 0.600 ;
 END
 ANTENNAPARTIALMETALAREA                  1.918 LAYER ME2 ;
 ANTENNAGATEAREA                          0.101 LAYER ME2 ;
 ANTENNAGATEAREA                          0.101 LAYER ME3 ;
 ANTENNAGATEAREA                          0.101 LAYER ME4 ;
 ANTENNADIFFAREA                          0.160 LAYER ME2 ;
 ANTENNADIFFAREA                          0.160 LAYER ME3 ;
 ANTENNADIFFAREA                          0.160 LAYER ME4 ;
 ANTENNAMAXAREACAR                       22.361 LAYER ME2 ;
 ANTENNAMAXAREACAR                       24.266 LAYER ME3 ;
 ANTENNAMAXAREACAR                       26.171 LAYER ME4 ;
END DI46
PIN DI45
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 364.750 0.000 365.070 0.600 ;
  LAYER ME3 ;
  RECT 364.750 0.000 365.070 0.600 ;
  LAYER ME2 ;
  RECT 364.750 0.000 365.070 0.600 ;
  LAYER ME1 ;
  RECT 364.750 0.000 365.070 0.600 ;
 END
 ANTENNAPARTIALMETALAREA                  1.904 LAYER ME2 ;
 ANTENNAGATEAREA                          0.101 LAYER ME2 ;
 ANTENNAGATEAREA                          0.101 LAYER ME3 ;
 ANTENNAGATEAREA                          0.101 LAYER ME4 ;
 ANTENNADIFFAREA                          0.160 LAYER ME2 ;
 ANTENNADIFFAREA                          0.160 LAYER ME3 ;
 ANTENNADIFFAREA                          0.160 LAYER ME4 ;
 ANTENNAMAXAREACAR                       22.222 LAYER ME2 ;
 ANTENNAMAXAREACAR                       24.127 LAYER ME3 ;
 ANTENNAMAXAREACAR                       26.032 LAYER ME4 ;
END DI45
PIN WEB5
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 359.380 0.000 359.700 0.600 ;
  LAYER ME3 ;
  RECT 359.380 0.000 359.700 0.600 ;
  LAYER ME2 ;
  RECT 359.380 0.000 359.700 0.600 ;
  LAYER ME1 ;
  RECT 359.380 0.000 359.700 0.600 ;
 END
 ANTENNAPARTIALMETALAREA                  0.436 LAYER ME2 ;
 ANTENNAPARTIALMETALAREA                  0.310 LAYER ME3 ;
 ANTENNAGATEAREA                          0.322 LAYER ME2 ;
 ANTENNAGATEAREA                          0.322 LAYER ME3 ;
 ANTENNAGATEAREA                          0.322 LAYER ME4 ;
 ANTENNADIFFAREA                          0.160 LAYER ME2 ;
 ANTENNADIFFAREA                          0.160 LAYER ME3 ;
 ANTENNADIFFAREA                          0.160 LAYER ME4 ;
 ANTENNAMAXAREACAR                        3.197 LAYER ME2 ;
 ANTENNAMAXAREACAR                        4.757 LAYER ME3 ;
 ANTENNAMAXAREACAR                        5.354 LAYER ME4 ;
END WEB5
PIN DI44
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 358.150 0.000 358.470 0.600 ;
  LAYER ME3 ;
  RECT 358.150 0.000 358.470 0.600 ;
  LAYER ME2 ;
  RECT 358.150 0.000 358.470 0.600 ;
  LAYER ME1 ;
  RECT 358.150 0.000 358.470 0.600 ;
 END
 ANTENNAPARTIALMETALAREA                  1.918 LAYER ME2 ;
 ANTENNAGATEAREA                          0.101 LAYER ME2 ;
 ANTENNAGATEAREA                          0.101 LAYER ME3 ;
 ANTENNAGATEAREA                          0.101 LAYER ME4 ;
 ANTENNADIFFAREA                          0.160 LAYER ME2 ;
 ANTENNADIFFAREA                          0.160 LAYER ME3 ;
 ANTENNADIFFAREA                          0.160 LAYER ME4 ;
 ANTENNAMAXAREACAR                       22.361 LAYER ME2 ;
 ANTENNAMAXAREACAR                       24.266 LAYER ME3 ;
 ANTENNAMAXAREACAR                       26.171 LAYER ME4 ;
END DI44
PIN DI43
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 351.550 0.000 351.870 0.600 ;
  LAYER ME3 ;
  RECT 351.550 0.000 351.870 0.600 ;
  LAYER ME2 ;
  RECT 351.550 0.000 351.870 0.600 ;
  LAYER ME1 ;
  RECT 351.550 0.000 351.870 0.600 ;
 END
 ANTENNAPARTIALMETALAREA                  1.918 LAYER ME2 ;
 ANTENNAGATEAREA                          0.101 LAYER ME2 ;
 ANTENNAGATEAREA                          0.101 LAYER ME3 ;
 ANTENNAGATEAREA                          0.101 LAYER ME4 ;
 ANTENNADIFFAREA                          0.160 LAYER ME2 ;
 ANTENNADIFFAREA                          0.160 LAYER ME3 ;
 ANTENNADIFFAREA                          0.160 LAYER ME4 ;
 ANTENNAMAXAREACAR                       22.361 LAYER ME2 ;
 ANTENNAMAXAREACAR                       24.266 LAYER ME3 ;
 ANTENNAMAXAREACAR                       26.171 LAYER ME4 ;
END DI43
PIN DI42
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 344.950 0.000 345.270 0.600 ;
  LAYER ME3 ;
  RECT 344.950 0.000 345.270 0.600 ;
  LAYER ME2 ;
  RECT 344.950 0.000 345.270 0.600 ;
  LAYER ME1 ;
  RECT 344.950 0.000 345.270 0.600 ;
 END
 ANTENNAPARTIALMETALAREA                  1.918 LAYER ME2 ;
 ANTENNAGATEAREA                          0.101 LAYER ME2 ;
 ANTENNAGATEAREA                          0.101 LAYER ME3 ;
 ANTENNAGATEAREA                          0.101 LAYER ME4 ;
 ANTENNADIFFAREA                          0.160 LAYER ME2 ;
 ANTENNADIFFAREA                          0.160 LAYER ME3 ;
 ANTENNADIFFAREA                          0.160 LAYER ME4 ;
 ANTENNAMAXAREACAR                       22.361 LAYER ME2 ;
 ANTENNAMAXAREACAR                       24.266 LAYER ME3 ;
 ANTENNAMAXAREACAR                       26.171 LAYER ME4 ;
END DI42
PIN DI41
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 338.350 0.000 338.670 0.600 ;
  LAYER ME3 ;
  RECT 338.350 0.000 338.670 0.600 ;
  LAYER ME2 ;
  RECT 338.350 0.000 338.670 0.600 ;
  LAYER ME1 ;
  RECT 338.350 0.000 338.670 0.600 ;
 END
 ANTENNAPARTIALMETALAREA                  1.918 LAYER ME2 ;
 ANTENNAGATEAREA                          0.101 LAYER ME2 ;
 ANTENNAGATEAREA                          0.101 LAYER ME3 ;
 ANTENNAGATEAREA                          0.101 LAYER ME4 ;
 ANTENNADIFFAREA                          0.160 LAYER ME2 ;
 ANTENNADIFFAREA                          0.160 LAYER ME3 ;
 ANTENNADIFFAREA                          0.160 LAYER ME4 ;
 ANTENNAMAXAREACAR                       22.361 LAYER ME2 ;
 ANTENNAMAXAREACAR                       24.266 LAYER ME3 ;
 ANTENNAMAXAREACAR                       26.171 LAYER ME4 ;
END DI41
PIN DI40
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 331.750 0.000 332.070 0.600 ;
  LAYER ME3 ;
  RECT 331.750 0.000 332.070 0.600 ;
  LAYER ME2 ;
  RECT 331.750 0.000 332.070 0.600 ;
  LAYER ME1 ;
  RECT 331.750 0.000 332.070 0.600 ;
 END
 ANTENNAPARTIALMETALAREA                  1.918 LAYER ME2 ;
 ANTENNAGATEAREA                          0.101 LAYER ME2 ;
 ANTENNAGATEAREA                          0.101 LAYER ME3 ;
 ANTENNAGATEAREA                          0.101 LAYER ME4 ;
 ANTENNADIFFAREA                          0.160 LAYER ME2 ;
 ANTENNADIFFAREA                          0.160 LAYER ME3 ;
 ANTENNADIFFAREA                          0.160 LAYER ME4 ;
 ANTENNAMAXAREACAR                       22.361 LAYER ME2 ;
 ANTENNAMAXAREACAR                       24.266 LAYER ME3 ;
 ANTENNAMAXAREACAR                       26.171 LAYER ME4 ;
END DI40
PIN DI39
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 325.150 0.000 325.470 0.600 ;
  LAYER ME3 ;
  RECT 325.150 0.000 325.470 0.600 ;
  LAYER ME2 ;
  RECT 325.150 0.000 325.470 0.600 ;
  LAYER ME1 ;
  RECT 325.150 0.000 325.470 0.600 ;
 END
 ANTENNAPARTIALMETALAREA                  1.918 LAYER ME2 ;
 ANTENNAGATEAREA                          0.101 LAYER ME2 ;
 ANTENNAGATEAREA                          0.101 LAYER ME3 ;
 ANTENNAGATEAREA                          0.101 LAYER ME4 ;
 ANTENNADIFFAREA                          0.160 LAYER ME2 ;
 ANTENNADIFFAREA                          0.160 LAYER ME3 ;
 ANTENNADIFFAREA                          0.160 LAYER ME4 ;
 ANTENNAMAXAREACAR                       22.361 LAYER ME2 ;
 ANTENNAMAXAREACAR                       24.266 LAYER ME3 ;
 ANTENNAMAXAREACAR                       26.171 LAYER ME4 ;
END DI39
PIN DI38
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 318.550 0.000 318.870 0.600 ;
  LAYER ME3 ;
  RECT 318.550 0.000 318.870 0.600 ;
  LAYER ME2 ;
  RECT 318.550 0.000 318.870 0.600 ;
  LAYER ME1 ;
  RECT 318.550 0.000 318.870 0.600 ;
 END
 ANTENNAPARTIALMETALAREA                  1.918 LAYER ME2 ;
 ANTENNAGATEAREA                          0.101 LAYER ME2 ;
 ANTENNAGATEAREA                          0.101 LAYER ME3 ;
 ANTENNAGATEAREA                          0.101 LAYER ME4 ;
 ANTENNADIFFAREA                          0.160 LAYER ME2 ;
 ANTENNADIFFAREA                          0.160 LAYER ME3 ;
 ANTENNADIFFAREA                          0.160 LAYER ME4 ;
 ANTENNAMAXAREACAR                       22.361 LAYER ME2 ;
 ANTENNAMAXAREACAR                       24.266 LAYER ME3 ;
 ANTENNAMAXAREACAR                       26.171 LAYER ME4 ;
END DI38
PIN DI37
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 311.950 0.000 312.270 0.600 ;
  LAYER ME3 ;
  RECT 311.950 0.000 312.270 0.600 ;
  LAYER ME2 ;
  RECT 311.950 0.000 312.270 0.600 ;
  LAYER ME1 ;
  RECT 311.950 0.000 312.270 0.600 ;
 END
 ANTENNAPARTIALMETALAREA                  1.918 LAYER ME2 ;
 ANTENNAGATEAREA                          0.101 LAYER ME2 ;
 ANTENNAGATEAREA                          0.101 LAYER ME3 ;
 ANTENNAGATEAREA                          0.101 LAYER ME4 ;
 ANTENNADIFFAREA                          0.160 LAYER ME2 ;
 ANTENNADIFFAREA                          0.160 LAYER ME3 ;
 ANTENNADIFFAREA                          0.160 LAYER ME4 ;
 ANTENNAMAXAREACAR                       22.361 LAYER ME2 ;
 ANTENNAMAXAREACAR                       24.266 LAYER ME3 ;
 ANTENNAMAXAREACAR                       26.171 LAYER ME4 ;
END DI37
PIN DI36
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 305.350 0.000 305.670 0.600 ;
  LAYER ME3 ;
  RECT 305.350 0.000 305.670 0.600 ;
  LAYER ME2 ;
  RECT 305.350 0.000 305.670 0.600 ;
  LAYER ME1 ;
  RECT 305.350 0.000 305.670 0.600 ;
 END
 ANTENNAPARTIALMETALAREA                  1.904 LAYER ME2 ;
 ANTENNAGATEAREA                          0.101 LAYER ME2 ;
 ANTENNAGATEAREA                          0.101 LAYER ME3 ;
 ANTENNAGATEAREA                          0.101 LAYER ME4 ;
 ANTENNADIFFAREA                          0.160 LAYER ME2 ;
 ANTENNADIFFAREA                          0.160 LAYER ME3 ;
 ANTENNADIFFAREA                          0.160 LAYER ME4 ;
 ANTENNAMAXAREACAR                       22.222 LAYER ME2 ;
 ANTENNAMAXAREACAR                       24.127 LAYER ME3 ;
 ANTENNAMAXAREACAR                       26.032 LAYER ME4 ;
END DI36
PIN WEB4
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 299.980 0.000 300.300 0.600 ;
  LAYER ME3 ;
  RECT 299.980 0.000 300.300 0.600 ;
  LAYER ME2 ;
  RECT 299.980 0.000 300.300 0.600 ;
  LAYER ME1 ;
  RECT 299.980 0.000 300.300 0.600 ;
 END
 ANTENNAPARTIALMETALAREA                  0.436 LAYER ME2 ;
 ANTENNAPARTIALMETALAREA                  0.310 LAYER ME3 ;
 ANTENNAGATEAREA                          0.322 LAYER ME2 ;
 ANTENNAGATEAREA                          0.322 LAYER ME3 ;
 ANTENNAGATEAREA                          0.322 LAYER ME4 ;
 ANTENNADIFFAREA                          0.160 LAYER ME2 ;
 ANTENNADIFFAREA                          0.160 LAYER ME3 ;
 ANTENNADIFFAREA                          0.160 LAYER ME4 ;
 ANTENNAMAXAREACAR                        3.197 LAYER ME2 ;
 ANTENNAMAXAREACAR                        4.757 LAYER ME3 ;
 ANTENNAMAXAREACAR                        5.354 LAYER ME4 ;
END WEB4
OBS
  LAYER ME4 ;
  RECT 0.000 0.000 539.250 221.080 ;
  LAYER ME3 ;
  RECT 0.000 0.000 539.250 221.080 ;
  LAYER ME2 ;
  RECT 0.000 0.000 539.250 221.080 ;
  LAYER ME1 ;
  RECT 0.000 0.000 539.250 221.080 ;
END
END SZKD110_256X9X8CM2
END LIBRARY





