# ________________________________________________________________________________________________
# 
# 
#             Synchronous One-Port Register File Compiler
# 
#                 UMC 0.11um LL AE Logic Process
# 
# ________________________________________________________________________________________________
# 
#               
#         Copyright (C) 2024 Faraday Technology Corporation. All Rights Reserved.       
#                
#         This source code is an unpublished work belongs to Faraday Technology Corporation       
#         It is considered a trade secret and is not to be divulged or       
#         used by parties who have not received written authorization from       
#         Faraday Technology Corporation       
#                
#         Faraday's home page can be found at: http://www.faraday-tech.com/       
#                
# ________________________________________________________________________________________________
# 
#        IP Name            :  FSR0K_B_SY                
#        IP Version         :  1.4.0                     
#        IP Release Status  :  Active                    
#        Word               :  512                       
#        Bit                :  16                        
#        Byte               :  8                         
#        Mux                :  2                         
#        Output Loading     :  0.01                      
#        Clock Input Slew   :  0.016                     
#        Data Input Slew    :  0.016                     
#        Ring Type          :  Ringless Model            
#        Ring Width         :  0                         
#        Bus Format         :  0                         
#        Memaker Path       :  /home/mem/Desktop/memlib  
#        GUI Version        :  m20230904                 
#        Date               :  2024/09/23 13:16:55       
# ________________________________________________________________________________________________
# 

VERSION 5.5 ;
NAMESCASESENSITIVE ON ;
MACRO SYKB110_512X16X8CM2
CLASS BLOCK ;
FOREIGN SYKB110_512X16X8CM2 0.000 0.000 ;
ORIGIN 0.000 0.000 ;
SIZE 557.611 BY 293.175 ;
SYMMETRY x y r90 ;
SITE core ;
PIN GND
  DIRECTION INOUT ;
  USE GROUND ;
 PORT
  LAYER ME4 ;
  RECT 302.278 1.781 302.618 293.175 ;
 END
 PORT
  LAYER ME4 ;
  RECT 298.274 1.781 298.614 293.175 ;
 END
 PORT
  LAYER ME4 ;
  RECT 300.276 1.781 300.616 293.175 ;
 END
 PORT
  LAYER ME4 ;
  RECT 301.087 0.000 301.807 44.094 ;
 END
 PORT
  LAYER ME4 ;
  RECT 306.282 1.781 306.622 293.175 ;
 END
 PORT
  LAYER ME4 ;
  RECT 304.280 1.781 304.620 293.175 ;
 END
 PORT
  LAYER ME4 ;
  RECT 305.091 0.000 305.811 44.094 ;
 END
 PORT
  LAYER ME4 ;
  RECT 310.286 1.781 310.626 293.175 ;
 END
 PORT
  LAYER ME4 ;
  RECT 308.284 1.781 308.624 293.175 ;
 END
 PORT
  LAYER ME4 ;
  RECT 309.095 0.000 309.815 44.094 ;
 END
 PORT
  LAYER ME4 ;
  RECT 314.290 1.781 314.630 293.175 ;
 END
 PORT
  LAYER ME4 ;
  RECT 312.288 1.781 312.628 293.175 ;
 END
 PORT
  LAYER ME4 ;
  RECT 313.099 0.000 313.819 44.094 ;
 END
 PORT
  LAYER ME4 ;
  RECT 318.294 1.781 318.634 293.175 ;
 END
 PORT
  LAYER ME4 ;
  RECT 316.292 1.781 316.632 293.175 ;
 END
 PORT
  LAYER ME4 ;
  RECT 317.103 0.000 317.823 44.094 ;
 END
 PORT
  LAYER ME4 ;
  RECT 322.298 1.781 322.638 293.175 ;
 END
 PORT
  LAYER ME4 ;
  RECT 320.296 1.781 320.636 293.175 ;
 END
 PORT
  LAYER ME4 ;
  RECT 321.107 0.000 321.827 44.094 ;
 END
 PORT
  LAYER ME4 ;
  RECT 326.302 1.781 326.642 293.175 ;
 END
 PORT
  LAYER ME4 ;
  RECT 324.300 1.781 324.640 293.175 ;
 END
 PORT
  LAYER ME4 ;
  RECT 325.111 0.000 325.831 44.094 ;
 END
 PORT
  LAYER ME4 ;
  RECT 330.306 1.781 330.646 293.175 ;
 END
 PORT
  LAYER ME4 ;
  RECT 328.304 1.781 328.644 293.175 ;
 END
 PORT
  LAYER ME4 ;
  RECT 329.115 0.000 329.835 44.094 ;
 END
 PORT
  LAYER ME4 ;
  RECT 334.310 1.781 334.650 293.175 ;
 END
 PORT
  LAYER ME4 ;
  RECT 332.308 1.781 332.648 293.175 ;
 END
 PORT
  LAYER ME4 ;
  RECT 333.119 0.000 333.839 44.094 ;
 END
 PORT
  LAYER ME4 ;
  RECT 338.314 1.781 338.654 293.175 ;
 END
 PORT
  LAYER ME4 ;
  RECT 336.312 1.781 336.652 293.175 ;
 END
 PORT
  LAYER ME4 ;
  RECT 337.123 0.000 337.843 44.094 ;
 END
 PORT
  LAYER ME4 ;
  RECT 342.318 1.781 342.658 293.175 ;
 END
 PORT
  LAYER ME4 ;
  RECT 340.316 1.781 340.656 293.175 ;
 END
 PORT
  LAYER ME4 ;
  RECT 341.127 0.000 341.847 44.094 ;
 END
 PORT
  LAYER ME4 ;
  RECT 346.322 1.781 346.662 293.175 ;
 END
 PORT
  LAYER ME4 ;
  RECT 344.320 1.781 344.660 293.175 ;
 END
 PORT
  LAYER ME4 ;
  RECT 345.131 0.000 345.851 44.094 ;
 END
 PORT
  LAYER ME4 ;
  RECT 350.326 1.781 350.666 293.175 ;
 END
 PORT
  LAYER ME4 ;
  RECT 348.324 1.781 348.664 293.175 ;
 END
 PORT
  LAYER ME4 ;
  RECT 349.135 0.000 349.855 44.094 ;
 END
 PORT
  LAYER ME4 ;
  RECT 354.330 1.781 354.670 293.175 ;
 END
 PORT
  LAYER ME4 ;
  RECT 352.328 1.781 352.668 293.175 ;
 END
 PORT
  LAYER ME4 ;
  RECT 353.139 0.000 353.859 44.094 ;
 END
 PORT
  LAYER ME4 ;
  RECT 358.334 1.781 358.674 293.175 ;
 END
 PORT
  LAYER ME4 ;
  RECT 356.332 1.781 356.672 293.175 ;
 END
 PORT
  LAYER ME4 ;
  RECT 357.143 0.000 357.863 44.094 ;
 END
 PORT
  LAYER ME4 ;
  RECT 362.338 1.781 362.678 293.175 ;
 END
 PORT
  LAYER ME4 ;
  RECT 360.336 1.781 360.676 293.175 ;
 END
 PORT
  LAYER ME4 ;
  RECT 361.147 0.000 361.867 44.094 ;
 END
 PORT
  LAYER ME4 ;
  RECT 366.342 1.781 366.682 293.175 ;
 END
 PORT
  LAYER ME4 ;
  RECT 364.340 1.781 364.680 293.175 ;
 END
 PORT
  LAYER ME4 ;
  RECT 365.151 0.000 365.871 44.094 ;
 END
 PORT
  LAYER ME4 ;
  RECT 370.346 1.781 370.686 293.175 ;
 END
 PORT
  LAYER ME4 ;
  RECT 368.344 1.781 368.684 293.175 ;
 END
 PORT
  LAYER ME4 ;
  RECT 369.155 0.000 369.875 44.094 ;
 END
 PORT
  LAYER ME4 ;
  RECT 374.350 1.781 374.690 293.175 ;
 END
 PORT
  LAYER ME4 ;
  RECT 372.348 1.781 372.688 293.175 ;
 END
 PORT
  LAYER ME4 ;
  RECT 373.159 0.000 373.879 44.094 ;
 END
 PORT
  LAYER ME4 ;
  RECT 378.354 1.781 378.694 293.175 ;
 END
 PORT
  LAYER ME4 ;
  RECT 376.352 1.781 376.692 293.175 ;
 END
 PORT
  LAYER ME4 ;
  RECT 377.163 0.000 377.883 44.094 ;
 END
 PORT
  LAYER ME4 ;
  RECT 382.358 1.781 382.698 293.175 ;
 END
 PORT
  LAYER ME4 ;
  RECT 380.356 1.781 380.696 293.175 ;
 END
 PORT
  LAYER ME4 ;
  RECT 381.167 0.000 381.887 44.094 ;
 END
 PORT
  LAYER ME4 ;
  RECT 386.362 1.781 386.702 293.175 ;
 END
 PORT
  LAYER ME4 ;
  RECT 384.360 1.781 384.700 293.175 ;
 END
 PORT
  LAYER ME4 ;
  RECT 385.171 0.000 385.891 44.094 ;
 END
 PORT
  LAYER ME4 ;
  RECT 390.366 1.781 390.706 293.175 ;
 END
 PORT
  LAYER ME4 ;
  RECT 388.364 1.781 388.704 293.175 ;
 END
 PORT
  LAYER ME4 ;
  RECT 389.175 0.000 389.895 44.094 ;
 END
 PORT
  LAYER ME4 ;
  RECT 394.370 1.781 394.710 293.175 ;
 END
 PORT
  LAYER ME4 ;
  RECT 392.368 1.781 392.708 293.175 ;
 END
 PORT
  LAYER ME4 ;
  RECT 393.179 0.000 393.899 44.094 ;
 END
 PORT
  LAYER ME4 ;
  RECT 398.374 1.781 398.714 293.175 ;
 END
 PORT
  LAYER ME4 ;
  RECT 396.372 1.781 396.712 293.175 ;
 END
 PORT
  LAYER ME4 ;
  RECT 397.183 0.000 397.903 44.094 ;
 END
 PORT
  LAYER ME4 ;
  RECT 402.378 1.781 402.718 293.175 ;
 END
 PORT
  LAYER ME4 ;
  RECT 400.376 1.781 400.716 293.175 ;
 END
 PORT
  LAYER ME4 ;
  RECT 401.187 0.000 401.907 44.094 ;
 END
 PORT
  LAYER ME4 ;
  RECT 406.382 1.781 406.722 293.175 ;
 END
 PORT
  LAYER ME4 ;
  RECT 404.380 1.781 404.720 293.175 ;
 END
 PORT
  LAYER ME4 ;
  RECT 405.191 0.000 405.911 44.094 ;
 END
 PORT
  LAYER ME4 ;
  RECT 410.386 1.781 410.726 293.175 ;
 END
 PORT
  LAYER ME4 ;
  RECT 408.384 1.781 408.724 293.175 ;
 END
 PORT
  LAYER ME4 ;
  RECT 409.195 0.000 409.915 44.094 ;
 END
 PORT
  LAYER ME4 ;
  RECT 414.390 1.781 414.730 293.175 ;
 END
 PORT
  LAYER ME4 ;
  RECT 412.388 1.781 412.728 293.175 ;
 END
 PORT
  LAYER ME4 ;
  RECT 413.199 0.000 413.919 44.094 ;
 END
 PORT
  LAYER ME4 ;
  RECT 418.394 1.781 418.734 293.175 ;
 END
 PORT
  LAYER ME4 ;
  RECT 416.392 1.781 416.732 293.175 ;
 END
 PORT
  LAYER ME4 ;
  RECT 417.203 0.000 417.923 44.094 ;
 END
 PORT
  LAYER ME4 ;
  RECT 422.398 1.781 422.738 293.175 ;
 END
 PORT
  LAYER ME4 ;
  RECT 420.396 1.781 420.736 293.175 ;
 END
 PORT
  LAYER ME4 ;
  RECT 421.207 0.000 421.927 44.094 ;
 END
 PORT
  LAYER ME4 ;
  RECT 426.402 1.781 426.742 293.175 ;
 END
 PORT
  LAYER ME4 ;
  RECT 424.400 1.781 424.740 293.175 ;
 END
 PORT
  LAYER ME4 ;
  RECT 425.211 0.000 425.931 44.094 ;
 END
 PORT
  LAYER ME4 ;
  RECT 430.406 1.781 430.746 293.175 ;
 END
 PORT
  LAYER ME4 ;
  RECT 428.404 1.781 428.744 293.175 ;
 END
 PORT
  LAYER ME4 ;
  RECT 429.215 0.000 429.935 44.094 ;
 END
 PORT
  LAYER ME4 ;
  RECT 434.410 1.781 434.750 293.175 ;
 END
 PORT
  LAYER ME4 ;
  RECT 432.408 1.781 432.748 293.175 ;
 END
 PORT
  LAYER ME4 ;
  RECT 433.219 0.000 433.939 44.094 ;
 END
 PORT
  LAYER ME4 ;
  RECT 438.414 1.781 438.754 293.175 ;
 END
 PORT
  LAYER ME4 ;
  RECT 436.412 1.781 436.752 293.175 ;
 END
 PORT
  LAYER ME4 ;
  RECT 437.223 0.000 437.943 44.094 ;
 END
 PORT
  LAYER ME4 ;
  RECT 442.418 1.781 442.758 293.175 ;
 END
 PORT
  LAYER ME4 ;
  RECT 440.416 1.781 440.756 293.175 ;
 END
 PORT
  LAYER ME4 ;
  RECT 441.227 0.000 441.947 44.094 ;
 END
 PORT
  LAYER ME4 ;
  RECT 446.422 1.781 446.762 293.175 ;
 END
 PORT
  LAYER ME4 ;
  RECT 444.420 1.781 444.760 293.175 ;
 END
 PORT
  LAYER ME4 ;
  RECT 445.231 0.000 445.951 44.094 ;
 END
 PORT
  LAYER ME4 ;
  RECT 450.426 1.781 450.766 293.175 ;
 END
 PORT
  LAYER ME4 ;
  RECT 448.424 1.781 448.764 293.175 ;
 END
 PORT
  LAYER ME4 ;
  RECT 449.235 0.000 449.955 44.094 ;
 END
 PORT
  LAYER ME4 ;
  RECT 454.430 1.781 454.770 293.175 ;
 END
 PORT
  LAYER ME4 ;
  RECT 452.428 1.781 452.768 293.175 ;
 END
 PORT
  LAYER ME4 ;
  RECT 453.239 0.000 453.959 44.094 ;
 END
 PORT
  LAYER ME4 ;
  RECT 458.434 1.781 458.774 293.175 ;
 END
 PORT
  LAYER ME4 ;
  RECT 456.432 1.781 456.772 293.175 ;
 END
 PORT
  LAYER ME4 ;
  RECT 457.243 0.000 457.963 44.094 ;
 END
 PORT
  LAYER ME4 ;
  RECT 462.438 1.781 462.778 293.175 ;
 END
 PORT
  LAYER ME4 ;
  RECT 460.436 1.781 460.776 293.175 ;
 END
 PORT
  LAYER ME4 ;
  RECT 461.247 0.000 461.967 44.094 ;
 END
 PORT
  LAYER ME4 ;
  RECT 466.442 1.781 466.782 293.175 ;
 END
 PORT
  LAYER ME4 ;
  RECT 464.440 1.781 464.780 293.175 ;
 END
 PORT
  LAYER ME4 ;
  RECT 465.251 0.000 465.971 44.094 ;
 END
 PORT
  LAYER ME4 ;
  RECT 470.446 1.781 470.786 293.175 ;
 END
 PORT
  LAYER ME4 ;
  RECT 468.444 1.781 468.784 293.175 ;
 END
 PORT
  LAYER ME4 ;
  RECT 469.255 0.000 469.975 44.094 ;
 END
 PORT
  LAYER ME4 ;
  RECT 474.450 1.781 474.790 293.175 ;
 END
 PORT
  LAYER ME4 ;
  RECT 472.448 1.781 472.788 293.175 ;
 END
 PORT
  LAYER ME4 ;
  RECT 473.259 0.000 473.979 44.094 ;
 END
 PORT
  LAYER ME4 ;
  RECT 478.454 1.781 478.794 293.175 ;
 END
 PORT
  LAYER ME4 ;
  RECT 476.452 1.781 476.792 293.175 ;
 END
 PORT
  LAYER ME4 ;
  RECT 477.263 0.000 477.983 44.094 ;
 END
 PORT
  LAYER ME4 ;
  RECT 482.458 1.781 482.798 293.175 ;
 END
 PORT
  LAYER ME4 ;
  RECT 480.456 1.781 480.796 293.175 ;
 END
 PORT
  LAYER ME4 ;
  RECT 481.267 0.000 481.987 44.094 ;
 END
 PORT
  LAYER ME4 ;
  RECT 486.462 1.781 486.802 293.175 ;
 END
 PORT
  LAYER ME4 ;
  RECT 484.460 1.781 484.800 293.175 ;
 END
 PORT
  LAYER ME4 ;
  RECT 485.271 0.000 485.991 44.094 ;
 END
 PORT
  LAYER ME4 ;
  RECT 490.466 1.781 490.806 293.175 ;
 END
 PORT
  LAYER ME4 ;
  RECT 488.464 1.781 488.804 293.175 ;
 END
 PORT
  LAYER ME4 ;
  RECT 489.275 0.000 489.995 44.094 ;
 END
 PORT
  LAYER ME4 ;
  RECT 494.470 1.781 494.810 293.175 ;
 END
 PORT
  LAYER ME4 ;
  RECT 492.468 1.781 492.808 293.175 ;
 END
 PORT
  LAYER ME4 ;
  RECT 493.279 0.000 493.999 44.094 ;
 END
 PORT
  LAYER ME4 ;
  RECT 498.474 1.781 498.814 293.175 ;
 END
 PORT
  LAYER ME4 ;
  RECT 496.472 1.781 496.812 293.175 ;
 END
 PORT
  LAYER ME4 ;
  RECT 497.283 0.000 498.003 44.094 ;
 END
 PORT
  LAYER ME4 ;
  RECT 502.478 1.781 502.818 293.175 ;
 END
 PORT
  LAYER ME4 ;
  RECT 500.476 1.781 500.816 293.175 ;
 END
 PORT
  LAYER ME4 ;
  RECT 501.287 0.000 502.007 44.094 ;
 END
 PORT
  LAYER ME4 ;
  RECT 506.482 1.781 506.822 293.175 ;
 END
 PORT
  LAYER ME4 ;
  RECT 504.480 1.781 504.820 293.175 ;
 END
 PORT
  LAYER ME4 ;
  RECT 505.291 0.000 506.011 44.094 ;
 END
 PORT
  LAYER ME4 ;
  RECT 510.486 1.781 510.826 293.175 ;
 END
 PORT
  LAYER ME4 ;
  RECT 508.484 1.781 508.824 293.175 ;
 END
 PORT
  LAYER ME4 ;
  RECT 509.295 0.000 510.015 44.094 ;
 END
 PORT
  LAYER ME4 ;
  RECT 514.490 1.781 514.830 293.175 ;
 END
 PORT
  LAYER ME4 ;
  RECT 512.488 1.781 512.828 293.175 ;
 END
 PORT
  LAYER ME4 ;
  RECT 513.299 0.000 514.019 44.094 ;
 END
 PORT
  LAYER ME4 ;
  RECT 518.494 1.781 518.834 293.175 ;
 END
 PORT
  LAYER ME4 ;
  RECT 516.492 1.781 516.832 293.175 ;
 END
 PORT
  LAYER ME4 ;
  RECT 517.303 0.000 518.023 44.094 ;
 END
 PORT
  LAYER ME4 ;
  RECT 522.498 1.781 522.838 293.175 ;
 END
 PORT
  LAYER ME4 ;
  RECT 520.496 1.781 520.836 293.175 ;
 END
 PORT
  LAYER ME4 ;
  RECT 521.307 0.000 522.027 44.094 ;
 END
 PORT
  LAYER ME4 ;
  RECT 526.502 1.781 526.842 293.175 ;
 END
 PORT
  LAYER ME4 ;
  RECT 524.500 1.781 524.840 293.175 ;
 END
 PORT
  LAYER ME4 ;
  RECT 525.311 0.000 526.031 44.094 ;
 END
 PORT
  LAYER ME4 ;
  RECT 530.506 1.781 530.846 293.175 ;
 END
 PORT
  LAYER ME4 ;
  RECT 528.504 1.781 528.844 293.175 ;
 END
 PORT
  LAYER ME4 ;
  RECT 529.315 0.000 530.035 44.094 ;
 END
 PORT
  LAYER ME4 ;
  RECT 534.510 1.781 534.850 293.175 ;
 END
 PORT
  LAYER ME4 ;
  RECT 532.508 1.781 532.848 293.175 ;
 END
 PORT
  LAYER ME4 ;
  RECT 533.319 0.000 534.039 44.094 ;
 END
 PORT
  LAYER ME4 ;
  RECT 538.514 1.781 538.854 293.175 ;
 END
 PORT
  LAYER ME4 ;
  RECT 536.512 1.781 536.852 293.175 ;
 END
 PORT
  LAYER ME4 ;
  RECT 537.323 0.000 538.043 44.094 ;
 END
 PORT
  LAYER ME4 ;
  RECT 542.518 1.781 542.858 293.175 ;
 END
 PORT
  LAYER ME4 ;
  RECT 540.516 1.781 540.856 293.175 ;
 END
 PORT
  LAYER ME4 ;
  RECT 541.327 0.000 542.047 44.094 ;
 END
 PORT
  LAYER ME4 ;
  RECT 546.522 1.781 546.862 293.175 ;
 END
 PORT
  LAYER ME4 ;
  RECT 544.520 1.781 544.860 293.175 ;
 END
 PORT
  LAYER ME4 ;
  RECT 545.331 0.000 546.051 44.094 ;
 END
 PORT
  LAYER ME4 ;
  RECT 550.526 1.781 550.866 293.175 ;
 END
 PORT
  LAYER ME4 ;
  RECT 548.524 1.781 548.864 293.175 ;
 END
 PORT
  LAYER ME4 ;
  RECT 549.335 0.000 550.055 44.094 ;
 END
 PORT
  LAYER ME4 ;
  RECT 554.530 1.781 554.870 293.175 ;
 END
 PORT
  LAYER ME4 ;
  RECT 552.528 1.781 552.868 293.175 ;
 END
 PORT
  LAYER ME4 ;
  RECT 553.339 0.000 554.059 44.094 ;
 END
 PORT
  LAYER ME4 ;
  RECT 555.531 0.000 555.871 293.175 ;
 END
 PORT
  LAYER ME4 ;
  RECT 279.417 0.000 280.137 293.175 ;
 END
 PORT
  LAYER ME4 ;
  RECT 285.411 0.000 286.131 293.175 ;
 END
 PORT
  LAYER ME4 ;
  RECT 290.882 0.000 291.602 293.175 ;
 END
 PORT
  LAYER ME4 ;
  RECT 292.597 0.000 293.317 293.175 ;
 END
 PORT
  LAYER ME4 ;
  RECT 295.593 0.000 296.193 293.175 ;
 END
 PORT
  LAYER ME4 ;
  RECT 297.273 1.781 297.613 293.175 ;
 END
 PORT
  LAYER ME4 ;
  RECT 271.858 0.000 272.578 293.175 ;
 END
 PORT
  LAYER ME4 ;
  RECT 269.818 1.781 270.538 292.295 ;
 END
 PORT
  LAYER ME4 ;
  RECT 267.698 0.000 268.418 293.175 ;
 END
 PORT
  LAYER ME4 ;
  RECT 265.658 1.781 266.378 293.175 ;
 END
 PORT
  LAYER ME4 ;
  RECT 263.538 0.000 264.258 293.175 ;
 END
 PORT
  LAYER ME4 ;
  RECT 261.498 1.781 262.218 293.175 ;
 END
 PORT
  LAYER ME4 ;
  RECT 1.740 0.000 2.080 293.175 ;
 END
 PORT
  LAYER ME4 ;
  RECT 6.745 1.781 7.085 293.175 ;
 END
 PORT
  LAYER ME4 ;
  RECT 2.741 1.781 3.081 293.175 ;
 END
 PORT
  LAYER ME4 ;
  RECT 4.743 1.781 5.083 293.175 ;
 END
 PORT
  LAYER ME4 ;
  RECT 5.554 0.000 6.274 44.094 ;
 END
 PORT
  LAYER ME4 ;
  RECT 10.749 1.781 11.089 293.175 ;
 END
 PORT
  LAYER ME4 ;
  RECT 8.747 1.781 9.087 293.175 ;
 END
 PORT
  LAYER ME4 ;
  RECT 9.558 0.000 10.278 44.094 ;
 END
 PORT
  LAYER ME4 ;
  RECT 14.753 1.781 15.093 293.175 ;
 END
 PORT
  LAYER ME4 ;
  RECT 12.751 1.781 13.091 293.175 ;
 END
 PORT
  LAYER ME4 ;
  RECT 13.562 0.000 14.282 44.094 ;
 END
 PORT
  LAYER ME4 ;
  RECT 18.757 1.781 19.097 293.175 ;
 END
 PORT
  LAYER ME4 ;
  RECT 16.755 1.781 17.095 293.175 ;
 END
 PORT
  LAYER ME4 ;
  RECT 17.566 0.000 18.286 44.094 ;
 END
 PORT
  LAYER ME4 ;
  RECT 22.761 1.781 23.101 293.175 ;
 END
 PORT
  LAYER ME4 ;
  RECT 20.759 1.781 21.099 293.175 ;
 END
 PORT
  LAYER ME4 ;
  RECT 21.570 0.000 22.290 44.094 ;
 END
 PORT
  LAYER ME4 ;
  RECT 26.765 1.781 27.105 293.175 ;
 END
 PORT
  LAYER ME4 ;
  RECT 24.763 1.781 25.103 293.175 ;
 END
 PORT
  LAYER ME4 ;
  RECT 25.574 0.000 26.294 44.094 ;
 END
 PORT
  LAYER ME4 ;
  RECT 30.769 1.781 31.109 293.175 ;
 END
 PORT
  LAYER ME4 ;
  RECT 28.767 1.781 29.107 293.175 ;
 END
 PORT
  LAYER ME4 ;
  RECT 29.578 0.000 30.298 44.094 ;
 END
 PORT
  LAYER ME4 ;
  RECT 34.773 1.781 35.113 293.175 ;
 END
 PORT
  LAYER ME4 ;
  RECT 32.771 1.781 33.111 293.175 ;
 END
 PORT
  LAYER ME4 ;
  RECT 33.582 0.000 34.302 44.094 ;
 END
 PORT
  LAYER ME4 ;
  RECT 38.777 1.781 39.117 293.175 ;
 END
 PORT
  LAYER ME4 ;
  RECT 36.775 1.781 37.115 293.175 ;
 END
 PORT
  LAYER ME4 ;
  RECT 37.586 0.000 38.306 44.094 ;
 END
 PORT
  LAYER ME4 ;
  RECT 42.781 1.781 43.121 293.175 ;
 END
 PORT
  LAYER ME4 ;
  RECT 40.779 1.781 41.119 293.175 ;
 END
 PORT
  LAYER ME4 ;
  RECT 41.590 0.000 42.310 44.094 ;
 END
 PORT
  LAYER ME4 ;
  RECT 46.785 1.781 47.125 293.175 ;
 END
 PORT
  LAYER ME4 ;
  RECT 44.783 1.781 45.123 293.175 ;
 END
 PORT
  LAYER ME4 ;
  RECT 45.594 0.000 46.314 44.094 ;
 END
 PORT
  LAYER ME4 ;
  RECT 50.789 1.781 51.129 293.175 ;
 END
 PORT
  LAYER ME4 ;
  RECT 48.787 1.781 49.127 293.175 ;
 END
 PORT
  LAYER ME4 ;
  RECT 49.598 0.000 50.318 44.094 ;
 END
 PORT
  LAYER ME4 ;
  RECT 54.793 1.781 55.133 293.175 ;
 END
 PORT
  LAYER ME4 ;
  RECT 52.791 1.781 53.131 293.175 ;
 END
 PORT
  LAYER ME4 ;
  RECT 53.602 0.000 54.322 44.094 ;
 END
 PORT
  LAYER ME4 ;
  RECT 58.797 1.781 59.137 293.175 ;
 END
 PORT
  LAYER ME4 ;
  RECT 56.795 1.781 57.135 293.175 ;
 END
 PORT
  LAYER ME4 ;
  RECT 57.606 0.000 58.326 44.094 ;
 END
 PORT
  LAYER ME4 ;
  RECT 62.801 1.781 63.141 293.175 ;
 END
 PORT
  LAYER ME4 ;
  RECT 60.799 1.781 61.139 293.175 ;
 END
 PORT
  LAYER ME4 ;
  RECT 61.610 0.000 62.330 44.094 ;
 END
 PORT
  LAYER ME4 ;
  RECT 66.805 1.781 67.145 293.175 ;
 END
 PORT
  LAYER ME4 ;
  RECT 64.803 1.781 65.143 293.175 ;
 END
 PORT
  LAYER ME4 ;
  RECT 65.614 0.000 66.334 44.094 ;
 END
 PORT
  LAYER ME4 ;
  RECT 70.809 1.781 71.149 293.175 ;
 END
 PORT
  LAYER ME4 ;
  RECT 68.807 1.781 69.147 293.175 ;
 END
 PORT
  LAYER ME4 ;
  RECT 69.618 0.000 70.338 44.094 ;
 END
 PORT
  LAYER ME4 ;
  RECT 74.813 1.781 75.153 293.175 ;
 END
 PORT
  LAYER ME4 ;
  RECT 72.811 1.781 73.151 293.175 ;
 END
 PORT
  LAYER ME4 ;
  RECT 73.622 0.000 74.342 44.094 ;
 END
 PORT
  LAYER ME4 ;
  RECT 78.817 1.781 79.157 293.175 ;
 END
 PORT
  LAYER ME4 ;
  RECT 76.815 1.781 77.155 293.175 ;
 END
 PORT
  LAYER ME4 ;
  RECT 77.626 0.000 78.346 44.094 ;
 END
 PORT
  LAYER ME4 ;
  RECT 82.821 1.781 83.161 293.175 ;
 END
 PORT
  LAYER ME4 ;
  RECT 80.819 1.781 81.159 293.175 ;
 END
 PORT
  LAYER ME4 ;
  RECT 81.630 0.000 82.350 44.094 ;
 END
 PORT
  LAYER ME4 ;
  RECT 86.825 1.781 87.165 293.175 ;
 END
 PORT
  LAYER ME4 ;
  RECT 84.823 1.781 85.163 293.175 ;
 END
 PORT
  LAYER ME4 ;
  RECT 85.634 0.000 86.354 44.094 ;
 END
 PORT
  LAYER ME4 ;
  RECT 90.829 1.781 91.169 293.175 ;
 END
 PORT
  LAYER ME4 ;
  RECT 88.827 1.781 89.167 293.175 ;
 END
 PORT
  LAYER ME4 ;
  RECT 89.638 0.000 90.358 44.094 ;
 END
 PORT
  LAYER ME4 ;
  RECT 94.833 1.781 95.173 293.175 ;
 END
 PORT
  LAYER ME4 ;
  RECT 92.831 1.781 93.171 293.175 ;
 END
 PORT
  LAYER ME4 ;
  RECT 93.642 0.000 94.362 44.094 ;
 END
 PORT
  LAYER ME4 ;
  RECT 98.837 1.781 99.177 293.175 ;
 END
 PORT
  LAYER ME4 ;
  RECT 96.835 1.781 97.175 293.175 ;
 END
 PORT
  LAYER ME4 ;
  RECT 97.646 0.000 98.366 44.094 ;
 END
 PORT
  LAYER ME4 ;
  RECT 102.841 1.781 103.181 293.175 ;
 END
 PORT
  LAYER ME4 ;
  RECT 100.839 1.781 101.179 293.175 ;
 END
 PORT
  LAYER ME4 ;
  RECT 101.650 0.000 102.370 44.094 ;
 END
 PORT
  LAYER ME4 ;
  RECT 106.845 1.781 107.185 293.175 ;
 END
 PORT
  LAYER ME4 ;
  RECT 104.843 1.781 105.183 293.175 ;
 END
 PORT
  LAYER ME4 ;
  RECT 105.654 0.000 106.374 44.094 ;
 END
 PORT
  LAYER ME4 ;
  RECT 110.849 1.781 111.189 293.175 ;
 END
 PORT
  LAYER ME4 ;
  RECT 108.847 1.781 109.187 293.175 ;
 END
 PORT
  LAYER ME4 ;
  RECT 109.658 0.000 110.378 44.094 ;
 END
 PORT
  LAYER ME4 ;
  RECT 114.853 1.781 115.193 293.175 ;
 END
 PORT
  LAYER ME4 ;
  RECT 112.851 1.781 113.191 293.175 ;
 END
 PORT
  LAYER ME4 ;
  RECT 113.662 0.000 114.382 44.094 ;
 END
 PORT
  LAYER ME4 ;
  RECT 118.857 1.781 119.197 293.175 ;
 END
 PORT
  LAYER ME4 ;
  RECT 116.855 1.781 117.195 293.175 ;
 END
 PORT
  LAYER ME4 ;
  RECT 117.666 0.000 118.386 44.094 ;
 END
 PORT
  LAYER ME4 ;
  RECT 122.861 1.781 123.201 293.175 ;
 END
 PORT
  LAYER ME4 ;
  RECT 120.859 1.781 121.199 293.175 ;
 END
 PORT
  LAYER ME4 ;
  RECT 121.670 0.000 122.390 44.094 ;
 END
 PORT
  LAYER ME4 ;
  RECT 126.865 1.781 127.205 293.175 ;
 END
 PORT
  LAYER ME4 ;
  RECT 124.863 1.781 125.203 293.175 ;
 END
 PORT
  LAYER ME4 ;
  RECT 125.674 0.000 126.394 44.094 ;
 END
 PORT
  LAYER ME4 ;
  RECT 130.869 1.781 131.209 293.175 ;
 END
 PORT
  LAYER ME4 ;
  RECT 128.867 1.781 129.207 293.175 ;
 END
 PORT
  LAYER ME4 ;
  RECT 129.678 0.000 130.398 44.094 ;
 END
 PORT
  LAYER ME4 ;
  RECT 134.873 1.781 135.213 293.175 ;
 END
 PORT
  LAYER ME4 ;
  RECT 132.871 1.781 133.211 293.175 ;
 END
 PORT
  LAYER ME4 ;
  RECT 133.682 0.000 134.402 44.094 ;
 END
 PORT
  LAYER ME4 ;
  RECT 138.877 1.781 139.217 293.175 ;
 END
 PORT
  LAYER ME4 ;
  RECT 136.875 1.781 137.215 293.175 ;
 END
 PORT
  LAYER ME4 ;
  RECT 137.686 0.000 138.406 44.094 ;
 END
 PORT
  LAYER ME4 ;
  RECT 142.881 1.781 143.221 293.175 ;
 END
 PORT
  LAYER ME4 ;
  RECT 140.879 1.781 141.219 293.175 ;
 END
 PORT
  LAYER ME4 ;
  RECT 141.690 0.000 142.410 44.094 ;
 END
 PORT
  LAYER ME4 ;
  RECT 146.885 1.781 147.225 293.175 ;
 END
 PORT
  LAYER ME4 ;
  RECT 144.883 1.781 145.223 293.175 ;
 END
 PORT
  LAYER ME4 ;
  RECT 145.694 0.000 146.414 44.094 ;
 END
 PORT
  LAYER ME4 ;
  RECT 150.889 1.781 151.229 293.175 ;
 END
 PORT
  LAYER ME4 ;
  RECT 148.887 1.781 149.227 293.175 ;
 END
 PORT
  LAYER ME4 ;
  RECT 149.698 0.000 150.418 44.094 ;
 END
 PORT
  LAYER ME4 ;
  RECT 154.893 1.781 155.233 293.175 ;
 END
 PORT
  LAYER ME4 ;
  RECT 152.891 1.781 153.231 293.175 ;
 END
 PORT
  LAYER ME4 ;
  RECT 153.702 0.000 154.422 44.094 ;
 END
 PORT
  LAYER ME4 ;
  RECT 158.897 1.781 159.237 293.175 ;
 END
 PORT
  LAYER ME4 ;
  RECT 156.895 1.781 157.235 293.175 ;
 END
 PORT
  LAYER ME4 ;
  RECT 157.706 0.000 158.426 44.094 ;
 END
 PORT
  LAYER ME4 ;
  RECT 162.901 1.781 163.241 293.175 ;
 END
 PORT
  LAYER ME4 ;
  RECT 160.899 1.781 161.239 293.175 ;
 END
 PORT
  LAYER ME4 ;
  RECT 161.710 0.000 162.430 44.094 ;
 END
 PORT
  LAYER ME4 ;
  RECT 166.905 1.781 167.245 293.175 ;
 END
 PORT
  LAYER ME4 ;
  RECT 164.903 1.781 165.243 293.175 ;
 END
 PORT
  LAYER ME4 ;
  RECT 165.714 0.000 166.434 44.094 ;
 END
 PORT
  LAYER ME4 ;
  RECT 170.909 1.781 171.249 293.175 ;
 END
 PORT
  LAYER ME4 ;
  RECT 168.907 1.781 169.247 293.175 ;
 END
 PORT
  LAYER ME4 ;
  RECT 169.718 0.000 170.438 44.094 ;
 END
 PORT
  LAYER ME4 ;
  RECT 174.913 1.781 175.253 293.175 ;
 END
 PORT
  LAYER ME4 ;
  RECT 172.911 1.781 173.251 293.175 ;
 END
 PORT
  LAYER ME4 ;
  RECT 173.722 0.000 174.442 44.094 ;
 END
 PORT
  LAYER ME4 ;
  RECT 178.917 1.781 179.257 293.175 ;
 END
 PORT
  LAYER ME4 ;
  RECT 176.915 1.781 177.255 293.175 ;
 END
 PORT
  LAYER ME4 ;
  RECT 177.726 0.000 178.446 44.094 ;
 END
 PORT
  LAYER ME4 ;
  RECT 182.921 1.781 183.261 293.175 ;
 END
 PORT
  LAYER ME4 ;
  RECT 180.919 1.781 181.259 293.175 ;
 END
 PORT
  LAYER ME4 ;
  RECT 181.730 0.000 182.450 44.094 ;
 END
 PORT
  LAYER ME4 ;
  RECT 186.925 1.781 187.265 293.175 ;
 END
 PORT
  LAYER ME4 ;
  RECT 184.923 1.781 185.263 293.175 ;
 END
 PORT
  LAYER ME4 ;
  RECT 185.734 0.000 186.454 44.094 ;
 END
 PORT
  LAYER ME4 ;
  RECT 190.929 1.781 191.269 293.175 ;
 END
 PORT
  LAYER ME4 ;
  RECT 188.927 1.781 189.267 293.175 ;
 END
 PORT
  LAYER ME4 ;
  RECT 189.738 0.000 190.458 44.094 ;
 END
 PORT
  LAYER ME4 ;
  RECT 194.933 1.781 195.273 293.175 ;
 END
 PORT
  LAYER ME4 ;
  RECT 192.931 1.781 193.271 293.175 ;
 END
 PORT
  LAYER ME4 ;
  RECT 193.742 0.000 194.462 44.094 ;
 END
 PORT
  LAYER ME4 ;
  RECT 198.937 1.781 199.277 293.175 ;
 END
 PORT
  LAYER ME4 ;
  RECT 196.935 1.781 197.275 293.175 ;
 END
 PORT
  LAYER ME4 ;
  RECT 197.746 0.000 198.466 44.094 ;
 END
 PORT
  LAYER ME4 ;
  RECT 202.941 1.781 203.281 293.175 ;
 END
 PORT
  LAYER ME4 ;
  RECT 200.939 1.781 201.279 293.175 ;
 END
 PORT
  LAYER ME4 ;
  RECT 201.750 0.000 202.470 44.094 ;
 END
 PORT
  LAYER ME4 ;
  RECT 206.945 1.781 207.285 293.175 ;
 END
 PORT
  LAYER ME4 ;
  RECT 204.943 1.781 205.283 293.175 ;
 END
 PORT
  LAYER ME4 ;
  RECT 205.754 0.000 206.474 44.094 ;
 END
 PORT
  LAYER ME4 ;
  RECT 210.949 1.781 211.289 293.175 ;
 END
 PORT
  LAYER ME4 ;
  RECT 208.947 1.781 209.287 293.175 ;
 END
 PORT
  LAYER ME4 ;
  RECT 209.758 0.000 210.478 44.094 ;
 END
 PORT
  LAYER ME4 ;
  RECT 214.953 1.781 215.293 293.175 ;
 END
 PORT
  LAYER ME4 ;
  RECT 212.951 1.781 213.291 293.175 ;
 END
 PORT
  LAYER ME4 ;
  RECT 213.762 0.000 214.482 44.094 ;
 END
 PORT
  LAYER ME4 ;
  RECT 218.957 1.781 219.297 293.175 ;
 END
 PORT
  LAYER ME4 ;
  RECT 216.955 1.781 217.295 293.175 ;
 END
 PORT
  LAYER ME4 ;
  RECT 217.766 0.000 218.486 44.094 ;
 END
 PORT
  LAYER ME4 ;
  RECT 222.961 1.781 223.301 293.175 ;
 END
 PORT
  LAYER ME4 ;
  RECT 220.959 1.781 221.299 293.175 ;
 END
 PORT
  LAYER ME4 ;
  RECT 221.770 0.000 222.490 44.094 ;
 END
 PORT
  LAYER ME4 ;
  RECT 226.965 1.781 227.305 293.175 ;
 END
 PORT
  LAYER ME4 ;
  RECT 224.963 1.781 225.303 293.175 ;
 END
 PORT
  LAYER ME4 ;
  RECT 225.774 0.000 226.494 44.094 ;
 END
 PORT
  LAYER ME4 ;
  RECT 230.969 1.781 231.309 293.175 ;
 END
 PORT
  LAYER ME4 ;
  RECT 228.967 1.781 229.307 293.175 ;
 END
 PORT
  LAYER ME4 ;
  RECT 229.778 0.000 230.498 44.094 ;
 END
 PORT
  LAYER ME4 ;
  RECT 234.973 1.781 235.313 293.175 ;
 END
 PORT
  LAYER ME4 ;
  RECT 232.971 1.781 233.311 293.175 ;
 END
 PORT
  LAYER ME4 ;
  RECT 233.782 0.000 234.502 44.094 ;
 END
 PORT
  LAYER ME4 ;
  RECT 238.977 1.781 239.317 293.175 ;
 END
 PORT
  LAYER ME4 ;
  RECT 236.975 1.781 237.315 293.175 ;
 END
 PORT
  LAYER ME4 ;
  RECT 237.786 0.000 238.506 44.094 ;
 END
 PORT
  LAYER ME4 ;
  RECT 242.981 1.781 243.321 293.175 ;
 END
 PORT
  LAYER ME4 ;
  RECT 240.979 1.781 241.319 293.175 ;
 END
 PORT
  LAYER ME4 ;
  RECT 241.790 0.000 242.510 44.094 ;
 END
 PORT
  LAYER ME4 ;
  RECT 246.985 1.781 247.325 293.175 ;
 END
 PORT
  LAYER ME4 ;
  RECT 244.983 1.781 245.323 293.175 ;
 END
 PORT
  LAYER ME4 ;
  RECT 245.794 0.000 246.514 44.094 ;
 END
 PORT
  LAYER ME4 ;
  RECT 250.989 1.781 251.329 293.175 ;
 END
 PORT
  LAYER ME4 ;
  RECT 248.987 1.781 249.327 293.175 ;
 END
 PORT
  LAYER ME4 ;
  RECT 249.798 0.000 250.518 44.094 ;
 END
 PORT
  LAYER ME4 ;
  RECT 254.993 1.781 255.333 293.175 ;
 END
 PORT
  LAYER ME4 ;
  RECT 252.991 1.781 253.331 293.175 ;
 END
 PORT
  LAYER ME4 ;
  RECT 253.802 0.000 254.522 44.094 ;
 END
 PORT
  LAYER ME4 ;
  RECT 258.997 1.781 259.337 293.175 ;
 END
 PORT
  LAYER ME4 ;
  RECT 256.995 1.781 257.335 293.175 ;
 END
 PORT
  LAYER ME4 ;
  RECT 257.806 0.000 258.526 44.094 ;
 END
 PORT
  LAYER ME4 ;
  RECT 259.998 0.000 260.338 293.175 ;
 END
END GND
PIN VCC
  DIRECTION INOUT ;
  USE POWER ;
 PORT
  LAYER ME4 ;
  RECT 301.277 45.394 301.617 293.175 ;
 END
 PORT
  LAYER ME4 ;
  RECT 299.085 0.000 299.805 46.394 ;
 END
 PORT
  LAYER ME4 ;
  RECT 305.281 45.394 305.621 293.175 ;
 END
 PORT
  LAYER ME4 ;
  RECT 303.089 0.000 303.809 46.394 ;
 END
 PORT
  LAYER ME4 ;
  RECT 309.285 45.394 309.625 293.175 ;
 END
 PORT
  LAYER ME4 ;
  RECT 307.093 0.000 307.813 46.394 ;
 END
 PORT
  LAYER ME4 ;
  RECT 313.289 45.394 313.629 293.175 ;
 END
 PORT
  LAYER ME4 ;
  RECT 311.097 0.000 311.817 46.394 ;
 END
 PORT
  LAYER ME4 ;
  RECT 317.293 45.394 317.633 293.175 ;
 END
 PORT
  LAYER ME4 ;
  RECT 315.101 0.000 315.821 46.394 ;
 END
 PORT
  LAYER ME4 ;
  RECT 321.297 45.394 321.637 293.175 ;
 END
 PORT
  LAYER ME4 ;
  RECT 319.105 0.000 319.825 46.394 ;
 END
 PORT
  LAYER ME4 ;
  RECT 325.301 45.394 325.641 293.175 ;
 END
 PORT
  LAYER ME4 ;
  RECT 323.109 0.000 323.829 46.394 ;
 END
 PORT
  LAYER ME4 ;
  RECT 329.305 45.394 329.645 293.175 ;
 END
 PORT
  LAYER ME4 ;
  RECT 327.113 0.000 327.833 46.394 ;
 END
 PORT
  LAYER ME4 ;
  RECT 333.309 45.394 333.649 293.175 ;
 END
 PORT
  LAYER ME4 ;
  RECT 331.117 0.000 331.837 46.394 ;
 END
 PORT
  LAYER ME4 ;
  RECT 337.313 45.394 337.653 293.175 ;
 END
 PORT
  LAYER ME4 ;
  RECT 335.121 0.000 335.841 46.394 ;
 END
 PORT
  LAYER ME4 ;
  RECT 341.317 45.394 341.657 293.175 ;
 END
 PORT
  LAYER ME4 ;
  RECT 339.125 0.000 339.845 46.394 ;
 END
 PORT
  LAYER ME4 ;
  RECT 345.321 45.394 345.661 293.175 ;
 END
 PORT
  LAYER ME4 ;
  RECT 343.129 0.000 343.849 46.394 ;
 END
 PORT
  LAYER ME4 ;
  RECT 349.325 45.394 349.665 293.175 ;
 END
 PORT
  LAYER ME4 ;
  RECT 347.133 0.000 347.853 46.394 ;
 END
 PORT
  LAYER ME4 ;
  RECT 353.329 45.394 353.669 293.175 ;
 END
 PORT
  LAYER ME4 ;
  RECT 351.137 0.000 351.857 46.394 ;
 END
 PORT
  LAYER ME4 ;
  RECT 357.333 45.394 357.673 293.175 ;
 END
 PORT
  LAYER ME4 ;
  RECT 355.141 0.000 355.861 46.394 ;
 END
 PORT
  LAYER ME4 ;
  RECT 361.337 45.394 361.677 293.175 ;
 END
 PORT
  LAYER ME4 ;
  RECT 359.145 0.000 359.865 46.394 ;
 END
 PORT
  LAYER ME4 ;
  RECT 365.341 45.394 365.681 293.175 ;
 END
 PORT
  LAYER ME4 ;
  RECT 363.149 0.000 363.869 46.394 ;
 END
 PORT
  LAYER ME4 ;
  RECT 369.345 45.394 369.685 293.175 ;
 END
 PORT
  LAYER ME4 ;
  RECT 367.153 0.000 367.873 46.394 ;
 END
 PORT
  LAYER ME4 ;
  RECT 373.349 45.394 373.689 293.175 ;
 END
 PORT
  LAYER ME4 ;
  RECT 371.157 0.000 371.877 46.394 ;
 END
 PORT
  LAYER ME4 ;
  RECT 377.353 45.394 377.693 293.175 ;
 END
 PORT
  LAYER ME4 ;
  RECT 375.161 0.000 375.881 46.394 ;
 END
 PORT
  LAYER ME4 ;
  RECT 381.357 45.394 381.697 293.175 ;
 END
 PORT
  LAYER ME4 ;
  RECT 379.165 0.000 379.885 46.394 ;
 END
 PORT
  LAYER ME4 ;
  RECT 385.361 45.394 385.701 293.175 ;
 END
 PORT
  LAYER ME4 ;
  RECT 383.169 0.000 383.889 46.394 ;
 END
 PORT
  LAYER ME4 ;
  RECT 389.365 45.394 389.705 293.175 ;
 END
 PORT
  LAYER ME4 ;
  RECT 387.173 0.000 387.893 46.394 ;
 END
 PORT
  LAYER ME4 ;
  RECT 393.369 45.394 393.709 293.175 ;
 END
 PORT
  LAYER ME4 ;
  RECT 391.177 0.000 391.897 46.394 ;
 END
 PORT
  LAYER ME4 ;
  RECT 397.373 45.394 397.713 293.175 ;
 END
 PORT
  LAYER ME4 ;
  RECT 395.181 0.000 395.901 46.394 ;
 END
 PORT
  LAYER ME4 ;
  RECT 401.377 45.394 401.717 293.175 ;
 END
 PORT
  LAYER ME4 ;
  RECT 399.185 0.000 399.905 46.394 ;
 END
 PORT
  LAYER ME4 ;
  RECT 405.381 45.394 405.721 293.175 ;
 END
 PORT
  LAYER ME4 ;
  RECT 403.189 0.000 403.909 46.394 ;
 END
 PORT
  LAYER ME4 ;
  RECT 409.385 45.394 409.725 293.175 ;
 END
 PORT
  LAYER ME4 ;
  RECT 407.193 0.000 407.913 46.394 ;
 END
 PORT
  LAYER ME4 ;
  RECT 413.389 45.394 413.729 293.175 ;
 END
 PORT
  LAYER ME4 ;
  RECT 411.197 0.000 411.917 46.394 ;
 END
 PORT
  LAYER ME4 ;
  RECT 417.393 45.394 417.733 293.175 ;
 END
 PORT
  LAYER ME4 ;
  RECT 415.201 0.000 415.921 46.394 ;
 END
 PORT
  LAYER ME4 ;
  RECT 421.397 45.394 421.737 293.175 ;
 END
 PORT
  LAYER ME4 ;
  RECT 419.205 0.000 419.925 46.394 ;
 END
 PORT
  LAYER ME4 ;
  RECT 425.401 45.394 425.741 293.175 ;
 END
 PORT
  LAYER ME4 ;
  RECT 423.209 0.000 423.929 46.394 ;
 END
 PORT
  LAYER ME4 ;
  RECT 429.405 45.394 429.745 293.175 ;
 END
 PORT
  LAYER ME4 ;
  RECT 427.213 0.000 427.933 46.394 ;
 END
 PORT
  LAYER ME4 ;
  RECT 433.409 45.394 433.749 293.175 ;
 END
 PORT
  LAYER ME4 ;
  RECT 431.217 0.000 431.937 46.394 ;
 END
 PORT
  LAYER ME4 ;
  RECT 437.413 45.394 437.753 293.175 ;
 END
 PORT
  LAYER ME4 ;
  RECT 435.221 0.000 435.941 46.394 ;
 END
 PORT
  LAYER ME4 ;
  RECT 441.417 45.394 441.757 293.175 ;
 END
 PORT
  LAYER ME4 ;
  RECT 439.225 0.000 439.945 46.394 ;
 END
 PORT
  LAYER ME4 ;
  RECT 445.421 45.394 445.761 293.175 ;
 END
 PORT
  LAYER ME4 ;
  RECT 443.229 0.000 443.949 46.394 ;
 END
 PORT
  LAYER ME4 ;
  RECT 449.425 45.394 449.765 293.175 ;
 END
 PORT
  LAYER ME4 ;
  RECT 447.233 0.000 447.953 46.394 ;
 END
 PORT
  LAYER ME4 ;
  RECT 453.429 45.394 453.769 293.175 ;
 END
 PORT
  LAYER ME4 ;
  RECT 451.237 0.000 451.957 46.394 ;
 END
 PORT
  LAYER ME4 ;
  RECT 457.433 45.394 457.773 293.175 ;
 END
 PORT
  LAYER ME4 ;
  RECT 455.241 0.000 455.961 46.394 ;
 END
 PORT
  LAYER ME4 ;
  RECT 461.437 45.394 461.777 293.175 ;
 END
 PORT
  LAYER ME4 ;
  RECT 459.245 0.000 459.965 46.394 ;
 END
 PORT
  LAYER ME4 ;
  RECT 465.441 45.394 465.781 293.175 ;
 END
 PORT
  LAYER ME4 ;
  RECT 463.249 0.000 463.969 46.394 ;
 END
 PORT
  LAYER ME4 ;
  RECT 469.445 45.394 469.785 293.175 ;
 END
 PORT
  LAYER ME4 ;
  RECT 467.253 0.000 467.973 46.394 ;
 END
 PORT
  LAYER ME4 ;
  RECT 473.449 45.394 473.789 293.175 ;
 END
 PORT
  LAYER ME4 ;
  RECT 471.257 0.000 471.977 46.394 ;
 END
 PORT
  LAYER ME4 ;
  RECT 477.453 45.394 477.793 293.175 ;
 END
 PORT
  LAYER ME4 ;
  RECT 475.261 0.000 475.981 46.394 ;
 END
 PORT
  LAYER ME4 ;
  RECT 481.457 45.394 481.797 293.175 ;
 END
 PORT
  LAYER ME4 ;
  RECT 479.265 0.000 479.985 46.394 ;
 END
 PORT
  LAYER ME4 ;
  RECT 485.461 45.394 485.801 293.175 ;
 END
 PORT
  LAYER ME4 ;
  RECT 483.269 0.000 483.989 46.394 ;
 END
 PORT
  LAYER ME4 ;
  RECT 489.465 45.394 489.805 293.175 ;
 END
 PORT
  LAYER ME4 ;
  RECT 487.273 0.000 487.993 46.394 ;
 END
 PORT
  LAYER ME4 ;
  RECT 493.469 45.394 493.809 293.175 ;
 END
 PORT
  LAYER ME4 ;
  RECT 491.277 0.000 491.997 46.394 ;
 END
 PORT
  LAYER ME4 ;
  RECT 497.473 45.394 497.813 293.175 ;
 END
 PORT
  LAYER ME4 ;
  RECT 495.281 0.000 496.001 46.394 ;
 END
 PORT
  LAYER ME4 ;
  RECT 501.477 45.394 501.817 293.175 ;
 END
 PORT
  LAYER ME4 ;
  RECT 499.285 0.000 500.005 46.394 ;
 END
 PORT
  LAYER ME4 ;
  RECT 505.481 45.394 505.821 293.175 ;
 END
 PORT
  LAYER ME4 ;
  RECT 503.289 0.000 504.009 46.394 ;
 END
 PORT
  LAYER ME4 ;
  RECT 509.485 45.394 509.825 293.175 ;
 END
 PORT
  LAYER ME4 ;
  RECT 507.293 0.000 508.013 46.394 ;
 END
 PORT
  LAYER ME4 ;
  RECT 513.489 45.394 513.829 293.175 ;
 END
 PORT
  LAYER ME4 ;
  RECT 511.297 0.000 512.017 46.394 ;
 END
 PORT
  LAYER ME4 ;
  RECT 517.493 45.394 517.833 293.175 ;
 END
 PORT
  LAYER ME4 ;
  RECT 515.301 0.000 516.021 46.394 ;
 END
 PORT
  LAYER ME4 ;
  RECT 521.497 45.394 521.837 293.175 ;
 END
 PORT
  LAYER ME4 ;
  RECT 519.305 0.000 520.025 46.394 ;
 END
 PORT
  LAYER ME4 ;
  RECT 525.501 45.394 525.841 293.175 ;
 END
 PORT
  LAYER ME4 ;
  RECT 523.309 0.000 524.029 46.394 ;
 END
 PORT
  LAYER ME4 ;
  RECT 529.505 45.394 529.845 293.175 ;
 END
 PORT
  LAYER ME4 ;
  RECT 527.313 0.000 528.033 46.394 ;
 END
 PORT
  LAYER ME4 ;
  RECT 533.509 45.394 533.849 293.175 ;
 END
 PORT
  LAYER ME4 ;
  RECT 531.317 0.000 532.037 46.394 ;
 END
 PORT
  LAYER ME4 ;
  RECT 537.513 45.394 537.853 293.175 ;
 END
 PORT
  LAYER ME4 ;
  RECT 535.321 0.000 536.041 46.394 ;
 END
 PORT
  LAYER ME4 ;
  RECT 541.517 45.394 541.857 293.175 ;
 END
 PORT
  LAYER ME4 ;
  RECT 539.325 0.000 540.045 46.394 ;
 END
 PORT
  LAYER ME4 ;
  RECT 545.521 45.394 545.861 293.175 ;
 END
 PORT
  LAYER ME4 ;
  RECT 543.329 0.000 544.049 46.394 ;
 END
 PORT
  LAYER ME4 ;
  RECT 549.525 45.394 549.865 293.175 ;
 END
 PORT
  LAYER ME4 ;
  RECT 547.333 0.000 548.053 46.394 ;
 END
 PORT
  LAYER ME4 ;
  RECT 553.529 45.394 553.869 293.175 ;
 END
 PORT
  LAYER ME4 ;
  RECT 551.337 0.000 552.057 46.394 ;
 END
 PORT
  LAYER ME4 ;
  RECT 556.311 0.000 556.691 293.175 ;
 END
 PORT
  LAYER ME4 ;
  RECT 282.197 0.000 282.797 293.175 ;
 END
 PORT
  LAYER ME4 ;
  RECT 286.377 0.000 287.097 293.175 ;
 END
 PORT
  LAYER ME4 ;
  RECT 288.487 0.000 289.607 293.175 ;
 END
 PORT
  LAYER ME4 ;
  RECT 294.517 0.000 295.237 293.175 ;
 END
 PORT
  LAYER ME4 ;
  RECT 296.453 1.781 296.833 293.175 ;
 END
 PORT
  LAYER ME4 ;
  RECT 277.967 0.000 278.687 293.175 ;
 END
 PORT
  LAYER ME4 ;
  RECT 275.252 0.000 276.372 293.175 ;
 END
 PORT
  LAYER ME4 ;
  RECT 272.878 0.000 273.598 292.295 ;
 END
 PORT
  LAYER ME4 ;
  RECT 270.838 1.781 271.558 293.175 ;
 END
 PORT
  LAYER ME4 ;
  RECT 268.718 0.000 269.438 293.175 ;
 END
 PORT
  LAYER ME4 ;
  RECT 266.678 1.781 267.398 293.175 ;
 END
 PORT
  LAYER ME4 ;
  RECT 264.558 0.000 265.278 293.175 ;
 END
 PORT
  LAYER ME4 ;
  RECT 262.518 1.781 263.238 293.175 ;
 END
 PORT
  LAYER ME4 ;
  RECT 0.920 0.000 1.300 293.175 ;
 END
 PORT
  LAYER ME4 ;
  RECT 5.744 45.394 6.084 293.175 ;
 END
 PORT
  LAYER ME4 ;
  RECT 3.552 0.000 4.272 46.394 ;
 END
 PORT
  LAYER ME4 ;
  RECT 9.748 45.394 10.088 293.175 ;
 END
 PORT
  LAYER ME4 ;
  RECT 7.556 0.000 8.276 46.394 ;
 END
 PORT
  LAYER ME4 ;
  RECT 13.752 45.394 14.092 293.175 ;
 END
 PORT
  LAYER ME4 ;
  RECT 11.560 0.000 12.280 46.394 ;
 END
 PORT
  LAYER ME4 ;
  RECT 17.756 45.394 18.096 293.175 ;
 END
 PORT
  LAYER ME4 ;
  RECT 15.564 0.000 16.284 46.394 ;
 END
 PORT
  LAYER ME4 ;
  RECT 21.760 45.394 22.100 293.175 ;
 END
 PORT
  LAYER ME4 ;
  RECT 19.568 0.000 20.288 46.394 ;
 END
 PORT
  LAYER ME4 ;
  RECT 25.764 45.394 26.104 293.175 ;
 END
 PORT
  LAYER ME4 ;
  RECT 23.572 0.000 24.292 46.394 ;
 END
 PORT
  LAYER ME4 ;
  RECT 29.768 45.394 30.108 293.175 ;
 END
 PORT
  LAYER ME4 ;
  RECT 27.576 0.000 28.296 46.394 ;
 END
 PORT
  LAYER ME4 ;
  RECT 33.772 45.394 34.112 293.175 ;
 END
 PORT
  LAYER ME4 ;
  RECT 31.580 0.000 32.300 46.394 ;
 END
 PORT
  LAYER ME4 ;
  RECT 37.776 45.394 38.116 293.175 ;
 END
 PORT
  LAYER ME4 ;
  RECT 35.584 0.000 36.304 46.394 ;
 END
 PORT
  LAYER ME4 ;
  RECT 41.780 45.394 42.120 293.175 ;
 END
 PORT
  LAYER ME4 ;
  RECT 39.588 0.000 40.308 46.394 ;
 END
 PORT
  LAYER ME4 ;
  RECT 45.784 45.394 46.124 293.175 ;
 END
 PORT
  LAYER ME4 ;
  RECT 43.592 0.000 44.312 46.394 ;
 END
 PORT
  LAYER ME4 ;
  RECT 49.788 45.394 50.128 293.175 ;
 END
 PORT
  LAYER ME4 ;
  RECT 47.596 0.000 48.316 46.394 ;
 END
 PORT
  LAYER ME4 ;
  RECT 53.792 45.394 54.132 293.175 ;
 END
 PORT
  LAYER ME4 ;
  RECT 51.600 0.000 52.320 46.394 ;
 END
 PORT
  LAYER ME4 ;
  RECT 57.796 45.394 58.136 293.175 ;
 END
 PORT
  LAYER ME4 ;
  RECT 55.604 0.000 56.324 46.394 ;
 END
 PORT
  LAYER ME4 ;
  RECT 61.800 45.394 62.140 293.175 ;
 END
 PORT
  LAYER ME4 ;
  RECT 59.608 0.000 60.328 46.394 ;
 END
 PORT
  LAYER ME4 ;
  RECT 65.804 45.394 66.144 293.175 ;
 END
 PORT
  LAYER ME4 ;
  RECT 63.612 0.000 64.332 46.394 ;
 END
 PORT
  LAYER ME4 ;
  RECT 69.808 45.394 70.148 293.175 ;
 END
 PORT
  LAYER ME4 ;
  RECT 67.616 0.000 68.336 46.394 ;
 END
 PORT
  LAYER ME4 ;
  RECT 73.812 45.394 74.152 293.175 ;
 END
 PORT
  LAYER ME4 ;
  RECT 71.620 0.000 72.340 46.394 ;
 END
 PORT
  LAYER ME4 ;
  RECT 77.816 45.394 78.156 293.175 ;
 END
 PORT
  LAYER ME4 ;
  RECT 75.624 0.000 76.344 46.394 ;
 END
 PORT
  LAYER ME4 ;
  RECT 81.820 45.394 82.160 293.175 ;
 END
 PORT
  LAYER ME4 ;
  RECT 79.628 0.000 80.348 46.394 ;
 END
 PORT
  LAYER ME4 ;
  RECT 85.824 45.394 86.164 293.175 ;
 END
 PORT
  LAYER ME4 ;
  RECT 83.632 0.000 84.352 46.394 ;
 END
 PORT
  LAYER ME4 ;
  RECT 89.828 45.394 90.168 293.175 ;
 END
 PORT
  LAYER ME4 ;
  RECT 87.636 0.000 88.356 46.394 ;
 END
 PORT
  LAYER ME4 ;
  RECT 93.832 45.394 94.172 293.175 ;
 END
 PORT
  LAYER ME4 ;
  RECT 91.640 0.000 92.360 46.394 ;
 END
 PORT
  LAYER ME4 ;
  RECT 97.836 45.394 98.176 293.175 ;
 END
 PORT
  LAYER ME4 ;
  RECT 95.644 0.000 96.364 46.394 ;
 END
 PORT
  LAYER ME4 ;
  RECT 101.840 45.394 102.180 293.175 ;
 END
 PORT
  LAYER ME4 ;
  RECT 99.648 0.000 100.368 46.394 ;
 END
 PORT
  LAYER ME4 ;
  RECT 105.844 45.394 106.184 293.175 ;
 END
 PORT
  LAYER ME4 ;
  RECT 103.652 0.000 104.372 46.394 ;
 END
 PORT
  LAYER ME4 ;
  RECT 109.848 45.394 110.188 293.175 ;
 END
 PORT
  LAYER ME4 ;
  RECT 107.656 0.000 108.376 46.394 ;
 END
 PORT
  LAYER ME4 ;
  RECT 113.852 45.394 114.192 293.175 ;
 END
 PORT
  LAYER ME4 ;
  RECT 111.660 0.000 112.380 46.394 ;
 END
 PORT
  LAYER ME4 ;
  RECT 117.856 45.394 118.196 293.175 ;
 END
 PORT
  LAYER ME4 ;
  RECT 115.664 0.000 116.384 46.394 ;
 END
 PORT
  LAYER ME4 ;
  RECT 121.860 45.394 122.200 293.175 ;
 END
 PORT
  LAYER ME4 ;
  RECT 119.668 0.000 120.388 46.394 ;
 END
 PORT
  LAYER ME4 ;
  RECT 125.864 45.394 126.204 293.175 ;
 END
 PORT
  LAYER ME4 ;
  RECT 123.672 0.000 124.392 46.394 ;
 END
 PORT
  LAYER ME4 ;
  RECT 129.868 45.394 130.208 293.175 ;
 END
 PORT
  LAYER ME4 ;
  RECT 127.676 0.000 128.396 46.394 ;
 END
 PORT
  LAYER ME4 ;
  RECT 133.872 45.394 134.212 293.175 ;
 END
 PORT
  LAYER ME4 ;
  RECT 131.680 0.000 132.400 46.394 ;
 END
 PORT
  LAYER ME4 ;
  RECT 137.876 45.394 138.216 293.175 ;
 END
 PORT
  LAYER ME4 ;
  RECT 135.684 0.000 136.404 46.394 ;
 END
 PORT
  LAYER ME4 ;
  RECT 141.880 45.394 142.220 293.175 ;
 END
 PORT
  LAYER ME4 ;
  RECT 139.688 0.000 140.408 46.394 ;
 END
 PORT
  LAYER ME4 ;
  RECT 145.884 45.394 146.224 293.175 ;
 END
 PORT
  LAYER ME4 ;
  RECT 143.692 0.000 144.412 46.394 ;
 END
 PORT
  LAYER ME4 ;
  RECT 149.888 45.394 150.228 293.175 ;
 END
 PORT
  LAYER ME4 ;
  RECT 147.696 0.000 148.416 46.394 ;
 END
 PORT
  LAYER ME4 ;
  RECT 153.892 45.394 154.232 293.175 ;
 END
 PORT
  LAYER ME4 ;
  RECT 151.700 0.000 152.420 46.394 ;
 END
 PORT
  LAYER ME4 ;
  RECT 157.896 45.394 158.236 293.175 ;
 END
 PORT
  LAYER ME4 ;
  RECT 155.704 0.000 156.424 46.394 ;
 END
 PORT
  LAYER ME4 ;
  RECT 161.900 45.394 162.240 293.175 ;
 END
 PORT
  LAYER ME4 ;
  RECT 159.708 0.000 160.428 46.394 ;
 END
 PORT
  LAYER ME4 ;
  RECT 165.904 45.394 166.244 293.175 ;
 END
 PORT
  LAYER ME4 ;
  RECT 163.712 0.000 164.432 46.394 ;
 END
 PORT
  LAYER ME4 ;
  RECT 169.908 45.394 170.248 293.175 ;
 END
 PORT
  LAYER ME4 ;
  RECT 167.716 0.000 168.436 46.394 ;
 END
 PORT
  LAYER ME4 ;
  RECT 173.912 45.394 174.252 293.175 ;
 END
 PORT
  LAYER ME4 ;
  RECT 171.720 0.000 172.440 46.394 ;
 END
 PORT
  LAYER ME4 ;
  RECT 177.916 45.394 178.256 293.175 ;
 END
 PORT
  LAYER ME4 ;
  RECT 175.724 0.000 176.444 46.394 ;
 END
 PORT
  LAYER ME4 ;
  RECT 181.920 45.394 182.260 293.175 ;
 END
 PORT
  LAYER ME4 ;
  RECT 179.728 0.000 180.448 46.394 ;
 END
 PORT
  LAYER ME4 ;
  RECT 185.924 45.394 186.264 293.175 ;
 END
 PORT
  LAYER ME4 ;
  RECT 183.732 0.000 184.452 46.394 ;
 END
 PORT
  LAYER ME4 ;
  RECT 189.928 45.394 190.268 293.175 ;
 END
 PORT
  LAYER ME4 ;
  RECT 187.736 0.000 188.456 46.394 ;
 END
 PORT
  LAYER ME4 ;
  RECT 193.932 45.394 194.272 293.175 ;
 END
 PORT
  LAYER ME4 ;
  RECT 191.740 0.000 192.460 46.394 ;
 END
 PORT
  LAYER ME4 ;
  RECT 197.936 45.394 198.276 293.175 ;
 END
 PORT
  LAYER ME4 ;
  RECT 195.744 0.000 196.464 46.394 ;
 END
 PORT
  LAYER ME4 ;
  RECT 201.940 45.394 202.280 293.175 ;
 END
 PORT
  LAYER ME4 ;
  RECT 199.748 0.000 200.468 46.394 ;
 END
 PORT
  LAYER ME4 ;
  RECT 205.944 45.394 206.284 293.175 ;
 END
 PORT
  LAYER ME4 ;
  RECT 203.752 0.000 204.472 46.394 ;
 END
 PORT
  LAYER ME4 ;
  RECT 209.948 45.394 210.288 293.175 ;
 END
 PORT
  LAYER ME4 ;
  RECT 207.756 0.000 208.476 46.394 ;
 END
 PORT
  LAYER ME4 ;
  RECT 213.952 45.394 214.292 293.175 ;
 END
 PORT
  LAYER ME4 ;
  RECT 211.760 0.000 212.480 46.394 ;
 END
 PORT
  LAYER ME4 ;
  RECT 217.956 45.394 218.296 293.175 ;
 END
 PORT
  LAYER ME4 ;
  RECT 215.764 0.000 216.484 46.394 ;
 END
 PORT
  LAYER ME4 ;
  RECT 221.960 45.394 222.300 293.175 ;
 END
 PORT
  LAYER ME4 ;
  RECT 219.768 0.000 220.488 46.394 ;
 END
 PORT
  LAYER ME4 ;
  RECT 225.964 45.394 226.304 293.175 ;
 END
 PORT
  LAYER ME4 ;
  RECT 223.772 0.000 224.492 46.394 ;
 END
 PORT
  LAYER ME4 ;
  RECT 229.968 45.394 230.308 293.175 ;
 END
 PORT
  LAYER ME4 ;
  RECT 227.776 0.000 228.496 46.394 ;
 END
 PORT
  LAYER ME4 ;
  RECT 233.972 45.394 234.312 293.175 ;
 END
 PORT
  LAYER ME4 ;
  RECT 231.780 0.000 232.500 46.394 ;
 END
 PORT
  LAYER ME4 ;
  RECT 237.976 45.394 238.316 293.175 ;
 END
 PORT
  LAYER ME4 ;
  RECT 235.784 0.000 236.504 46.394 ;
 END
 PORT
  LAYER ME4 ;
  RECT 241.980 45.394 242.320 293.175 ;
 END
 PORT
  LAYER ME4 ;
  RECT 239.788 0.000 240.508 46.394 ;
 END
 PORT
  LAYER ME4 ;
  RECT 245.984 45.394 246.324 293.175 ;
 END
 PORT
  LAYER ME4 ;
  RECT 243.792 0.000 244.512 46.394 ;
 END
 PORT
  LAYER ME4 ;
  RECT 249.988 45.394 250.328 293.175 ;
 END
 PORT
  LAYER ME4 ;
  RECT 247.796 0.000 248.516 46.394 ;
 END
 PORT
  LAYER ME4 ;
  RECT 253.992 45.394 254.332 293.175 ;
 END
 PORT
  LAYER ME4 ;
  RECT 251.800 0.000 252.520 46.394 ;
 END
 PORT
  LAYER ME4 ;
  RECT 257.996 45.394 258.336 293.175 ;
 END
 PORT
  LAYER ME4 ;
  RECT 255.804 0.000 256.524 46.394 ;
 END
 PORT
  LAYER ME4 ;
  RECT 260.778 0.000 261.158 293.175 ;
 END
 PORT
  LAYER ME4 ;
  RECT 299.275 47.744 299.615 293.175 ;
 END
 PORT
  LAYER ME4 ;
  RECT 303.279 47.744 303.619 293.175 ;
 END
 PORT
  LAYER ME4 ;
  RECT 307.283 47.744 307.623 293.175 ;
 END
 PORT
  LAYER ME4 ;
  RECT 311.287 47.744 311.627 293.175 ;
 END
 PORT
  LAYER ME4 ;
  RECT 315.291 47.744 315.631 293.175 ;
 END
 PORT
  LAYER ME4 ;
  RECT 319.295 47.744 319.635 293.175 ;
 END
 PORT
  LAYER ME4 ;
  RECT 323.299 47.744 323.639 293.175 ;
 END
 PORT
  LAYER ME4 ;
  RECT 327.303 47.744 327.643 293.175 ;
 END
 PORT
  LAYER ME4 ;
  RECT 331.307 47.744 331.647 293.175 ;
 END
 PORT
  LAYER ME4 ;
  RECT 335.311 47.744 335.651 293.175 ;
 END
 PORT
  LAYER ME4 ;
  RECT 339.315 47.744 339.655 293.175 ;
 END
 PORT
  LAYER ME4 ;
  RECT 343.319 47.744 343.659 293.175 ;
 END
 PORT
  LAYER ME4 ;
  RECT 347.323 47.744 347.663 293.175 ;
 END
 PORT
  LAYER ME4 ;
  RECT 351.327 47.744 351.667 293.175 ;
 END
 PORT
  LAYER ME4 ;
  RECT 355.331 47.744 355.671 293.175 ;
 END
 PORT
  LAYER ME4 ;
  RECT 359.335 47.744 359.675 293.175 ;
 END
 PORT
  LAYER ME4 ;
  RECT 363.339 47.744 363.679 293.175 ;
 END
 PORT
  LAYER ME4 ;
  RECT 367.343 47.744 367.683 293.175 ;
 END
 PORT
  LAYER ME4 ;
  RECT 371.347 47.744 371.687 293.175 ;
 END
 PORT
  LAYER ME4 ;
  RECT 375.351 47.744 375.691 293.175 ;
 END
 PORT
  LAYER ME4 ;
  RECT 379.355 47.744 379.695 293.175 ;
 END
 PORT
  LAYER ME4 ;
  RECT 383.359 47.744 383.699 293.175 ;
 END
 PORT
  LAYER ME4 ;
  RECT 387.363 47.744 387.703 293.175 ;
 END
 PORT
  LAYER ME4 ;
  RECT 391.367 47.744 391.707 293.175 ;
 END
 PORT
  LAYER ME4 ;
  RECT 395.371 47.744 395.711 293.175 ;
 END
 PORT
  LAYER ME4 ;
  RECT 399.375 47.744 399.715 293.175 ;
 END
 PORT
  LAYER ME4 ;
  RECT 403.379 47.744 403.719 293.175 ;
 END
 PORT
  LAYER ME4 ;
  RECT 407.383 47.744 407.723 293.175 ;
 END
 PORT
  LAYER ME4 ;
  RECT 411.387 47.744 411.727 293.175 ;
 END
 PORT
  LAYER ME4 ;
  RECT 415.391 47.744 415.731 293.175 ;
 END
 PORT
  LAYER ME4 ;
  RECT 419.395 47.744 419.735 293.175 ;
 END
 PORT
  LAYER ME4 ;
  RECT 423.399 47.744 423.739 293.175 ;
 END
 PORT
  LAYER ME4 ;
  RECT 427.403 47.744 427.743 293.175 ;
 END
 PORT
  LAYER ME4 ;
  RECT 431.407 47.744 431.747 293.175 ;
 END
 PORT
  LAYER ME4 ;
  RECT 435.411 47.744 435.751 293.175 ;
 END
 PORT
  LAYER ME4 ;
  RECT 439.415 47.744 439.755 293.175 ;
 END
 PORT
  LAYER ME4 ;
  RECT 443.419 47.744 443.759 293.175 ;
 END
 PORT
  LAYER ME4 ;
  RECT 447.423 47.744 447.763 293.175 ;
 END
 PORT
  LAYER ME4 ;
  RECT 451.427 47.744 451.767 293.175 ;
 END
 PORT
  LAYER ME4 ;
  RECT 455.431 47.744 455.771 293.175 ;
 END
 PORT
  LAYER ME4 ;
  RECT 459.435 47.744 459.775 293.175 ;
 END
 PORT
  LAYER ME4 ;
  RECT 463.439 47.744 463.779 293.175 ;
 END
 PORT
  LAYER ME4 ;
  RECT 467.443 47.744 467.783 293.175 ;
 END
 PORT
  LAYER ME4 ;
  RECT 471.447 47.744 471.787 293.175 ;
 END
 PORT
  LAYER ME4 ;
  RECT 475.451 47.744 475.791 293.175 ;
 END
 PORT
  LAYER ME4 ;
  RECT 479.455 47.744 479.795 293.175 ;
 END
 PORT
  LAYER ME4 ;
  RECT 483.459 47.744 483.799 293.175 ;
 END
 PORT
  LAYER ME4 ;
  RECT 487.463 47.744 487.803 293.175 ;
 END
 PORT
  LAYER ME4 ;
  RECT 491.467 47.744 491.807 293.175 ;
 END
 PORT
  LAYER ME4 ;
  RECT 495.471 47.744 495.811 293.175 ;
 END
 PORT
  LAYER ME4 ;
  RECT 499.475 47.744 499.815 293.175 ;
 END
 PORT
  LAYER ME4 ;
  RECT 503.479 47.744 503.819 293.175 ;
 END
 PORT
  LAYER ME4 ;
  RECT 507.483 47.744 507.823 293.175 ;
 END
 PORT
  LAYER ME4 ;
  RECT 511.487 47.744 511.827 293.175 ;
 END
 PORT
  LAYER ME4 ;
  RECT 515.491 47.744 515.831 293.175 ;
 END
 PORT
  LAYER ME4 ;
  RECT 519.495 47.744 519.835 293.175 ;
 END
 PORT
  LAYER ME4 ;
  RECT 523.499 47.744 523.839 293.175 ;
 END
 PORT
  LAYER ME4 ;
  RECT 527.503 47.744 527.843 293.175 ;
 END
 PORT
  LAYER ME4 ;
  RECT 531.507 47.744 531.847 293.175 ;
 END
 PORT
  LAYER ME4 ;
  RECT 535.511 47.744 535.851 293.175 ;
 END
 PORT
  LAYER ME4 ;
  RECT 539.515 47.744 539.855 293.175 ;
 END
 PORT
  LAYER ME4 ;
  RECT 543.519 47.744 543.859 293.175 ;
 END
 PORT
  LAYER ME4 ;
  RECT 547.523 47.744 547.863 293.175 ;
 END
 PORT
  LAYER ME4 ;
  RECT 551.527 47.744 551.867 293.175 ;
 END
 PORT
  LAYER ME4 ;
  RECT 3.742 47.744 4.082 293.175 ;
 END
 PORT
  LAYER ME4 ;
  RECT 7.746 47.744 8.086 293.175 ;
 END
 PORT
  LAYER ME4 ;
  RECT 11.750 47.744 12.090 293.175 ;
 END
 PORT
  LAYER ME4 ;
  RECT 15.754 47.744 16.094 293.175 ;
 END
 PORT
  LAYER ME4 ;
  RECT 19.758 47.744 20.098 293.175 ;
 END
 PORT
  LAYER ME4 ;
  RECT 23.762 47.744 24.102 293.175 ;
 END
 PORT
  LAYER ME4 ;
  RECT 27.766 47.744 28.106 293.175 ;
 END
 PORT
  LAYER ME4 ;
  RECT 31.770 47.744 32.110 293.175 ;
 END
 PORT
  LAYER ME4 ;
  RECT 35.774 47.744 36.114 293.175 ;
 END
 PORT
  LAYER ME4 ;
  RECT 39.778 47.744 40.118 293.175 ;
 END
 PORT
  LAYER ME4 ;
  RECT 43.782 47.744 44.122 293.175 ;
 END
 PORT
  LAYER ME4 ;
  RECT 47.786 47.744 48.126 293.175 ;
 END
 PORT
  LAYER ME4 ;
  RECT 51.790 47.744 52.130 293.175 ;
 END
 PORT
  LAYER ME4 ;
  RECT 55.794 47.744 56.134 293.175 ;
 END
 PORT
  LAYER ME4 ;
  RECT 59.798 47.744 60.138 293.175 ;
 END
 PORT
  LAYER ME4 ;
  RECT 63.802 47.744 64.142 293.175 ;
 END
 PORT
  LAYER ME4 ;
  RECT 67.806 47.744 68.146 293.175 ;
 END
 PORT
  LAYER ME4 ;
  RECT 71.810 47.744 72.150 293.175 ;
 END
 PORT
  LAYER ME4 ;
  RECT 75.814 47.744 76.154 293.175 ;
 END
 PORT
  LAYER ME4 ;
  RECT 79.818 47.744 80.158 293.175 ;
 END
 PORT
  LAYER ME4 ;
  RECT 83.822 47.744 84.162 293.175 ;
 END
 PORT
  LAYER ME4 ;
  RECT 87.826 47.744 88.166 293.175 ;
 END
 PORT
  LAYER ME4 ;
  RECT 91.830 47.744 92.170 293.175 ;
 END
 PORT
  LAYER ME4 ;
  RECT 95.834 47.744 96.174 293.175 ;
 END
 PORT
  LAYER ME4 ;
  RECT 99.838 47.744 100.178 293.175 ;
 END
 PORT
  LAYER ME4 ;
  RECT 103.842 47.744 104.182 293.175 ;
 END
 PORT
  LAYER ME4 ;
  RECT 107.846 47.744 108.186 293.175 ;
 END
 PORT
  LAYER ME4 ;
  RECT 111.850 47.744 112.190 293.175 ;
 END
 PORT
  LAYER ME4 ;
  RECT 115.854 47.744 116.194 293.175 ;
 END
 PORT
  LAYER ME4 ;
  RECT 119.858 47.744 120.198 293.175 ;
 END
 PORT
  LAYER ME4 ;
  RECT 123.862 47.744 124.202 293.175 ;
 END
 PORT
  LAYER ME4 ;
  RECT 127.866 47.744 128.206 293.175 ;
 END
 PORT
  LAYER ME4 ;
  RECT 131.870 47.744 132.210 293.175 ;
 END
 PORT
  LAYER ME4 ;
  RECT 135.874 47.744 136.214 293.175 ;
 END
 PORT
  LAYER ME4 ;
  RECT 139.878 47.744 140.218 293.175 ;
 END
 PORT
  LAYER ME4 ;
  RECT 143.882 47.744 144.222 293.175 ;
 END
 PORT
  LAYER ME4 ;
  RECT 147.886 47.744 148.226 293.175 ;
 END
 PORT
  LAYER ME4 ;
  RECT 151.890 47.744 152.230 293.175 ;
 END
 PORT
  LAYER ME4 ;
  RECT 155.894 47.744 156.234 293.175 ;
 END
 PORT
  LAYER ME4 ;
  RECT 159.898 47.744 160.238 293.175 ;
 END
 PORT
  LAYER ME4 ;
  RECT 163.902 47.744 164.242 293.175 ;
 END
 PORT
  LAYER ME4 ;
  RECT 167.906 47.744 168.246 293.175 ;
 END
 PORT
  LAYER ME4 ;
  RECT 171.910 47.744 172.250 293.175 ;
 END
 PORT
  LAYER ME4 ;
  RECT 175.914 47.744 176.254 293.175 ;
 END
 PORT
  LAYER ME4 ;
  RECT 179.918 47.744 180.258 293.175 ;
 END
 PORT
  LAYER ME4 ;
  RECT 183.922 47.744 184.262 293.175 ;
 END
 PORT
  LAYER ME4 ;
  RECT 187.926 47.744 188.266 293.175 ;
 END
 PORT
  LAYER ME4 ;
  RECT 191.930 47.744 192.270 293.175 ;
 END
 PORT
  LAYER ME4 ;
  RECT 195.934 47.744 196.274 293.175 ;
 END
 PORT
  LAYER ME4 ;
  RECT 199.938 47.744 200.278 293.175 ;
 END
 PORT
  LAYER ME4 ;
  RECT 203.942 47.744 204.282 293.175 ;
 END
 PORT
  LAYER ME4 ;
  RECT 207.946 47.744 208.286 293.175 ;
 END
 PORT
  LAYER ME4 ;
  RECT 211.950 47.744 212.290 293.175 ;
 END
 PORT
  LAYER ME4 ;
  RECT 215.954 47.744 216.294 293.175 ;
 END
 PORT
  LAYER ME4 ;
  RECT 219.958 47.744 220.298 293.175 ;
 END
 PORT
  LAYER ME4 ;
  RECT 223.962 47.744 224.302 293.175 ;
 END
 PORT
  LAYER ME4 ;
  RECT 227.966 47.744 228.306 293.175 ;
 END
 PORT
  LAYER ME4 ;
  RECT 231.970 47.744 232.310 293.175 ;
 END
 PORT
  LAYER ME4 ;
  RECT 235.974 47.744 236.314 293.175 ;
 END
 PORT
  LAYER ME4 ;
  RECT 239.978 47.744 240.318 293.175 ;
 END
 PORT
  LAYER ME4 ;
  RECT 243.982 47.744 244.322 293.175 ;
 END
 PORT
  LAYER ME4 ;
  RECT 247.986 47.744 248.326 293.175 ;
 END
 PORT
  LAYER ME4 ;
  RECT 251.990 47.744 252.330 293.175 ;
 END
 PORT
  LAYER ME4 ;
  RECT 255.994 47.744 256.334 293.175 ;
 END
END VCC
PIN DI63
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 257.286 0.000 257.606 0.600 ;
  LAYER ME3 ;
  RECT 257.286 0.000 257.606 0.600 ;
  LAYER ME2 ;
  RECT 257.286 0.000 257.606 0.600 ;
  LAYER ME1 ;
  RECT 257.286 0.000 257.606 0.600 ;
 END
 ANTENNAPARTIALMETALAREA                  1.058 LAYER ME2 ;
 ANTENNAGATEAREA                          0.072 LAYER ME2 ;
 ANTENNAGATEAREA                          0.072 LAYER ME3 ;
 ANTENNAGATEAREA                          0.072 LAYER ME4 ;
 ANTENNADIFFAREA                          0.160 LAYER ME2 ;
 ANTENNADIFFAREA                          0.160 LAYER ME3 ;
 ANTENNADIFFAREA                          0.160 LAYER ME4 ;
 ANTENNAMAXAREACAR                       21.782 LAYER ME2 ;
 ANTENNAMAXAREACAR                       24.449 LAYER ME3 ;
 ANTENNAMAXAREACAR                       27.116 LAYER ME4 ;
END DI63
PIN DO63
  DIRECTION OUTPUT ;
 PORT
  LAYER ME4 ;
  RECT 256.724 0.000 257.044 0.600 ;
  LAYER ME3 ;
  RECT 256.724 0.000 257.044 0.600 ;
  LAYER ME2 ;
  RECT 256.724 0.000 257.044 0.600 ;
  LAYER ME1 ;
  RECT 256.724 0.000 257.044 0.600 ;
 END
 ANTENNAPARTIALMETALAREA                  5.273 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME3 ;
 ANTENNADIFFAREA                          1.293 LAYER ME4 ;
END DO63
PIN DI62
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 253.282 0.000 253.602 0.600 ;
  LAYER ME3 ;
  RECT 253.282 0.000 253.602 0.600 ;
  LAYER ME2 ;
  RECT 253.282 0.000 253.602 0.600 ;
  LAYER ME1 ;
  RECT 253.282 0.000 253.602 0.600 ;
 END
 ANTENNAPARTIALMETALAREA                  1.058 LAYER ME2 ;
 ANTENNAGATEAREA                          0.072 LAYER ME2 ;
 ANTENNAGATEAREA                          0.072 LAYER ME3 ;
 ANTENNAGATEAREA                          0.072 LAYER ME4 ;
 ANTENNADIFFAREA                          0.160 LAYER ME2 ;
 ANTENNADIFFAREA                          0.160 LAYER ME3 ;
 ANTENNADIFFAREA                          0.160 LAYER ME4 ;
 ANTENNAMAXAREACAR                       21.782 LAYER ME2 ;
 ANTENNAMAXAREACAR                       24.449 LAYER ME3 ;
 ANTENNAMAXAREACAR                       27.116 LAYER ME4 ;
END DI62
PIN DO62
  DIRECTION OUTPUT ;
 PORT
  LAYER ME4 ;
  RECT 252.720 0.000 253.040 0.600 ;
  LAYER ME3 ;
  RECT 252.720 0.000 253.040 0.600 ;
  LAYER ME2 ;
  RECT 252.720 0.000 253.040 0.600 ;
  LAYER ME1 ;
  RECT 252.720 0.000 253.040 0.600 ;
 END
 ANTENNAPARTIALMETALAREA                  5.273 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME3 ;
 ANTENNADIFFAREA                          1.293 LAYER ME4 ;
END DO62
PIN DI61
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 249.278 0.000 249.598 0.600 ;
  LAYER ME3 ;
  RECT 249.278 0.000 249.598 0.600 ;
  LAYER ME2 ;
  RECT 249.278 0.000 249.598 0.600 ;
  LAYER ME1 ;
  RECT 249.278 0.000 249.598 0.600 ;
 END
 ANTENNAPARTIALMETALAREA                  1.058 LAYER ME2 ;
 ANTENNAGATEAREA                          0.072 LAYER ME2 ;
 ANTENNAGATEAREA                          0.072 LAYER ME3 ;
 ANTENNAGATEAREA                          0.072 LAYER ME4 ;
 ANTENNADIFFAREA                          0.160 LAYER ME2 ;
 ANTENNADIFFAREA                          0.160 LAYER ME3 ;
 ANTENNADIFFAREA                          0.160 LAYER ME4 ;
 ANTENNAMAXAREACAR                       21.782 LAYER ME2 ;
 ANTENNAMAXAREACAR                       24.449 LAYER ME3 ;
 ANTENNAMAXAREACAR                       27.116 LAYER ME4 ;
END DI61
PIN DO61
  DIRECTION OUTPUT ;
 PORT
  LAYER ME4 ;
  RECT 248.716 0.000 249.036 0.600 ;
  LAYER ME3 ;
  RECT 248.716 0.000 249.036 0.600 ;
  LAYER ME2 ;
  RECT 248.716 0.000 249.036 0.600 ;
  LAYER ME1 ;
  RECT 248.716 0.000 249.036 0.600 ;
 END
 ANTENNAPARTIALMETALAREA                  5.273 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME3 ;
 ANTENNADIFFAREA                          1.293 LAYER ME4 ;
END DO61
PIN DI60
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 245.274 0.000 245.594 0.600 ;
  LAYER ME3 ;
  RECT 245.274 0.000 245.594 0.600 ;
  LAYER ME2 ;
  RECT 245.274 0.000 245.594 0.600 ;
  LAYER ME1 ;
  RECT 245.274 0.000 245.594 0.600 ;
 END
 ANTENNAPARTIALMETALAREA                  1.058 LAYER ME2 ;
 ANTENNAGATEAREA                          0.072 LAYER ME2 ;
 ANTENNAGATEAREA                          0.072 LAYER ME3 ;
 ANTENNAGATEAREA                          0.072 LAYER ME4 ;
 ANTENNADIFFAREA                          0.160 LAYER ME2 ;
 ANTENNADIFFAREA                          0.160 LAYER ME3 ;
 ANTENNADIFFAREA                          0.160 LAYER ME4 ;
 ANTENNAMAXAREACAR                       21.782 LAYER ME2 ;
 ANTENNAMAXAREACAR                       24.449 LAYER ME3 ;
 ANTENNAMAXAREACAR                       27.116 LAYER ME4 ;
END DI60
PIN DO60
  DIRECTION OUTPUT ;
 PORT
  LAYER ME4 ;
  RECT 244.712 0.000 245.032 0.600 ;
  LAYER ME3 ;
  RECT 244.712 0.000 245.032 0.600 ;
  LAYER ME2 ;
  RECT 244.712 0.000 245.032 0.600 ;
  LAYER ME1 ;
  RECT 244.712 0.000 245.032 0.600 ;
 END
 ANTENNAPARTIALMETALAREA                  5.273 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME3 ;
 ANTENNADIFFAREA                          1.293 LAYER ME4 ;
END DO60
PIN DI59
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 241.270 0.000 241.590 0.600 ;
  LAYER ME3 ;
  RECT 241.270 0.000 241.590 0.600 ;
  LAYER ME2 ;
  RECT 241.270 0.000 241.590 0.600 ;
  LAYER ME1 ;
  RECT 241.270 0.000 241.590 0.600 ;
 END
 ANTENNAPARTIALMETALAREA                  1.058 LAYER ME2 ;
 ANTENNAGATEAREA                          0.072 LAYER ME2 ;
 ANTENNAGATEAREA                          0.072 LAYER ME3 ;
 ANTENNAGATEAREA                          0.072 LAYER ME4 ;
 ANTENNADIFFAREA                          0.160 LAYER ME2 ;
 ANTENNADIFFAREA                          0.160 LAYER ME3 ;
 ANTENNADIFFAREA                          0.160 LAYER ME4 ;
 ANTENNAMAXAREACAR                       21.782 LAYER ME2 ;
 ANTENNAMAXAREACAR                       24.449 LAYER ME3 ;
 ANTENNAMAXAREACAR                       27.116 LAYER ME4 ;
END DI59
PIN DO59
  DIRECTION OUTPUT ;
 PORT
  LAYER ME4 ;
  RECT 240.708 0.000 241.028 0.600 ;
  LAYER ME3 ;
  RECT 240.708 0.000 241.028 0.600 ;
  LAYER ME2 ;
  RECT 240.708 0.000 241.028 0.600 ;
  LAYER ME1 ;
  RECT 240.708 0.000 241.028 0.600 ;
 END
 ANTENNAPARTIALMETALAREA                  5.273 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME3 ;
 ANTENNADIFFAREA                          1.293 LAYER ME4 ;
END DO59
PIN DI58
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 237.266 0.000 237.586 0.600 ;
  LAYER ME3 ;
  RECT 237.266 0.000 237.586 0.600 ;
  LAYER ME2 ;
  RECT 237.266 0.000 237.586 0.600 ;
  LAYER ME1 ;
  RECT 237.266 0.000 237.586 0.600 ;
 END
 ANTENNAPARTIALMETALAREA                  1.058 LAYER ME2 ;
 ANTENNAGATEAREA                          0.072 LAYER ME2 ;
 ANTENNAGATEAREA                          0.072 LAYER ME3 ;
 ANTENNAGATEAREA                          0.072 LAYER ME4 ;
 ANTENNADIFFAREA                          0.160 LAYER ME2 ;
 ANTENNADIFFAREA                          0.160 LAYER ME3 ;
 ANTENNADIFFAREA                          0.160 LAYER ME4 ;
 ANTENNAMAXAREACAR                       21.782 LAYER ME2 ;
 ANTENNAMAXAREACAR                       24.449 LAYER ME3 ;
 ANTENNAMAXAREACAR                       27.116 LAYER ME4 ;
END DI58
PIN DO58
  DIRECTION OUTPUT ;
 PORT
  LAYER ME4 ;
  RECT 236.704 0.000 237.024 0.600 ;
  LAYER ME3 ;
  RECT 236.704 0.000 237.024 0.600 ;
  LAYER ME2 ;
  RECT 236.704 0.000 237.024 0.600 ;
  LAYER ME1 ;
  RECT 236.704 0.000 237.024 0.600 ;
 END
 ANTENNAPARTIALMETALAREA                  5.273 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME3 ;
 ANTENNADIFFAREA                          1.293 LAYER ME4 ;
END DO58
PIN DI57
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 233.262 0.000 233.582 0.600 ;
  LAYER ME3 ;
  RECT 233.262 0.000 233.582 0.600 ;
  LAYER ME2 ;
  RECT 233.262 0.000 233.582 0.600 ;
  LAYER ME1 ;
  RECT 233.262 0.000 233.582 0.600 ;
 END
 ANTENNAPARTIALMETALAREA                  1.058 LAYER ME2 ;
 ANTENNAGATEAREA                          0.072 LAYER ME2 ;
 ANTENNAGATEAREA                          0.072 LAYER ME3 ;
 ANTENNAGATEAREA                          0.072 LAYER ME4 ;
 ANTENNADIFFAREA                          0.160 LAYER ME2 ;
 ANTENNADIFFAREA                          0.160 LAYER ME3 ;
 ANTENNADIFFAREA                          0.160 LAYER ME4 ;
 ANTENNAMAXAREACAR                       21.782 LAYER ME2 ;
 ANTENNAMAXAREACAR                       24.449 LAYER ME3 ;
 ANTENNAMAXAREACAR                       27.116 LAYER ME4 ;
END DI57
PIN DO57
  DIRECTION OUTPUT ;
 PORT
  LAYER ME4 ;
  RECT 232.700 0.000 233.020 0.600 ;
  LAYER ME3 ;
  RECT 232.700 0.000 233.020 0.600 ;
  LAYER ME2 ;
  RECT 232.700 0.000 233.020 0.600 ;
  LAYER ME1 ;
  RECT 232.700 0.000 233.020 0.600 ;
 END
 ANTENNAPARTIALMETALAREA                  5.273 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME3 ;
 ANTENNADIFFAREA                          1.293 LAYER ME4 ;
END DO57
PIN DI56
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 229.258 0.000 229.578 0.600 ;
  LAYER ME3 ;
  RECT 229.258 0.000 229.578 0.600 ;
  LAYER ME2 ;
  RECT 229.258 0.000 229.578 0.600 ;
  LAYER ME1 ;
  RECT 229.258 0.000 229.578 0.600 ;
 END
 ANTENNAPARTIALMETALAREA                  1.058 LAYER ME2 ;
 ANTENNAGATEAREA                          0.072 LAYER ME2 ;
 ANTENNAGATEAREA                          0.072 LAYER ME3 ;
 ANTENNAGATEAREA                          0.072 LAYER ME4 ;
 ANTENNADIFFAREA                          0.160 LAYER ME2 ;
 ANTENNADIFFAREA                          0.160 LAYER ME3 ;
 ANTENNADIFFAREA                          0.160 LAYER ME4 ;
 ANTENNAMAXAREACAR                       21.782 LAYER ME2 ;
 ANTENNAMAXAREACAR                       24.449 LAYER ME3 ;
 ANTENNAMAXAREACAR                       27.116 LAYER ME4 ;
END DI56
PIN DO56
  DIRECTION OUTPUT ;
 PORT
  LAYER ME4 ;
  RECT 228.696 0.000 229.016 0.600 ;
  LAYER ME3 ;
  RECT 228.696 0.000 229.016 0.600 ;
  LAYER ME2 ;
  RECT 228.696 0.000 229.016 0.600 ;
  LAYER ME1 ;
  RECT 228.696 0.000 229.016 0.600 ;
 END
 ANTENNAPARTIALMETALAREA                  5.273 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME3 ;
 ANTENNADIFFAREA                          1.293 LAYER ME4 ;
END DO56
PIN DI55
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 225.254 0.000 225.574 0.600 ;
  LAYER ME3 ;
  RECT 225.254 0.000 225.574 0.600 ;
  LAYER ME2 ;
  RECT 225.254 0.000 225.574 0.600 ;
  LAYER ME1 ;
  RECT 225.254 0.000 225.574 0.600 ;
 END
 ANTENNAPARTIALMETALAREA                  1.058 LAYER ME2 ;
 ANTENNAGATEAREA                          0.072 LAYER ME2 ;
 ANTENNAGATEAREA                          0.072 LAYER ME3 ;
 ANTENNAGATEAREA                          0.072 LAYER ME4 ;
 ANTENNADIFFAREA                          0.160 LAYER ME2 ;
 ANTENNADIFFAREA                          0.160 LAYER ME3 ;
 ANTENNADIFFAREA                          0.160 LAYER ME4 ;
 ANTENNAMAXAREACAR                       21.782 LAYER ME2 ;
 ANTENNAMAXAREACAR                       24.449 LAYER ME3 ;
 ANTENNAMAXAREACAR                       27.116 LAYER ME4 ;
END DI55
PIN DO55
  DIRECTION OUTPUT ;
 PORT
  LAYER ME4 ;
  RECT 224.692 0.000 225.012 0.600 ;
  LAYER ME3 ;
  RECT 224.692 0.000 225.012 0.600 ;
  LAYER ME2 ;
  RECT 224.692 0.000 225.012 0.600 ;
  LAYER ME1 ;
  RECT 224.692 0.000 225.012 0.600 ;
 END
 ANTENNAPARTIALMETALAREA                  5.273 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME3 ;
 ANTENNADIFFAREA                          1.293 LAYER ME4 ;
END DO55
PIN DI54
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 221.250 0.000 221.570 0.600 ;
  LAYER ME3 ;
  RECT 221.250 0.000 221.570 0.600 ;
  LAYER ME2 ;
  RECT 221.250 0.000 221.570 0.600 ;
  LAYER ME1 ;
  RECT 221.250 0.000 221.570 0.600 ;
 END
 ANTENNAPARTIALMETALAREA                  1.058 LAYER ME2 ;
 ANTENNAGATEAREA                          0.072 LAYER ME2 ;
 ANTENNAGATEAREA                          0.072 LAYER ME3 ;
 ANTENNAGATEAREA                          0.072 LAYER ME4 ;
 ANTENNADIFFAREA                          0.160 LAYER ME2 ;
 ANTENNADIFFAREA                          0.160 LAYER ME3 ;
 ANTENNADIFFAREA                          0.160 LAYER ME4 ;
 ANTENNAMAXAREACAR                       21.782 LAYER ME2 ;
 ANTENNAMAXAREACAR                       24.449 LAYER ME3 ;
 ANTENNAMAXAREACAR                       27.116 LAYER ME4 ;
END DI54
PIN DO54
  DIRECTION OUTPUT ;
 PORT
  LAYER ME4 ;
  RECT 220.688 0.000 221.008 0.600 ;
  LAYER ME3 ;
  RECT 220.688 0.000 221.008 0.600 ;
  LAYER ME2 ;
  RECT 220.688 0.000 221.008 0.600 ;
  LAYER ME1 ;
  RECT 220.688 0.000 221.008 0.600 ;
 END
 ANTENNAPARTIALMETALAREA                  5.273 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME3 ;
 ANTENNADIFFAREA                          1.293 LAYER ME4 ;
END DO54
PIN DI53
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 217.246 0.000 217.566 0.600 ;
  LAYER ME3 ;
  RECT 217.246 0.000 217.566 0.600 ;
  LAYER ME2 ;
  RECT 217.246 0.000 217.566 0.600 ;
  LAYER ME1 ;
  RECT 217.246 0.000 217.566 0.600 ;
 END
 ANTENNAPARTIALMETALAREA                  1.058 LAYER ME2 ;
 ANTENNAGATEAREA                          0.072 LAYER ME2 ;
 ANTENNAGATEAREA                          0.072 LAYER ME3 ;
 ANTENNAGATEAREA                          0.072 LAYER ME4 ;
 ANTENNADIFFAREA                          0.160 LAYER ME2 ;
 ANTENNADIFFAREA                          0.160 LAYER ME3 ;
 ANTENNADIFFAREA                          0.160 LAYER ME4 ;
 ANTENNAMAXAREACAR                       21.782 LAYER ME2 ;
 ANTENNAMAXAREACAR                       24.449 LAYER ME3 ;
 ANTENNAMAXAREACAR                       27.116 LAYER ME4 ;
END DI53
PIN DO53
  DIRECTION OUTPUT ;
 PORT
  LAYER ME4 ;
  RECT 216.684 0.000 217.004 0.600 ;
  LAYER ME3 ;
  RECT 216.684 0.000 217.004 0.600 ;
  LAYER ME2 ;
  RECT 216.684 0.000 217.004 0.600 ;
  LAYER ME1 ;
  RECT 216.684 0.000 217.004 0.600 ;
 END
 ANTENNAPARTIALMETALAREA                  5.273 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME3 ;
 ANTENNADIFFAREA                          1.293 LAYER ME4 ;
END DO53
PIN DI52
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 213.242 0.000 213.562 0.600 ;
  LAYER ME3 ;
  RECT 213.242 0.000 213.562 0.600 ;
  LAYER ME2 ;
  RECT 213.242 0.000 213.562 0.600 ;
  LAYER ME1 ;
  RECT 213.242 0.000 213.562 0.600 ;
 END
 ANTENNAPARTIALMETALAREA                  1.058 LAYER ME2 ;
 ANTENNAGATEAREA                          0.072 LAYER ME2 ;
 ANTENNAGATEAREA                          0.072 LAYER ME3 ;
 ANTENNAGATEAREA                          0.072 LAYER ME4 ;
 ANTENNADIFFAREA                          0.160 LAYER ME2 ;
 ANTENNADIFFAREA                          0.160 LAYER ME3 ;
 ANTENNADIFFAREA                          0.160 LAYER ME4 ;
 ANTENNAMAXAREACAR                       21.782 LAYER ME2 ;
 ANTENNAMAXAREACAR                       24.449 LAYER ME3 ;
 ANTENNAMAXAREACAR                       27.116 LAYER ME4 ;
END DI52
PIN DO52
  DIRECTION OUTPUT ;
 PORT
  LAYER ME4 ;
  RECT 212.680 0.000 213.000 0.600 ;
  LAYER ME3 ;
  RECT 212.680 0.000 213.000 0.600 ;
  LAYER ME2 ;
  RECT 212.680 0.000 213.000 0.600 ;
  LAYER ME1 ;
  RECT 212.680 0.000 213.000 0.600 ;
 END
 ANTENNAPARTIALMETALAREA                  5.273 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME3 ;
 ANTENNADIFFAREA                          1.293 LAYER ME4 ;
END DO52
PIN DI51
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 209.238 0.000 209.558 0.600 ;
  LAYER ME3 ;
  RECT 209.238 0.000 209.558 0.600 ;
  LAYER ME2 ;
  RECT 209.238 0.000 209.558 0.600 ;
  LAYER ME1 ;
  RECT 209.238 0.000 209.558 0.600 ;
 END
 ANTENNAPARTIALMETALAREA                  1.058 LAYER ME2 ;
 ANTENNAGATEAREA                          0.072 LAYER ME2 ;
 ANTENNAGATEAREA                          0.072 LAYER ME3 ;
 ANTENNAGATEAREA                          0.072 LAYER ME4 ;
 ANTENNADIFFAREA                          0.160 LAYER ME2 ;
 ANTENNADIFFAREA                          0.160 LAYER ME3 ;
 ANTENNADIFFAREA                          0.160 LAYER ME4 ;
 ANTENNAMAXAREACAR                       21.782 LAYER ME2 ;
 ANTENNAMAXAREACAR                       24.449 LAYER ME3 ;
 ANTENNAMAXAREACAR                       27.116 LAYER ME4 ;
END DI51
PIN DO51
  DIRECTION OUTPUT ;
 PORT
  LAYER ME4 ;
  RECT 208.676 0.000 208.996 0.600 ;
  LAYER ME3 ;
  RECT 208.676 0.000 208.996 0.600 ;
  LAYER ME2 ;
  RECT 208.676 0.000 208.996 0.600 ;
  LAYER ME1 ;
  RECT 208.676 0.000 208.996 0.600 ;
 END
 ANTENNAPARTIALMETALAREA                  5.273 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME3 ;
 ANTENNADIFFAREA                          1.293 LAYER ME4 ;
END DO51
PIN DI50
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 205.234 0.000 205.554 0.600 ;
  LAYER ME3 ;
  RECT 205.234 0.000 205.554 0.600 ;
  LAYER ME2 ;
  RECT 205.234 0.000 205.554 0.600 ;
  LAYER ME1 ;
  RECT 205.234 0.000 205.554 0.600 ;
 END
 ANTENNAPARTIALMETALAREA                  1.058 LAYER ME2 ;
 ANTENNAGATEAREA                          0.072 LAYER ME2 ;
 ANTENNAGATEAREA                          0.072 LAYER ME3 ;
 ANTENNAGATEAREA                          0.072 LAYER ME4 ;
 ANTENNADIFFAREA                          0.160 LAYER ME2 ;
 ANTENNADIFFAREA                          0.160 LAYER ME3 ;
 ANTENNADIFFAREA                          0.160 LAYER ME4 ;
 ANTENNAMAXAREACAR                       21.782 LAYER ME2 ;
 ANTENNAMAXAREACAR                       24.449 LAYER ME3 ;
 ANTENNAMAXAREACAR                       27.116 LAYER ME4 ;
END DI50
PIN DO50
  DIRECTION OUTPUT ;
 PORT
  LAYER ME4 ;
  RECT 204.672 0.000 204.992 0.600 ;
  LAYER ME3 ;
  RECT 204.672 0.000 204.992 0.600 ;
  LAYER ME2 ;
  RECT 204.672 0.000 204.992 0.600 ;
  LAYER ME1 ;
  RECT 204.672 0.000 204.992 0.600 ;
 END
 ANTENNAPARTIALMETALAREA                  5.273 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME3 ;
 ANTENNADIFFAREA                          1.293 LAYER ME4 ;
END DO50
PIN DI49
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 201.230 0.000 201.550 0.600 ;
  LAYER ME3 ;
  RECT 201.230 0.000 201.550 0.600 ;
  LAYER ME2 ;
  RECT 201.230 0.000 201.550 0.600 ;
  LAYER ME1 ;
  RECT 201.230 0.000 201.550 0.600 ;
 END
 ANTENNAPARTIALMETALAREA                  1.058 LAYER ME2 ;
 ANTENNAGATEAREA                          0.072 LAYER ME2 ;
 ANTENNAGATEAREA                          0.072 LAYER ME3 ;
 ANTENNAGATEAREA                          0.072 LAYER ME4 ;
 ANTENNADIFFAREA                          0.160 LAYER ME2 ;
 ANTENNADIFFAREA                          0.160 LAYER ME3 ;
 ANTENNADIFFAREA                          0.160 LAYER ME4 ;
 ANTENNAMAXAREACAR                       21.782 LAYER ME2 ;
 ANTENNAMAXAREACAR                       24.449 LAYER ME3 ;
 ANTENNAMAXAREACAR                       27.116 LAYER ME4 ;
END DI49
PIN DO49
  DIRECTION OUTPUT ;
 PORT
  LAYER ME4 ;
  RECT 200.668 0.000 200.988 0.600 ;
  LAYER ME3 ;
  RECT 200.668 0.000 200.988 0.600 ;
  LAYER ME2 ;
  RECT 200.668 0.000 200.988 0.600 ;
  LAYER ME1 ;
  RECT 200.668 0.000 200.988 0.600 ;
 END
 ANTENNAPARTIALMETALAREA                  5.273 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME3 ;
 ANTENNADIFFAREA                          1.293 LAYER ME4 ;
END DO49
PIN DI48
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 196.664 0.000 196.984 0.600 ;
  LAYER ME3 ;
  RECT 196.664 0.000 196.984 0.600 ;
  LAYER ME2 ;
  RECT 196.664 0.000 196.984 0.600 ;
  LAYER ME1 ;
  RECT 196.664 0.000 196.984 0.600 ;
 END
 ANTENNAPARTIALMETALAREA                  0.346 LAYER ME1 ;
 ANTENNAPARTIALMETALAREA                  1.466 LAYER ME2 ;
 ANTENNAPARTIALMETALAREA                  0.508 LAYER ME3 ;
 ANTENNAGATEAREA                          0.072 LAYER ME3 ;
 ANTENNAGATEAREA                          0.072 LAYER ME4 ;
 ANTENNADIFFAREA                          0.218 LAYER ME1 ;
 ANTENNADIFFAREA                          0.218 LAYER ME2 ;
 ANTENNADIFFAREA                          0.218 LAYER ME3 ;
 ANTENNADIFFAREA                          0.218 LAYER ME4 ;
 ANTENNAMAXAREACAR                       17.267 LAYER ME3 ;
 ANTENNAMAXAREACAR                       19.933 LAYER ME4 ;
END DI48
PIN DO48
  DIRECTION OUTPUT ;
 PORT
  LAYER ME4 ;
  RECT 197.226 0.000 197.546 0.600 ;
  LAYER ME3 ;
  RECT 197.226 0.000 197.546 0.600 ;
  LAYER ME2 ;
  RECT 197.226 0.000 197.546 0.600 ;
  LAYER ME1 ;
  RECT 197.226 0.000 197.546 0.600 ;
 END
 ANTENNAPARTIALMETALAREA                  5.602 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME3 ;
 ANTENNADIFFAREA                          1.293 LAYER ME4 ;
END DO48
PIN WEB3
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 195.224 0.000 195.544 0.600 ;
  LAYER ME3 ;
  RECT 195.224 0.000 195.544 0.600 ;
  LAYER ME2 ;
  RECT 195.224 0.000 195.544 0.600 ;
  LAYER ME1 ;
  RECT 195.224 0.000 195.544 0.600 ;
 END
 ANTENNAPARTIALMETALAREA                  1.036 LAYER ME2 ;
 ANTENNAGATEAREA                          0.288 LAYER ME2 ;
 ANTENNAGATEAREA                          0.288 LAYER ME3 ;
 ANTENNAGATEAREA                          0.288 LAYER ME4 ;
 ANTENNADIFFAREA                          0.206 LAYER ME2 ;
 ANTENNADIFFAREA                          0.206 LAYER ME3 ;
 ANTENNADIFFAREA                          0.206 LAYER ME4 ;
 ANTENNAMAXAREACAR                        5.844 LAYER ME2 ;
 ANTENNAMAXAREACAR                        6.511 LAYER ME3 ;
 ANTENNAMAXAREACAR                        7.178 LAYER ME4 ;
END WEB3
PIN DI47
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 193.222 0.000 193.542 0.600 ;
  LAYER ME3 ;
  RECT 193.222 0.000 193.542 0.600 ;
  LAYER ME2 ;
  RECT 193.222 0.000 193.542 0.600 ;
  LAYER ME1 ;
  RECT 193.222 0.000 193.542 0.600 ;
 END
 ANTENNAPARTIALMETALAREA                  1.058 LAYER ME2 ;
 ANTENNAGATEAREA                          0.072 LAYER ME2 ;
 ANTENNAGATEAREA                          0.072 LAYER ME3 ;
 ANTENNAGATEAREA                          0.072 LAYER ME4 ;
 ANTENNADIFFAREA                          0.160 LAYER ME2 ;
 ANTENNADIFFAREA                          0.160 LAYER ME3 ;
 ANTENNADIFFAREA                          0.160 LAYER ME4 ;
 ANTENNAMAXAREACAR                       21.782 LAYER ME2 ;
 ANTENNAMAXAREACAR                       24.449 LAYER ME3 ;
 ANTENNAMAXAREACAR                       27.116 LAYER ME4 ;
END DI47
PIN DO47
  DIRECTION OUTPUT ;
 PORT
  LAYER ME4 ;
  RECT 192.660 0.000 192.980 0.600 ;
  LAYER ME3 ;
  RECT 192.660 0.000 192.980 0.600 ;
  LAYER ME2 ;
  RECT 192.660 0.000 192.980 0.600 ;
  LAYER ME1 ;
  RECT 192.660 0.000 192.980 0.600 ;
 END
 ANTENNAPARTIALMETALAREA                  5.273 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME3 ;
 ANTENNADIFFAREA                          1.293 LAYER ME4 ;
END DO47
PIN DI46
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 189.218 0.000 189.538 0.600 ;
  LAYER ME3 ;
  RECT 189.218 0.000 189.538 0.600 ;
  LAYER ME2 ;
  RECT 189.218 0.000 189.538 0.600 ;
  LAYER ME1 ;
  RECT 189.218 0.000 189.538 0.600 ;
 END
 ANTENNAPARTIALMETALAREA                  1.058 LAYER ME2 ;
 ANTENNAGATEAREA                          0.072 LAYER ME2 ;
 ANTENNAGATEAREA                          0.072 LAYER ME3 ;
 ANTENNAGATEAREA                          0.072 LAYER ME4 ;
 ANTENNADIFFAREA                          0.160 LAYER ME2 ;
 ANTENNADIFFAREA                          0.160 LAYER ME3 ;
 ANTENNADIFFAREA                          0.160 LAYER ME4 ;
 ANTENNAMAXAREACAR                       21.782 LAYER ME2 ;
 ANTENNAMAXAREACAR                       24.449 LAYER ME3 ;
 ANTENNAMAXAREACAR                       27.116 LAYER ME4 ;
END DI46
PIN DO46
  DIRECTION OUTPUT ;
 PORT
  LAYER ME4 ;
  RECT 188.656 0.000 188.976 0.600 ;
  LAYER ME3 ;
  RECT 188.656 0.000 188.976 0.600 ;
  LAYER ME2 ;
  RECT 188.656 0.000 188.976 0.600 ;
  LAYER ME1 ;
  RECT 188.656 0.000 188.976 0.600 ;
 END
 ANTENNAPARTIALMETALAREA                  5.273 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME3 ;
 ANTENNADIFFAREA                          1.293 LAYER ME4 ;
END DO46
PIN DI45
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 185.214 0.000 185.534 0.600 ;
  LAYER ME3 ;
  RECT 185.214 0.000 185.534 0.600 ;
  LAYER ME2 ;
  RECT 185.214 0.000 185.534 0.600 ;
  LAYER ME1 ;
  RECT 185.214 0.000 185.534 0.600 ;
 END
 ANTENNAPARTIALMETALAREA                  1.058 LAYER ME2 ;
 ANTENNAGATEAREA                          0.072 LAYER ME2 ;
 ANTENNAGATEAREA                          0.072 LAYER ME3 ;
 ANTENNAGATEAREA                          0.072 LAYER ME4 ;
 ANTENNADIFFAREA                          0.160 LAYER ME2 ;
 ANTENNADIFFAREA                          0.160 LAYER ME3 ;
 ANTENNADIFFAREA                          0.160 LAYER ME4 ;
 ANTENNAMAXAREACAR                       21.782 LAYER ME2 ;
 ANTENNAMAXAREACAR                       24.449 LAYER ME3 ;
 ANTENNAMAXAREACAR                       27.116 LAYER ME4 ;
END DI45
PIN DO45
  DIRECTION OUTPUT ;
 PORT
  LAYER ME4 ;
  RECT 184.652 0.000 184.972 0.600 ;
  LAYER ME3 ;
  RECT 184.652 0.000 184.972 0.600 ;
  LAYER ME2 ;
  RECT 184.652 0.000 184.972 0.600 ;
  LAYER ME1 ;
  RECT 184.652 0.000 184.972 0.600 ;
 END
 ANTENNAPARTIALMETALAREA                  5.273 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME3 ;
 ANTENNADIFFAREA                          1.293 LAYER ME4 ;
END DO45
PIN DI44
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 181.210 0.000 181.530 0.600 ;
  LAYER ME3 ;
  RECT 181.210 0.000 181.530 0.600 ;
  LAYER ME2 ;
  RECT 181.210 0.000 181.530 0.600 ;
  LAYER ME1 ;
  RECT 181.210 0.000 181.530 0.600 ;
 END
 ANTENNAPARTIALMETALAREA                  1.058 LAYER ME2 ;
 ANTENNAGATEAREA                          0.072 LAYER ME2 ;
 ANTENNAGATEAREA                          0.072 LAYER ME3 ;
 ANTENNAGATEAREA                          0.072 LAYER ME4 ;
 ANTENNADIFFAREA                          0.160 LAYER ME2 ;
 ANTENNADIFFAREA                          0.160 LAYER ME3 ;
 ANTENNADIFFAREA                          0.160 LAYER ME4 ;
 ANTENNAMAXAREACAR                       21.782 LAYER ME2 ;
 ANTENNAMAXAREACAR                       24.449 LAYER ME3 ;
 ANTENNAMAXAREACAR                       27.116 LAYER ME4 ;
END DI44
PIN DO44
  DIRECTION OUTPUT ;
 PORT
  LAYER ME4 ;
  RECT 180.648 0.000 180.968 0.600 ;
  LAYER ME3 ;
  RECT 180.648 0.000 180.968 0.600 ;
  LAYER ME2 ;
  RECT 180.648 0.000 180.968 0.600 ;
  LAYER ME1 ;
  RECT 180.648 0.000 180.968 0.600 ;
 END
 ANTENNAPARTIALMETALAREA                  5.273 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME3 ;
 ANTENNADIFFAREA                          1.293 LAYER ME4 ;
END DO44
PIN DI43
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 177.206 0.000 177.526 0.600 ;
  LAYER ME3 ;
  RECT 177.206 0.000 177.526 0.600 ;
  LAYER ME2 ;
  RECT 177.206 0.000 177.526 0.600 ;
  LAYER ME1 ;
  RECT 177.206 0.000 177.526 0.600 ;
 END
 ANTENNAPARTIALMETALAREA                  1.058 LAYER ME2 ;
 ANTENNAGATEAREA                          0.072 LAYER ME2 ;
 ANTENNAGATEAREA                          0.072 LAYER ME3 ;
 ANTENNAGATEAREA                          0.072 LAYER ME4 ;
 ANTENNADIFFAREA                          0.160 LAYER ME2 ;
 ANTENNADIFFAREA                          0.160 LAYER ME3 ;
 ANTENNADIFFAREA                          0.160 LAYER ME4 ;
 ANTENNAMAXAREACAR                       21.782 LAYER ME2 ;
 ANTENNAMAXAREACAR                       24.449 LAYER ME3 ;
 ANTENNAMAXAREACAR                       27.116 LAYER ME4 ;
END DI43
PIN DO43
  DIRECTION OUTPUT ;
 PORT
  LAYER ME4 ;
  RECT 176.644 0.000 176.964 0.600 ;
  LAYER ME3 ;
  RECT 176.644 0.000 176.964 0.600 ;
  LAYER ME2 ;
  RECT 176.644 0.000 176.964 0.600 ;
  LAYER ME1 ;
  RECT 176.644 0.000 176.964 0.600 ;
 END
 ANTENNAPARTIALMETALAREA                  5.273 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME3 ;
 ANTENNADIFFAREA                          1.293 LAYER ME4 ;
END DO43
PIN DI42
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 173.202 0.000 173.522 0.600 ;
  LAYER ME3 ;
  RECT 173.202 0.000 173.522 0.600 ;
  LAYER ME2 ;
  RECT 173.202 0.000 173.522 0.600 ;
  LAYER ME1 ;
  RECT 173.202 0.000 173.522 0.600 ;
 END
 ANTENNAPARTIALMETALAREA                  1.058 LAYER ME2 ;
 ANTENNAGATEAREA                          0.072 LAYER ME2 ;
 ANTENNAGATEAREA                          0.072 LAYER ME3 ;
 ANTENNAGATEAREA                          0.072 LAYER ME4 ;
 ANTENNADIFFAREA                          0.160 LAYER ME2 ;
 ANTENNADIFFAREA                          0.160 LAYER ME3 ;
 ANTENNADIFFAREA                          0.160 LAYER ME4 ;
 ANTENNAMAXAREACAR                       21.782 LAYER ME2 ;
 ANTENNAMAXAREACAR                       24.449 LAYER ME3 ;
 ANTENNAMAXAREACAR                       27.116 LAYER ME4 ;
END DI42
PIN DO42
  DIRECTION OUTPUT ;
 PORT
  LAYER ME4 ;
  RECT 172.640 0.000 172.960 0.600 ;
  LAYER ME3 ;
  RECT 172.640 0.000 172.960 0.600 ;
  LAYER ME2 ;
  RECT 172.640 0.000 172.960 0.600 ;
  LAYER ME1 ;
  RECT 172.640 0.000 172.960 0.600 ;
 END
 ANTENNAPARTIALMETALAREA                  5.273 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME3 ;
 ANTENNADIFFAREA                          1.293 LAYER ME4 ;
END DO42
PIN DI41
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 169.198 0.000 169.518 0.600 ;
  LAYER ME3 ;
  RECT 169.198 0.000 169.518 0.600 ;
  LAYER ME2 ;
  RECT 169.198 0.000 169.518 0.600 ;
  LAYER ME1 ;
  RECT 169.198 0.000 169.518 0.600 ;
 END
 ANTENNAPARTIALMETALAREA                  1.058 LAYER ME2 ;
 ANTENNAGATEAREA                          0.072 LAYER ME2 ;
 ANTENNAGATEAREA                          0.072 LAYER ME3 ;
 ANTENNAGATEAREA                          0.072 LAYER ME4 ;
 ANTENNADIFFAREA                          0.160 LAYER ME2 ;
 ANTENNADIFFAREA                          0.160 LAYER ME3 ;
 ANTENNADIFFAREA                          0.160 LAYER ME4 ;
 ANTENNAMAXAREACAR                       21.782 LAYER ME2 ;
 ANTENNAMAXAREACAR                       24.449 LAYER ME3 ;
 ANTENNAMAXAREACAR                       27.116 LAYER ME4 ;
END DI41
PIN DO41
  DIRECTION OUTPUT ;
 PORT
  LAYER ME4 ;
  RECT 168.636 0.000 168.956 0.600 ;
  LAYER ME3 ;
  RECT 168.636 0.000 168.956 0.600 ;
  LAYER ME2 ;
  RECT 168.636 0.000 168.956 0.600 ;
  LAYER ME1 ;
  RECT 168.636 0.000 168.956 0.600 ;
 END
 ANTENNAPARTIALMETALAREA                  5.273 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME3 ;
 ANTENNADIFFAREA                          1.293 LAYER ME4 ;
END DO41
PIN DI40
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 165.194 0.000 165.514 0.600 ;
  LAYER ME3 ;
  RECT 165.194 0.000 165.514 0.600 ;
  LAYER ME2 ;
  RECT 165.194 0.000 165.514 0.600 ;
  LAYER ME1 ;
  RECT 165.194 0.000 165.514 0.600 ;
 END
 ANTENNAPARTIALMETALAREA                  1.058 LAYER ME2 ;
 ANTENNAGATEAREA                          0.072 LAYER ME2 ;
 ANTENNAGATEAREA                          0.072 LAYER ME3 ;
 ANTENNAGATEAREA                          0.072 LAYER ME4 ;
 ANTENNADIFFAREA                          0.160 LAYER ME2 ;
 ANTENNADIFFAREA                          0.160 LAYER ME3 ;
 ANTENNADIFFAREA                          0.160 LAYER ME4 ;
 ANTENNAMAXAREACAR                       21.782 LAYER ME2 ;
 ANTENNAMAXAREACAR                       24.449 LAYER ME3 ;
 ANTENNAMAXAREACAR                       27.116 LAYER ME4 ;
END DI40
PIN DO40
  DIRECTION OUTPUT ;
 PORT
  LAYER ME4 ;
  RECT 164.632 0.000 164.952 0.600 ;
  LAYER ME3 ;
  RECT 164.632 0.000 164.952 0.600 ;
  LAYER ME2 ;
  RECT 164.632 0.000 164.952 0.600 ;
  LAYER ME1 ;
  RECT 164.632 0.000 164.952 0.600 ;
 END
 ANTENNAPARTIALMETALAREA                  5.273 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME3 ;
 ANTENNADIFFAREA                          1.293 LAYER ME4 ;
END DO40
PIN DI39
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 161.190 0.000 161.510 0.600 ;
  LAYER ME3 ;
  RECT 161.190 0.000 161.510 0.600 ;
  LAYER ME2 ;
  RECT 161.190 0.000 161.510 0.600 ;
  LAYER ME1 ;
  RECT 161.190 0.000 161.510 0.600 ;
 END
 ANTENNAPARTIALMETALAREA                  1.058 LAYER ME2 ;
 ANTENNAGATEAREA                          0.072 LAYER ME2 ;
 ANTENNAGATEAREA                          0.072 LAYER ME3 ;
 ANTENNAGATEAREA                          0.072 LAYER ME4 ;
 ANTENNADIFFAREA                          0.160 LAYER ME2 ;
 ANTENNADIFFAREA                          0.160 LAYER ME3 ;
 ANTENNADIFFAREA                          0.160 LAYER ME4 ;
 ANTENNAMAXAREACAR                       21.782 LAYER ME2 ;
 ANTENNAMAXAREACAR                       24.449 LAYER ME3 ;
 ANTENNAMAXAREACAR                       27.116 LAYER ME4 ;
END DI39
PIN DO39
  DIRECTION OUTPUT ;
 PORT
  LAYER ME4 ;
  RECT 160.628 0.000 160.948 0.600 ;
  LAYER ME3 ;
  RECT 160.628 0.000 160.948 0.600 ;
  LAYER ME2 ;
  RECT 160.628 0.000 160.948 0.600 ;
  LAYER ME1 ;
  RECT 160.628 0.000 160.948 0.600 ;
 END
 ANTENNAPARTIALMETALAREA                  5.273 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME3 ;
 ANTENNADIFFAREA                          1.293 LAYER ME4 ;
END DO39
PIN DI38
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 157.186 0.000 157.506 0.600 ;
  LAYER ME3 ;
  RECT 157.186 0.000 157.506 0.600 ;
  LAYER ME2 ;
  RECT 157.186 0.000 157.506 0.600 ;
  LAYER ME1 ;
  RECT 157.186 0.000 157.506 0.600 ;
 END
 ANTENNAPARTIALMETALAREA                  1.058 LAYER ME2 ;
 ANTENNAGATEAREA                          0.072 LAYER ME2 ;
 ANTENNAGATEAREA                          0.072 LAYER ME3 ;
 ANTENNAGATEAREA                          0.072 LAYER ME4 ;
 ANTENNADIFFAREA                          0.160 LAYER ME2 ;
 ANTENNADIFFAREA                          0.160 LAYER ME3 ;
 ANTENNADIFFAREA                          0.160 LAYER ME4 ;
 ANTENNAMAXAREACAR                       21.782 LAYER ME2 ;
 ANTENNAMAXAREACAR                       24.449 LAYER ME3 ;
 ANTENNAMAXAREACAR                       27.116 LAYER ME4 ;
END DI38
PIN DO38
  DIRECTION OUTPUT ;
 PORT
  LAYER ME4 ;
  RECT 156.624 0.000 156.944 0.600 ;
  LAYER ME3 ;
  RECT 156.624 0.000 156.944 0.600 ;
  LAYER ME2 ;
  RECT 156.624 0.000 156.944 0.600 ;
  LAYER ME1 ;
  RECT 156.624 0.000 156.944 0.600 ;
 END
 ANTENNAPARTIALMETALAREA                  5.273 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME3 ;
 ANTENNADIFFAREA                          1.293 LAYER ME4 ;
END DO38
PIN DI37
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 153.182 0.000 153.502 0.600 ;
  LAYER ME3 ;
  RECT 153.182 0.000 153.502 0.600 ;
  LAYER ME2 ;
  RECT 153.182 0.000 153.502 0.600 ;
  LAYER ME1 ;
  RECT 153.182 0.000 153.502 0.600 ;
 END
 ANTENNAPARTIALMETALAREA                  1.058 LAYER ME2 ;
 ANTENNAGATEAREA                          0.072 LAYER ME2 ;
 ANTENNAGATEAREA                          0.072 LAYER ME3 ;
 ANTENNAGATEAREA                          0.072 LAYER ME4 ;
 ANTENNADIFFAREA                          0.160 LAYER ME2 ;
 ANTENNADIFFAREA                          0.160 LAYER ME3 ;
 ANTENNADIFFAREA                          0.160 LAYER ME4 ;
 ANTENNAMAXAREACAR                       21.782 LAYER ME2 ;
 ANTENNAMAXAREACAR                       24.449 LAYER ME3 ;
 ANTENNAMAXAREACAR                       27.116 LAYER ME4 ;
END DI37
PIN DO37
  DIRECTION OUTPUT ;
 PORT
  LAYER ME4 ;
  RECT 152.620 0.000 152.940 0.600 ;
  LAYER ME3 ;
  RECT 152.620 0.000 152.940 0.600 ;
  LAYER ME2 ;
  RECT 152.620 0.000 152.940 0.600 ;
  LAYER ME1 ;
  RECT 152.620 0.000 152.940 0.600 ;
 END
 ANTENNAPARTIALMETALAREA                  5.273 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME3 ;
 ANTENNADIFFAREA                          1.293 LAYER ME4 ;
END DO37
PIN DI36
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 149.178 0.000 149.498 0.600 ;
  LAYER ME3 ;
  RECT 149.178 0.000 149.498 0.600 ;
  LAYER ME2 ;
  RECT 149.178 0.000 149.498 0.600 ;
  LAYER ME1 ;
  RECT 149.178 0.000 149.498 0.600 ;
 END
 ANTENNAPARTIALMETALAREA                  1.058 LAYER ME2 ;
 ANTENNAGATEAREA                          0.072 LAYER ME2 ;
 ANTENNAGATEAREA                          0.072 LAYER ME3 ;
 ANTENNAGATEAREA                          0.072 LAYER ME4 ;
 ANTENNADIFFAREA                          0.160 LAYER ME2 ;
 ANTENNADIFFAREA                          0.160 LAYER ME3 ;
 ANTENNADIFFAREA                          0.160 LAYER ME4 ;
 ANTENNAMAXAREACAR                       21.782 LAYER ME2 ;
 ANTENNAMAXAREACAR                       24.449 LAYER ME3 ;
 ANTENNAMAXAREACAR                       27.116 LAYER ME4 ;
END DI36
PIN DO36
  DIRECTION OUTPUT ;
 PORT
  LAYER ME4 ;
  RECT 148.616 0.000 148.936 0.600 ;
  LAYER ME3 ;
  RECT 148.616 0.000 148.936 0.600 ;
  LAYER ME2 ;
  RECT 148.616 0.000 148.936 0.600 ;
  LAYER ME1 ;
  RECT 148.616 0.000 148.936 0.600 ;
 END
 ANTENNAPARTIALMETALAREA                  5.273 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME3 ;
 ANTENNADIFFAREA                          1.293 LAYER ME4 ;
END DO36
PIN DI35
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 145.174 0.000 145.494 0.600 ;
  LAYER ME3 ;
  RECT 145.174 0.000 145.494 0.600 ;
  LAYER ME2 ;
  RECT 145.174 0.000 145.494 0.600 ;
  LAYER ME1 ;
  RECT 145.174 0.000 145.494 0.600 ;
 END
 ANTENNAPARTIALMETALAREA                  1.058 LAYER ME2 ;
 ANTENNAGATEAREA                          0.072 LAYER ME2 ;
 ANTENNAGATEAREA                          0.072 LAYER ME3 ;
 ANTENNAGATEAREA                          0.072 LAYER ME4 ;
 ANTENNADIFFAREA                          0.160 LAYER ME2 ;
 ANTENNADIFFAREA                          0.160 LAYER ME3 ;
 ANTENNADIFFAREA                          0.160 LAYER ME4 ;
 ANTENNAMAXAREACAR                       21.782 LAYER ME2 ;
 ANTENNAMAXAREACAR                       24.449 LAYER ME3 ;
 ANTENNAMAXAREACAR                       27.116 LAYER ME4 ;
END DI35
PIN DO35
  DIRECTION OUTPUT ;
 PORT
  LAYER ME4 ;
  RECT 144.612 0.000 144.932 0.600 ;
  LAYER ME3 ;
  RECT 144.612 0.000 144.932 0.600 ;
  LAYER ME2 ;
  RECT 144.612 0.000 144.932 0.600 ;
  LAYER ME1 ;
  RECT 144.612 0.000 144.932 0.600 ;
 END
 ANTENNAPARTIALMETALAREA                  5.273 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME3 ;
 ANTENNADIFFAREA                          1.293 LAYER ME4 ;
END DO35
PIN DI34
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 141.170 0.000 141.490 0.600 ;
  LAYER ME3 ;
  RECT 141.170 0.000 141.490 0.600 ;
  LAYER ME2 ;
  RECT 141.170 0.000 141.490 0.600 ;
  LAYER ME1 ;
  RECT 141.170 0.000 141.490 0.600 ;
 END
 ANTENNAPARTIALMETALAREA                  1.058 LAYER ME2 ;
 ANTENNAGATEAREA                          0.072 LAYER ME2 ;
 ANTENNAGATEAREA                          0.072 LAYER ME3 ;
 ANTENNAGATEAREA                          0.072 LAYER ME4 ;
 ANTENNADIFFAREA                          0.160 LAYER ME2 ;
 ANTENNADIFFAREA                          0.160 LAYER ME3 ;
 ANTENNADIFFAREA                          0.160 LAYER ME4 ;
 ANTENNAMAXAREACAR                       21.782 LAYER ME2 ;
 ANTENNAMAXAREACAR                       24.449 LAYER ME3 ;
 ANTENNAMAXAREACAR                       27.116 LAYER ME4 ;
END DI34
PIN DO34
  DIRECTION OUTPUT ;
 PORT
  LAYER ME4 ;
  RECT 140.608 0.000 140.928 0.600 ;
  LAYER ME3 ;
  RECT 140.608 0.000 140.928 0.600 ;
  LAYER ME2 ;
  RECT 140.608 0.000 140.928 0.600 ;
  LAYER ME1 ;
  RECT 140.608 0.000 140.928 0.600 ;
 END
 ANTENNAPARTIALMETALAREA                  5.273 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME3 ;
 ANTENNADIFFAREA                          1.293 LAYER ME4 ;
END DO34
PIN DI33
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 137.166 0.000 137.486 0.600 ;
  LAYER ME3 ;
  RECT 137.166 0.000 137.486 0.600 ;
  LAYER ME2 ;
  RECT 137.166 0.000 137.486 0.600 ;
  LAYER ME1 ;
  RECT 137.166 0.000 137.486 0.600 ;
 END
 ANTENNAPARTIALMETALAREA                  1.058 LAYER ME2 ;
 ANTENNAGATEAREA                          0.072 LAYER ME2 ;
 ANTENNAGATEAREA                          0.072 LAYER ME3 ;
 ANTENNAGATEAREA                          0.072 LAYER ME4 ;
 ANTENNADIFFAREA                          0.160 LAYER ME2 ;
 ANTENNADIFFAREA                          0.160 LAYER ME3 ;
 ANTENNADIFFAREA                          0.160 LAYER ME4 ;
 ANTENNAMAXAREACAR                       21.782 LAYER ME2 ;
 ANTENNAMAXAREACAR                       24.449 LAYER ME3 ;
 ANTENNAMAXAREACAR                       27.116 LAYER ME4 ;
END DI33
PIN DO33
  DIRECTION OUTPUT ;
 PORT
  LAYER ME4 ;
  RECT 136.604 0.000 136.924 0.600 ;
  LAYER ME3 ;
  RECT 136.604 0.000 136.924 0.600 ;
  LAYER ME2 ;
  RECT 136.604 0.000 136.924 0.600 ;
  LAYER ME1 ;
  RECT 136.604 0.000 136.924 0.600 ;
 END
 ANTENNAPARTIALMETALAREA                  5.273 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME3 ;
 ANTENNADIFFAREA                          1.293 LAYER ME4 ;
END DO33
PIN DI32
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 132.600 0.000 132.920 0.600 ;
  LAYER ME3 ;
  RECT 132.600 0.000 132.920 0.600 ;
  LAYER ME2 ;
  RECT 132.600 0.000 132.920 0.600 ;
  LAYER ME1 ;
  RECT 132.600 0.000 132.920 0.600 ;
 END
 ANTENNAPARTIALMETALAREA                  0.346 LAYER ME1 ;
 ANTENNAPARTIALMETALAREA                  1.466 LAYER ME2 ;
 ANTENNAPARTIALMETALAREA                  0.508 LAYER ME3 ;
 ANTENNAGATEAREA                          0.072 LAYER ME3 ;
 ANTENNAGATEAREA                          0.072 LAYER ME4 ;
 ANTENNADIFFAREA                          0.218 LAYER ME1 ;
 ANTENNADIFFAREA                          0.218 LAYER ME2 ;
 ANTENNADIFFAREA                          0.218 LAYER ME3 ;
 ANTENNADIFFAREA                          0.218 LAYER ME4 ;
 ANTENNAMAXAREACAR                       17.267 LAYER ME3 ;
 ANTENNAMAXAREACAR                       19.933 LAYER ME4 ;
END DI32
PIN DO32
  DIRECTION OUTPUT ;
 PORT
  LAYER ME4 ;
  RECT 133.162 0.000 133.482 0.600 ;
  LAYER ME3 ;
  RECT 133.162 0.000 133.482 0.600 ;
  LAYER ME2 ;
  RECT 133.162 0.000 133.482 0.600 ;
  LAYER ME1 ;
  RECT 133.162 0.000 133.482 0.600 ;
 END
 ANTENNAPARTIALMETALAREA                  5.602 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME3 ;
 ANTENNADIFFAREA                          1.293 LAYER ME4 ;
END DO32
PIN WEB2
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 131.160 0.000 131.480 0.600 ;
  LAYER ME3 ;
  RECT 131.160 0.000 131.480 0.600 ;
  LAYER ME2 ;
  RECT 131.160 0.000 131.480 0.600 ;
  LAYER ME1 ;
  RECT 131.160 0.000 131.480 0.600 ;
 END
 ANTENNAPARTIALMETALAREA                  1.036 LAYER ME2 ;
 ANTENNAGATEAREA                          0.288 LAYER ME2 ;
 ANTENNAGATEAREA                          0.288 LAYER ME3 ;
 ANTENNAGATEAREA                          0.288 LAYER ME4 ;
 ANTENNADIFFAREA                          0.206 LAYER ME2 ;
 ANTENNADIFFAREA                          0.206 LAYER ME3 ;
 ANTENNADIFFAREA                          0.206 LAYER ME4 ;
 ANTENNAMAXAREACAR                        5.844 LAYER ME2 ;
 ANTENNAMAXAREACAR                        6.511 LAYER ME3 ;
 ANTENNAMAXAREACAR                        7.178 LAYER ME4 ;
END WEB2
PIN DI31
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 129.158 0.000 129.478 0.600 ;
  LAYER ME3 ;
  RECT 129.158 0.000 129.478 0.600 ;
  LAYER ME2 ;
  RECT 129.158 0.000 129.478 0.600 ;
  LAYER ME1 ;
  RECT 129.158 0.000 129.478 0.600 ;
 END
 ANTENNAPARTIALMETALAREA                  1.058 LAYER ME2 ;
 ANTENNAGATEAREA                          0.072 LAYER ME2 ;
 ANTENNAGATEAREA                          0.072 LAYER ME3 ;
 ANTENNAGATEAREA                          0.072 LAYER ME4 ;
 ANTENNADIFFAREA                          0.160 LAYER ME2 ;
 ANTENNADIFFAREA                          0.160 LAYER ME3 ;
 ANTENNADIFFAREA                          0.160 LAYER ME4 ;
 ANTENNAMAXAREACAR                       21.782 LAYER ME2 ;
 ANTENNAMAXAREACAR                       24.449 LAYER ME3 ;
 ANTENNAMAXAREACAR                       27.116 LAYER ME4 ;
END DI31
PIN DO31
  DIRECTION OUTPUT ;
 PORT
  LAYER ME4 ;
  RECT 128.596 0.000 128.916 0.600 ;
  LAYER ME3 ;
  RECT 128.596 0.000 128.916 0.600 ;
  LAYER ME2 ;
  RECT 128.596 0.000 128.916 0.600 ;
  LAYER ME1 ;
  RECT 128.596 0.000 128.916 0.600 ;
 END
 ANTENNAPARTIALMETALAREA                  5.273 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME3 ;
 ANTENNADIFFAREA                          1.293 LAYER ME4 ;
END DO31
PIN DI30
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 125.154 0.000 125.474 0.600 ;
  LAYER ME3 ;
  RECT 125.154 0.000 125.474 0.600 ;
  LAYER ME2 ;
  RECT 125.154 0.000 125.474 0.600 ;
  LAYER ME1 ;
  RECT 125.154 0.000 125.474 0.600 ;
 END
 ANTENNAPARTIALMETALAREA                  1.058 LAYER ME2 ;
 ANTENNAGATEAREA                          0.072 LAYER ME2 ;
 ANTENNAGATEAREA                          0.072 LAYER ME3 ;
 ANTENNAGATEAREA                          0.072 LAYER ME4 ;
 ANTENNADIFFAREA                          0.160 LAYER ME2 ;
 ANTENNADIFFAREA                          0.160 LAYER ME3 ;
 ANTENNADIFFAREA                          0.160 LAYER ME4 ;
 ANTENNAMAXAREACAR                       21.782 LAYER ME2 ;
 ANTENNAMAXAREACAR                       24.449 LAYER ME3 ;
 ANTENNAMAXAREACAR                       27.116 LAYER ME4 ;
END DI30
PIN DO30
  DIRECTION OUTPUT ;
 PORT
  LAYER ME4 ;
  RECT 124.592 0.000 124.912 0.600 ;
  LAYER ME3 ;
  RECT 124.592 0.000 124.912 0.600 ;
  LAYER ME2 ;
  RECT 124.592 0.000 124.912 0.600 ;
  LAYER ME1 ;
  RECT 124.592 0.000 124.912 0.600 ;
 END
 ANTENNAPARTIALMETALAREA                  5.273 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME3 ;
 ANTENNADIFFAREA                          1.293 LAYER ME4 ;
END DO30
PIN DI29
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 121.150 0.000 121.470 0.600 ;
  LAYER ME3 ;
  RECT 121.150 0.000 121.470 0.600 ;
  LAYER ME2 ;
  RECT 121.150 0.000 121.470 0.600 ;
  LAYER ME1 ;
  RECT 121.150 0.000 121.470 0.600 ;
 END
 ANTENNAPARTIALMETALAREA                  1.058 LAYER ME2 ;
 ANTENNAGATEAREA                          0.072 LAYER ME2 ;
 ANTENNAGATEAREA                          0.072 LAYER ME3 ;
 ANTENNAGATEAREA                          0.072 LAYER ME4 ;
 ANTENNADIFFAREA                          0.160 LAYER ME2 ;
 ANTENNADIFFAREA                          0.160 LAYER ME3 ;
 ANTENNADIFFAREA                          0.160 LAYER ME4 ;
 ANTENNAMAXAREACAR                       21.782 LAYER ME2 ;
 ANTENNAMAXAREACAR                       24.449 LAYER ME3 ;
 ANTENNAMAXAREACAR                       27.116 LAYER ME4 ;
END DI29
PIN DO29
  DIRECTION OUTPUT ;
 PORT
  LAYER ME4 ;
  RECT 120.588 0.000 120.908 0.600 ;
  LAYER ME3 ;
  RECT 120.588 0.000 120.908 0.600 ;
  LAYER ME2 ;
  RECT 120.588 0.000 120.908 0.600 ;
  LAYER ME1 ;
  RECT 120.588 0.000 120.908 0.600 ;
 END
 ANTENNAPARTIALMETALAREA                  5.273 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME3 ;
 ANTENNADIFFAREA                          1.293 LAYER ME4 ;
END DO29
PIN DI28
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 117.146 0.000 117.466 0.600 ;
  LAYER ME3 ;
  RECT 117.146 0.000 117.466 0.600 ;
  LAYER ME2 ;
  RECT 117.146 0.000 117.466 0.600 ;
  LAYER ME1 ;
  RECT 117.146 0.000 117.466 0.600 ;
 END
 ANTENNAPARTIALMETALAREA                  1.058 LAYER ME2 ;
 ANTENNAGATEAREA                          0.072 LAYER ME2 ;
 ANTENNAGATEAREA                          0.072 LAYER ME3 ;
 ANTENNAGATEAREA                          0.072 LAYER ME4 ;
 ANTENNADIFFAREA                          0.160 LAYER ME2 ;
 ANTENNADIFFAREA                          0.160 LAYER ME3 ;
 ANTENNADIFFAREA                          0.160 LAYER ME4 ;
 ANTENNAMAXAREACAR                       21.782 LAYER ME2 ;
 ANTENNAMAXAREACAR                       24.449 LAYER ME3 ;
 ANTENNAMAXAREACAR                       27.116 LAYER ME4 ;
END DI28
PIN DO28
  DIRECTION OUTPUT ;
 PORT
  LAYER ME4 ;
  RECT 116.584 0.000 116.904 0.600 ;
  LAYER ME3 ;
  RECT 116.584 0.000 116.904 0.600 ;
  LAYER ME2 ;
  RECT 116.584 0.000 116.904 0.600 ;
  LAYER ME1 ;
  RECT 116.584 0.000 116.904 0.600 ;
 END
 ANTENNAPARTIALMETALAREA                  5.273 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME3 ;
 ANTENNADIFFAREA                          1.293 LAYER ME4 ;
END DO28
PIN DI27
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 113.142 0.000 113.462 0.600 ;
  LAYER ME3 ;
  RECT 113.142 0.000 113.462 0.600 ;
  LAYER ME2 ;
  RECT 113.142 0.000 113.462 0.600 ;
  LAYER ME1 ;
  RECT 113.142 0.000 113.462 0.600 ;
 END
 ANTENNAPARTIALMETALAREA                  1.058 LAYER ME2 ;
 ANTENNAGATEAREA                          0.072 LAYER ME2 ;
 ANTENNAGATEAREA                          0.072 LAYER ME3 ;
 ANTENNAGATEAREA                          0.072 LAYER ME4 ;
 ANTENNADIFFAREA                          0.160 LAYER ME2 ;
 ANTENNADIFFAREA                          0.160 LAYER ME3 ;
 ANTENNADIFFAREA                          0.160 LAYER ME4 ;
 ANTENNAMAXAREACAR                       21.782 LAYER ME2 ;
 ANTENNAMAXAREACAR                       24.449 LAYER ME3 ;
 ANTENNAMAXAREACAR                       27.116 LAYER ME4 ;
END DI27
PIN DO27
  DIRECTION OUTPUT ;
 PORT
  LAYER ME4 ;
  RECT 112.580 0.000 112.900 0.600 ;
  LAYER ME3 ;
  RECT 112.580 0.000 112.900 0.600 ;
  LAYER ME2 ;
  RECT 112.580 0.000 112.900 0.600 ;
  LAYER ME1 ;
  RECT 112.580 0.000 112.900 0.600 ;
 END
 ANTENNAPARTIALMETALAREA                  5.273 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME3 ;
 ANTENNADIFFAREA                          1.293 LAYER ME4 ;
END DO27
PIN DI26
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 109.138 0.000 109.458 0.600 ;
  LAYER ME3 ;
  RECT 109.138 0.000 109.458 0.600 ;
  LAYER ME2 ;
  RECT 109.138 0.000 109.458 0.600 ;
  LAYER ME1 ;
  RECT 109.138 0.000 109.458 0.600 ;
 END
 ANTENNAPARTIALMETALAREA                  1.058 LAYER ME2 ;
 ANTENNAGATEAREA                          0.072 LAYER ME2 ;
 ANTENNAGATEAREA                          0.072 LAYER ME3 ;
 ANTENNAGATEAREA                          0.072 LAYER ME4 ;
 ANTENNADIFFAREA                          0.160 LAYER ME2 ;
 ANTENNADIFFAREA                          0.160 LAYER ME3 ;
 ANTENNADIFFAREA                          0.160 LAYER ME4 ;
 ANTENNAMAXAREACAR                       21.782 LAYER ME2 ;
 ANTENNAMAXAREACAR                       24.449 LAYER ME3 ;
 ANTENNAMAXAREACAR                       27.116 LAYER ME4 ;
END DI26
PIN DO26
  DIRECTION OUTPUT ;
 PORT
  LAYER ME4 ;
  RECT 108.576 0.000 108.896 0.600 ;
  LAYER ME3 ;
  RECT 108.576 0.000 108.896 0.600 ;
  LAYER ME2 ;
  RECT 108.576 0.000 108.896 0.600 ;
  LAYER ME1 ;
  RECT 108.576 0.000 108.896 0.600 ;
 END
 ANTENNAPARTIALMETALAREA                  5.273 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME3 ;
 ANTENNADIFFAREA                          1.293 LAYER ME4 ;
END DO26
PIN DI25
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 105.134 0.000 105.454 0.600 ;
  LAYER ME3 ;
  RECT 105.134 0.000 105.454 0.600 ;
  LAYER ME2 ;
  RECT 105.134 0.000 105.454 0.600 ;
  LAYER ME1 ;
  RECT 105.134 0.000 105.454 0.600 ;
 END
 ANTENNAPARTIALMETALAREA                  1.058 LAYER ME2 ;
 ANTENNAGATEAREA                          0.072 LAYER ME2 ;
 ANTENNAGATEAREA                          0.072 LAYER ME3 ;
 ANTENNAGATEAREA                          0.072 LAYER ME4 ;
 ANTENNADIFFAREA                          0.160 LAYER ME2 ;
 ANTENNADIFFAREA                          0.160 LAYER ME3 ;
 ANTENNADIFFAREA                          0.160 LAYER ME4 ;
 ANTENNAMAXAREACAR                       21.782 LAYER ME2 ;
 ANTENNAMAXAREACAR                       24.449 LAYER ME3 ;
 ANTENNAMAXAREACAR                       27.116 LAYER ME4 ;
END DI25
PIN DO25
  DIRECTION OUTPUT ;
 PORT
  LAYER ME4 ;
  RECT 104.572 0.000 104.892 0.600 ;
  LAYER ME3 ;
  RECT 104.572 0.000 104.892 0.600 ;
  LAYER ME2 ;
  RECT 104.572 0.000 104.892 0.600 ;
  LAYER ME1 ;
  RECT 104.572 0.000 104.892 0.600 ;
 END
 ANTENNAPARTIALMETALAREA                  5.273 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME3 ;
 ANTENNADIFFAREA                          1.293 LAYER ME4 ;
END DO25
PIN DI24
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 101.130 0.000 101.450 0.600 ;
  LAYER ME3 ;
  RECT 101.130 0.000 101.450 0.600 ;
  LAYER ME2 ;
  RECT 101.130 0.000 101.450 0.600 ;
  LAYER ME1 ;
  RECT 101.130 0.000 101.450 0.600 ;
 END
 ANTENNAPARTIALMETALAREA                  1.058 LAYER ME2 ;
 ANTENNAGATEAREA                          0.072 LAYER ME2 ;
 ANTENNAGATEAREA                          0.072 LAYER ME3 ;
 ANTENNAGATEAREA                          0.072 LAYER ME4 ;
 ANTENNADIFFAREA                          0.160 LAYER ME2 ;
 ANTENNADIFFAREA                          0.160 LAYER ME3 ;
 ANTENNADIFFAREA                          0.160 LAYER ME4 ;
 ANTENNAMAXAREACAR                       21.782 LAYER ME2 ;
 ANTENNAMAXAREACAR                       24.449 LAYER ME3 ;
 ANTENNAMAXAREACAR                       27.116 LAYER ME4 ;
END DI24
PIN DO24
  DIRECTION OUTPUT ;
 PORT
  LAYER ME4 ;
  RECT 100.568 0.000 100.888 0.600 ;
  LAYER ME3 ;
  RECT 100.568 0.000 100.888 0.600 ;
  LAYER ME2 ;
  RECT 100.568 0.000 100.888 0.600 ;
  LAYER ME1 ;
  RECT 100.568 0.000 100.888 0.600 ;
 END
 ANTENNAPARTIALMETALAREA                  5.273 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME3 ;
 ANTENNADIFFAREA                          1.293 LAYER ME4 ;
END DO24
PIN DI23
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 97.126 0.000 97.446 0.600 ;
  LAYER ME3 ;
  RECT 97.126 0.000 97.446 0.600 ;
  LAYER ME2 ;
  RECT 97.126 0.000 97.446 0.600 ;
  LAYER ME1 ;
  RECT 97.126 0.000 97.446 0.600 ;
 END
 ANTENNAPARTIALMETALAREA                  1.058 LAYER ME2 ;
 ANTENNAGATEAREA                          0.072 LAYER ME2 ;
 ANTENNAGATEAREA                          0.072 LAYER ME3 ;
 ANTENNAGATEAREA                          0.072 LAYER ME4 ;
 ANTENNADIFFAREA                          0.160 LAYER ME2 ;
 ANTENNADIFFAREA                          0.160 LAYER ME3 ;
 ANTENNADIFFAREA                          0.160 LAYER ME4 ;
 ANTENNAMAXAREACAR                       21.782 LAYER ME2 ;
 ANTENNAMAXAREACAR                       24.449 LAYER ME3 ;
 ANTENNAMAXAREACAR                       27.116 LAYER ME4 ;
END DI23
PIN DO23
  DIRECTION OUTPUT ;
 PORT
  LAYER ME4 ;
  RECT 96.564 0.000 96.884 0.600 ;
  LAYER ME3 ;
  RECT 96.564 0.000 96.884 0.600 ;
  LAYER ME2 ;
  RECT 96.564 0.000 96.884 0.600 ;
  LAYER ME1 ;
  RECT 96.564 0.000 96.884 0.600 ;
 END
 ANTENNAPARTIALMETALAREA                  5.273 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME3 ;
 ANTENNADIFFAREA                          1.293 LAYER ME4 ;
END DO23
PIN DI22
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 93.122 0.000 93.442 0.600 ;
  LAYER ME3 ;
  RECT 93.122 0.000 93.442 0.600 ;
  LAYER ME2 ;
  RECT 93.122 0.000 93.442 0.600 ;
  LAYER ME1 ;
  RECT 93.122 0.000 93.442 0.600 ;
 END
 ANTENNAPARTIALMETALAREA                  1.058 LAYER ME2 ;
 ANTENNAGATEAREA                          0.072 LAYER ME2 ;
 ANTENNAGATEAREA                          0.072 LAYER ME3 ;
 ANTENNAGATEAREA                          0.072 LAYER ME4 ;
 ANTENNADIFFAREA                          0.160 LAYER ME2 ;
 ANTENNADIFFAREA                          0.160 LAYER ME3 ;
 ANTENNADIFFAREA                          0.160 LAYER ME4 ;
 ANTENNAMAXAREACAR                       21.782 LAYER ME2 ;
 ANTENNAMAXAREACAR                       24.449 LAYER ME3 ;
 ANTENNAMAXAREACAR                       27.116 LAYER ME4 ;
END DI22
PIN DO22
  DIRECTION OUTPUT ;
 PORT
  LAYER ME4 ;
  RECT 92.560 0.000 92.880 0.600 ;
  LAYER ME3 ;
  RECT 92.560 0.000 92.880 0.600 ;
  LAYER ME2 ;
  RECT 92.560 0.000 92.880 0.600 ;
  LAYER ME1 ;
  RECT 92.560 0.000 92.880 0.600 ;
 END
 ANTENNAPARTIALMETALAREA                  5.273 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME3 ;
 ANTENNADIFFAREA                          1.293 LAYER ME4 ;
END DO22
PIN DI21
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 89.118 0.000 89.438 0.600 ;
  LAYER ME3 ;
  RECT 89.118 0.000 89.438 0.600 ;
  LAYER ME2 ;
  RECT 89.118 0.000 89.438 0.600 ;
  LAYER ME1 ;
  RECT 89.118 0.000 89.438 0.600 ;
 END
 ANTENNAPARTIALMETALAREA                  1.058 LAYER ME2 ;
 ANTENNAGATEAREA                          0.072 LAYER ME2 ;
 ANTENNAGATEAREA                          0.072 LAYER ME3 ;
 ANTENNAGATEAREA                          0.072 LAYER ME4 ;
 ANTENNADIFFAREA                          0.160 LAYER ME2 ;
 ANTENNADIFFAREA                          0.160 LAYER ME3 ;
 ANTENNADIFFAREA                          0.160 LAYER ME4 ;
 ANTENNAMAXAREACAR                       21.782 LAYER ME2 ;
 ANTENNAMAXAREACAR                       24.449 LAYER ME3 ;
 ANTENNAMAXAREACAR                       27.116 LAYER ME4 ;
END DI21
PIN DO21
  DIRECTION OUTPUT ;
 PORT
  LAYER ME4 ;
  RECT 88.556 0.000 88.876 0.600 ;
  LAYER ME3 ;
  RECT 88.556 0.000 88.876 0.600 ;
  LAYER ME2 ;
  RECT 88.556 0.000 88.876 0.600 ;
  LAYER ME1 ;
  RECT 88.556 0.000 88.876 0.600 ;
 END
 ANTENNAPARTIALMETALAREA                  5.273 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME3 ;
 ANTENNADIFFAREA                          1.293 LAYER ME4 ;
END DO21
PIN DI20
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 85.114 0.000 85.434 0.600 ;
  LAYER ME3 ;
  RECT 85.114 0.000 85.434 0.600 ;
  LAYER ME2 ;
  RECT 85.114 0.000 85.434 0.600 ;
  LAYER ME1 ;
  RECT 85.114 0.000 85.434 0.600 ;
 END
 ANTENNAPARTIALMETALAREA                  1.058 LAYER ME2 ;
 ANTENNAGATEAREA                          0.072 LAYER ME2 ;
 ANTENNAGATEAREA                          0.072 LAYER ME3 ;
 ANTENNAGATEAREA                          0.072 LAYER ME4 ;
 ANTENNADIFFAREA                          0.160 LAYER ME2 ;
 ANTENNADIFFAREA                          0.160 LAYER ME3 ;
 ANTENNADIFFAREA                          0.160 LAYER ME4 ;
 ANTENNAMAXAREACAR                       21.782 LAYER ME2 ;
 ANTENNAMAXAREACAR                       24.449 LAYER ME3 ;
 ANTENNAMAXAREACAR                       27.116 LAYER ME4 ;
END DI20
PIN DO20
  DIRECTION OUTPUT ;
 PORT
  LAYER ME4 ;
  RECT 84.552 0.000 84.872 0.600 ;
  LAYER ME3 ;
  RECT 84.552 0.000 84.872 0.600 ;
  LAYER ME2 ;
  RECT 84.552 0.000 84.872 0.600 ;
  LAYER ME1 ;
  RECT 84.552 0.000 84.872 0.600 ;
 END
 ANTENNAPARTIALMETALAREA                  5.273 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME3 ;
 ANTENNADIFFAREA                          1.293 LAYER ME4 ;
END DO20
PIN DI19
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 81.110 0.000 81.430 0.600 ;
  LAYER ME3 ;
  RECT 81.110 0.000 81.430 0.600 ;
  LAYER ME2 ;
  RECT 81.110 0.000 81.430 0.600 ;
  LAYER ME1 ;
  RECT 81.110 0.000 81.430 0.600 ;
 END
 ANTENNAPARTIALMETALAREA                  1.058 LAYER ME2 ;
 ANTENNAGATEAREA                          0.072 LAYER ME2 ;
 ANTENNAGATEAREA                          0.072 LAYER ME3 ;
 ANTENNAGATEAREA                          0.072 LAYER ME4 ;
 ANTENNADIFFAREA                          0.160 LAYER ME2 ;
 ANTENNADIFFAREA                          0.160 LAYER ME3 ;
 ANTENNADIFFAREA                          0.160 LAYER ME4 ;
 ANTENNAMAXAREACAR                       21.782 LAYER ME2 ;
 ANTENNAMAXAREACAR                       24.449 LAYER ME3 ;
 ANTENNAMAXAREACAR                       27.116 LAYER ME4 ;
END DI19
PIN DO19
  DIRECTION OUTPUT ;
 PORT
  LAYER ME4 ;
  RECT 80.548 0.000 80.868 0.600 ;
  LAYER ME3 ;
  RECT 80.548 0.000 80.868 0.600 ;
  LAYER ME2 ;
  RECT 80.548 0.000 80.868 0.600 ;
  LAYER ME1 ;
  RECT 80.548 0.000 80.868 0.600 ;
 END
 ANTENNAPARTIALMETALAREA                  5.273 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME3 ;
 ANTENNADIFFAREA                          1.293 LAYER ME4 ;
END DO19
PIN DI18
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 77.106 0.000 77.426 0.600 ;
  LAYER ME3 ;
  RECT 77.106 0.000 77.426 0.600 ;
  LAYER ME2 ;
  RECT 77.106 0.000 77.426 0.600 ;
  LAYER ME1 ;
  RECT 77.106 0.000 77.426 0.600 ;
 END
 ANTENNAPARTIALMETALAREA                  1.058 LAYER ME2 ;
 ANTENNAGATEAREA                          0.072 LAYER ME2 ;
 ANTENNAGATEAREA                          0.072 LAYER ME3 ;
 ANTENNAGATEAREA                          0.072 LAYER ME4 ;
 ANTENNADIFFAREA                          0.160 LAYER ME2 ;
 ANTENNADIFFAREA                          0.160 LAYER ME3 ;
 ANTENNADIFFAREA                          0.160 LAYER ME4 ;
 ANTENNAMAXAREACAR                       21.782 LAYER ME2 ;
 ANTENNAMAXAREACAR                       24.449 LAYER ME3 ;
 ANTENNAMAXAREACAR                       27.116 LAYER ME4 ;
END DI18
PIN DO18
  DIRECTION OUTPUT ;
 PORT
  LAYER ME4 ;
  RECT 76.544 0.000 76.864 0.600 ;
  LAYER ME3 ;
  RECT 76.544 0.000 76.864 0.600 ;
  LAYER ME2 ;
  RECT 76.544 0.000 76.864 0.600 ;
  LAYER ME1 ;
  RECT 76.544 0.000 76.864 0.600 ;
 END
 ANTENNAPARTIALMETALAREA                  5.273 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME3 ;
 ANTENNADIFFAREA                          1.293 LAYER ME4 ;
END DO18
PIN DI17
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 73.102 0.000 73.422 0.600 ;
  LAYER ME3 ;
  RECT 73.102 0.000 73.422 0.600 ;
  LAYER ME2 ;
  RECT 73.102 0.000 73.422 0.600 ;
  LAYER ME1 ;
  RECT 73.102 0.000 73.422 0.600 ;
 END
 ANTENNAPARTIALMETALAREA                  1.058 LAYER ME2 ;
 ANTENNAGATEAREA                          0.072 LAYER ME2 ;
 ANTENNAGATEAREA                          0.072 LAYER ME3 ;
 ANTENNAGATEAREA                          0.072 LAYER ME4 ;
 ANTENNADIFFAREA                          0.160 LAYER ME2 ;
 ANTENNADIFFAREA                          0.160 LAYER ME3 ;
 ANTENNADIFFAREA                          0.160 LAYER ME4 ;
 ANTENNAMAXAREACAR                       21.782 LAYER ME2 ;
 ANTENNAMAXAREACAR                       24.449 LAYER ME3 ;
 ANTENNAMAXAREACAR                       27.116 LAYER ME4 ;
END DI17
PIN DO17
  DIRECTION OUTPUT ;
 PORT
  LAYER ME4 ;
  RECT 72.540 0.000 72.860 0.600 ;
  LAYER ME3 ;
  RECT 72.540 0.000 72.860 0.600 ;
  LAYER ME2 ;
  RECT 72.540 0.000 72.860 0.600 ;
  LAYER ME1 ;
  RECT 72.540 0.000 72.860 0.600 ;
 END
 ANTENNAPARTIALMETALAREA                  5.273 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME3 ;
 ANTENNADIFFAREA                          1.293 LAYER ME4 ;
END DO17
PIN DI16
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 68.536 0.000 68.856 0.600 ;
  LAYER ME3 ;
  RECT 68.536 0.000 68.856 0.600 ;
  LAYER ME2 ;
  RECT 68.536 0.000 68.856 0.600 ;
  LAYER ME1 ;
  RECT 68.536 0.000 68.856 0.600 ;
 END
 ANTENNAPARTIALMETALAREA                  0.346 LAYER ME1 ;
 ANTENNAPARTIALMETALAREA                  1.466 LAYER ME2 ;
 ANTENNAPARTIALMETALAREA                  0.508 LAYER ME3 ;
 ANTENNAGATEAREA                          0.072 LAYER ME3 ;
 ANTENNAGATEAREA                          0.072 LAYER ME4 ;
 ANTENNADIFFAREA                          0.218 LAYER ME1 ;
 ANTENNADIFFAREA                          0.218 LAYER ME2 ;
 ANTENNADIFFAREA                          0.218 LAYER ME3 ;
 ANTENNADIFFAREA                          0.218 LAYER ME4 ;
 ANTENNAMAXAREACAR                       17.267 LAYER ME3 ;
 ANTENNAMAXAREACAR                       19.933 LAYER ME4 ;
END DI16
PIN DO16
  DIRECTION OUTPUT ;
 PORT
  LAYER ME4 ;
  RECT 69.098 0.000 69.418 0.600 ;
  LAYER ME3 ;
  RECT 69.098 0.000 69.418 0.600 ;
  LAYER ME2 ;
  RECT 69.098 0.000 69.418 0.600 ;
  LAYER ME1 ;
  RECT 69.098 0.000 69.418 0.600 ;
 END
 ANTENNAPARTIALMETALAREA                  5.602 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME3 ;
 ANTENNADIFFAREA                          1.293 LAYER ME4 ;
END DO16
PIN WEB1
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 67.096 0.000 67.416 0.600 ;
  LAYER ME3 ;
  RECT 67.096 0.000 67.416 0.600 ;
  LAYER ME2 ;
  RECT 67.096 0.000 67.416 0.600 ;
  LAYER ME1 ;
  RECT 67.096 0.000 67.416 0.600 ;
 END
 ANTENNAPARTIALMETALAREA                  1.036 LAYER ME2 ;
 ANTENNAGATEAREA                          0.288 LAYER ME2 ;
 ANTENNAGATEAREA                          0.288 LAYER ME3 ;
 ANTENNAGATEAREA                          0.288 LAYER ME4 ;
 ANTENNADIFFAREA                          0.206 LAYER ME2 ;
 ANTENNADIFFAREA                          0.206 LAYER ME3 ;
 ANTENNADIFFAREA                          0.206 LAYER ME4 ;
 ANTENNAMAXAREACAR                        5.844 LAYER ME2 ;
 ANTENNAMAXAREACAR                        6.511 LAYER ME3 ;
 ANTENNAMAXAREACAR                        7.178 LAYER ME4 ;
END WEB1
PIN DI15
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 65.094 0.000 65.414 0.600 ;
  LAYER ME3 ;
  RECT 65.094 0.000 65.414 0.600 ;
  LAYER ME2 ;
  RECT 65.094 0.000 65.414 0.600 ;
  LAYER ME1 ;
  RECT 65.094 0.000 65.414 0.600 ;
 END
 ANTENNAPARTIALMETALAREA                  1.058 LAYER ME2 ;
 ANTENNAGATEAREA                          0.072 LAYER ME2 ;
 ANTENNAGATEAREA                          0.072 LAYER ME3 ;
 ANTENNAGATEAREA                          0.072 LAYER ME4 ;
 ANTENNADIFFAREA                          0.160 LAYER ME2 ;
 ANTENNADIFFAREA                          0.160 LAYER ME3 ;
 ANTENNADIFFAREA                          0.160 LAYER ME4 ;
 ANTENNAMAXAREACAR                       21.782 LAYER ME2 ;
 ANTENNAMAXAREACAR                       24.449 LAYER ME3 ;
 ANTENNAMAXAREACAR                       27.116 LAYER ME4 ;
END DI15
PIN DO15
  DIRECTION OUTPUT ;
 PORT
  LAYER ME4 ;
  RECT 64.532 0.000 64.852 0.600 ;
  LAYER ME3 ;
  RECT 64.532 0.000 64.852 0.600 ;
  LAYER ME2 ;
  RECT 64.532 0.000 64.852 0.600 ;
  LAYER ME1 ;
  RECT 64.532 0.000 64.852 0.600 ;
 END
 ANTENNAPARTIALMETALAREA                  5.273 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME3 ;
 ANTENNADIFFAREA                          1.293 LAYER ME4 ;
END DO15
PIN DI14
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 61.090 0.000 61.410 0.600 ;
  LAYER ME3 ;
  RECT 61.090 0.000 61.410 0.600 ;
  LAYER ME2 ;
  RECT 61.090 0.000 61.410 0.600 ;
  LAYER ME1 ;
  RECT 61.090 0.000 61.410 0.600 ;
 END
 ANTENNAPARTIALMETALAREA                  1.058 LAYER ME2 ;
 ANTENNAGATEAREA                          0.072 LAYER ME2 ;
 ANTENNAGATEAREA                          0.072 LAYER ME3 ;
 ANTENNAGATEAREA                          0.072 LAYER ME4 ;
 ANTENNADIFFAREA                          0.160 LAYER ME2 ;
 ANTENNADIFFAREA                          0.160 LAYER ME3 ;
 ANTENNADIFFAREA                          0.160 LAYER ME4 ;
 ANTENNAMAXAREACAR                       21.782 LAYER ME2 ;
 ANTENNAMAXAREACAR                       24.449 LAYER ME3 ;
 ANTENNAMAXAREACAR                       27.116 LAYER ME4 ;
END DI14
PIN DO14
  DIRECTION OUTPUT ;
 PORT
  LAYER ME4 ;
  RECT 60.528 0.000 60.848 0.600 ;
  LAYER ME3 ;
  RECT 60.528 0.000 60.848 0.600 ;
  LAYER ME2 ;
  RECT 60.528 0.000 60.848 0.600 ;
  LAYER ME1 ;
  RECT 60.528 0.000 60.848 0.600 ;
 END
 ANTENNAPARTIALMETALAREA                  5.273 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME3 ;
 ANTENNADIFFAREA                          1.293 LAYER ME4 ;
END DO14
PIN DI13
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 57.086 0.000 57.406 0.600 ;
  LAYER ME3 ;
  RECT 57.086 0.000 57.406 0.600 ;
  LAYER ME2 ;
  RECT 57.086 0.000 57.406 0.600 ;
  LAYER ME1 ;
  RECT 57.086 0.000 57.406 0.600 ;
 END
 ANTENNAPARTIALMETALAREA                  1.058 LAYER ME2 ;
 ANTENNAGATEAREA                          0.072 LAYER ME2 ;
 ANTENNAGATEAREA                          0.072 LAYER ME3 ;
 ANTENNAGATEAREA                          0.072 LAYER ME4 ;
 ANTENNADIFFAREA                          0.160 LAYER ME2 ;
 ANTENNADIFFAREA                          0.160 LAYER ME3 ;
 ANTENNADIFFAREA                          0.160 LAYER ME4 ;
 ANTENNAMAXAREACAR                       21.782 LAYER ME2 ;
 ANTENNAMAXAREACAR                       24.449 LAYER ME3 ;
 ANTENNAMAXAREACAR                       27.116 LAYER ME4 ;
END DI13
PIN DO13
  DIRECTION OUTPUT ;
 PORT
  LAYER ME4 ;
  RECT 56.524 0.000 56.844 0.600 ;
  LAYER ME3 ;
  RECT 56.524 0.000 56.844 0.600 ;
  LAYER ME2 ;
  RECT 56.524 0.000 56.844 0.600 ;
  LAYER ME1 ;
  RECT 56.524 0.000 56.844 0.600 ;
 END
 ANTENNAPARTIALMETALAREA                  5.273 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME3 ;
 ANTENNADIFFAREA                          1.293 LAYER ME4 ;
END DO13
PIN DI12
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 53.082 0.000 53.402 0.600 ;
  LAYER ME3 ;
  RECT 53.082 0.000 53.402 0.600 ;
  LAYER ME2 ;
  RECT 53.082 0.000 53.402 0.600 ;
  LAYER ME1 ;
  RECT 53.082 0.000 53.402 0.600 ;
 END
 ANTENNAPARTIALMETALAREA                  1.058 LAYER ME2 ;
 ANTENNAGATEAREA                          0.072 LAYER ME2 ;
 ANTENNAGATEAREA                          0.072 LAYER ME3 ;
 ANTENNAGATEAREA                          0.072 LAYER ME4 ;
 ANTENNADIFFAREA                          0.160 LAYER ME2 ;
 ANTENNADIFFAREA                          0.160 LAYER ME3 ;
 ANTENNADIFFAREA                          0.160 LAYER ME4 ;
 ANTENNAMAXAREACAR                       21.782 LAYER ME2 ;
 ANTENNAMAXAREACAR                       24.449 LAYER ME3 ;
 ANTENNAMAXAREACAR                       27.116 LAYER ME4 ;
END DI12
PIN DO12
  DIRECTION OUTPUT ;
 PORT
  LAYER ME4 ;
  RECT 52.520 0.000 52.840 0.600 ;
  LAYER ME3 ;
  RECT 52.520 0.000 52.840 0.600 ;
  LAYER ME2 ;
  RECT 52.520 0.000 52.840 0.600 ;
  LAYER ME1 ;
  RECT 52.520 0.000 52.840 0.600 ;
 END
 ANTENNAPARTIALMETALAREA                  5.273 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME3 ;
 ANTENNADIFFAREA                          1.293 LAYER ME4 ;
END DO12
PIN DI11
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 49.078 0.000 49.398 0.600 ;
  LAYER ME3 ;
  RECT 49.078 0.000 49.398 0.600 ;
  LAYER ME2 ;
  RECT 49.078 0.000 49.398 0.600 ;
  LAYER ME1 ;
  RECT 49.078 0.000 49.398 0.600 ;
 END
 ANTENNAPARTIALMETALAREA                  1.058 LAYER ME2 ;
 ANTENNAGATEAREA                          0.072 LAYER ME2 ;
 ANTENNAGATEAREA                          0.072 LAYER ME3 ;
 ANTENNAGATEAREA                          0.072 LAYER ME4 ;
 ANTENNADIFFAREA                          0.160 LAYER ME2 ;
 ANTENNADIFFAREA                          0.160 LAYER ME3 ;
 ANTENNADIFFAREA                          0.160 LAYER ME4 ;
 ANTENNAMAXAREACAR                       21.782 LAYER ME2 ;
 ANTENNAMAXAREACAR                       24.449 LAYER ME3 ;
 ANTENNAMAXAREACAR                       27.116 LAYER ME4 ;
END DI11
PIN DO11
  DIRECTION OUTPUT ;
 PORT
  LAYER ME4 ;
  RECT 48.516 0.000 48.836 0.600 ;
  LAYER ME3 ;
  RECT 48.516 0.000 48.836 0.600 ;
  LAYER ME2 ;
  RECT 48.516 0.000 48.836 0.600 ;
  LAYER ME1 ;
  RECT 48.516 0.000 48.836 0.600 ;
 END
 ANTENNAPARTIALMETALAREA                  5.273 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME3 ;
 ANTENNADIFFAREA                          1.293 LAYER ME4 ;
END DO11
PIN DI10
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 45.074 0.000 45.394 0.600 ;
  LAYER ME3 ;
  RECT 45.074 0.000 45.394 0.600 ;
  LAYER ME2 ;
  RECT 45.074 0.000 45.394 0.600 ;
  LAYER ME1 ;
  RECT 45.074 0.000 45.394 0.600 ;
 END
 ANTENNAPARTIALMETALAREA                  1.058 LAYER ME2 ;
 ANTENNAGATEAREA                          0.072 LAYER ME2 ;
 ANTENNAGATEAREA                          0.072 LAYER ME3 ;
 ANTENNAGATEAREA                          0.072 LAYER ME4 ;
 ANTENNADIFFAREA                          0.160 LAYER ME2 ;
 ANTENNADIFFAREA                          0.160 LAYER ME3 ;
 ANTENNADIFFAREA                          0.160 LAYER ME4 ;
 ANTENNAMAXAREACAR                       21.782 LAYER ME2 ;
 ANTENNAMAXAREACAR                       24.449 LAYER ME3 ;
 ANTENNAMAXAREACAR                       27.116 LAYER ME4 ;
END DI10
PIN DO10
  DIRECTION OUTPUT ;
 PORT
  LAYER ME4 ;
  RECT 44.512 0.000 44.832 0.600 ;
  LAYER ME3 ;
  RECT 44.512 0.000 44.832 0.600 ;
  LAYER ME2 ;
  RECT 44.512 0.000 44.832 0.600 ;
  LAYER ME1 ;
  RECT 44.512 0.000 44.832 0.600 ;
 END
 ANTENNAPARTIALMETALAREA                  5.273 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME3 ;
 ANTENNADIFFAREA                          1.293 LAYER ME4 ;
END DO10
PIN DI9
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 41.070 0.000 41.390 0.600 ;
  LAYER ME3 ;
  RECT 41.070 0.000 41.390 0.600 ;
  LAYER ME2 ;
  RECT 41.070 0.000 41.390 0.600 ;
  LAYER ME1 ;
  RECT 41.070 0.000 41.390 0.600 ;
 END
 ANTENNAPARTIALMETALAREA                  1.058 LAYER ME2 ;
 ANTENNAGATEAREA                          0.072 LAYER ME2 ;
 ANTENNAGATEAREA                          0.072 LAYER ME3 ;
 ANTENNAGATEAREA                          0.072 LAYER ME4 ;
 ANTENNADIFFAREA                          0.160 LAYER ME2 ;
 ANTENNADIFFAREA                          0.160 LAYER ME3 ;
 ANTENNADIFFAREA                          0.160 LAYER ME4 ;
 ANTENNAMAXAREACAR                       21.782 LAYER ME2 ;
 ANTENNAMAXAREACAR                       24.449 LAYER ME3 ;
 ANTENNAMAXAREACAR                       27.116 LAYER ME4 ;
END DI9
PIN DO9
  DIRECTION OUTPUT ;
 PORT
  LAYER ME4 ;
  RECT 40.508 0.000 40.828 0.600 ;
  LAYER ME3 ;
  RECT 40.508 0.000 40.828 0.600 ;
  LAYER ME2 ;
  RECT 40.508 0.000 40.828 0.600 ;
  LAYER ME1 ;
  RECT 40.508 0.000 40.828 0.600 ;
 END
 ANTENNAPARTIALMETALAREA                  5.273 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME3 ;
 ANTENNADIFFAREA                          1.293 LAYER ME4 ;
END DO9
PIN DI8
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 37.066 0.000 37.386 0.600 ;
  LAYER ME3 ;
  RECT 37.066 0.000 37.386 0.600 ;
  LAYER ME2 ;
  RECT 37.066 0.000 37.386 0.600 ;
  LAYER ME1 ;
  RECT 37.066 0.000 37.386 0.600 ;
 END
 ANTENNAPARTIALMETALAREA                  1.058 LAYER ME2 ;
 ANTENNAGATEAREA                          0.072 LAYER ME2 ;
 ANTENNAGATEAREA                          0.072 LAYER ME3 ;
 ANTENNAGATEAREA                          0.072 LAYER ME4 ;
 ANTENNADIFFAREA                          0.160 LAYER ME2 ;
 ANTENNADIFFAREA                          0.160 LAYER ME3 ;
 ANTENNADIFFAREA                          0.160 LAYER ME4 ;
 ANTENNAMAXAREACAR                       21.782 LAYER ME2 ;
 ANTENNAMAXAREACAR                       24.449 LAYER ME3 ;
 ANTENNAMAXAREACAR                       27.116 LAYER ME4 ;
END DI8
PIN DO8
  DIRECTION OUTPUT ;
 PORT
  LAYER ME4 ;
  RECT 36.504 0.000 36.824 0.600 ;
  LAYER ME3 ;
  RECT 36.504 0.000 36.824 0.600 ;
  LAYER ME2 ;
  RECT 36.504 0.000 36.824 0.600 ;
  LAYER ME1 ;
  RECT 36.504 0.000 36.824 0.600 ;
 END
 ANTENNAPARTIALMETALAREA                  5.273 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME3 ;
 ANTENNADIFFAREA                          1.293 LAYER ME4 ;
END DO8
PIN DI7
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 33.062 0.000 33.382 0.600 ;
  LAYER ME3 ;
  RECT 33.062 0.000 33.382 0.600 ;
  LAYER ME2 ;
  RECT 33.062 0.000 33.382 0.600 ;
  LAYER ME1 ;
  RECT 33.062 0.000 33.382 0.600 ;
 END
 ANTENNAPARTIALMETALAREA                  1.058 LAYER ME2 ;
 ANTENNAGATEAREA                          0.072 LAYER ME2 ;
 ANTENNAGATEAREA                          0.072 LAYER ME3 ;
 ANTENNAGATEAREA                          0.072 LAYER ME4 ;
 ANTENNADIFFAREA                          0.160 LAYER ME2 ;
 ANTENNADIFFAREA                          0.160 LAYER ME3 ;
 ANTENNADIFFAREA                          0.160 LAYER ME4 ;
 ANTENNAMAXAREACAR                       21.782 LAYER ME2 ;
 ANTENNAMAXAREACAR                       24.449 LAYER ME3 ;
 ANTENNAMAXAREACAR                       27.116 LAYER ME4 ;
END DI7
PIN DO7
  DIRECTION OUTPUT ;
 PORT
  LAYER ME4 ;
  RECT 32.500 0.000 32.820 0.600 ;
  LAYER ME3 ;
  RECT 32.500 0.000 32.820 0.600 ;
  LAYER ME2 ;
  RECT 32.500 0.000 32.820 0.600 ;
  LAYER ME1 ;
  RECT 32.500 0.000 32.820 0.600 ;
 END
 ANTENNAPARTIALMETALAREA                  5.273 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME3 ;
 ANTENNADIFFAREA                          1.293 LAYER ME4 ;
END DO7
PIN DI6
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 29.058 0.000 29.378 0.600 ;
  LAYER ME3 ;
  RECT 29.058 0.000 29.378 0.600 ;
  LAYER ME2 ;
  RECT 29.058 0.000 29.378 0.600 ;
  LAYER ME1 ;
  RECT 29.058 0.000 29.378 0.600 ;
 END
 ANTENNAPARTIALMETALAREA                  1.058 LAYER ME2 ;
 ANTENNAGATEAREA                          0.072 LAYER ME2 ;
 ANTENNAGATEAREA                          0.072 LAYER ME3 ;
 ANTENNAGATEAREA                          0.072 LAYER ME4 ;
 ANTENNADIFFAREA                          0.160 LAYER ME2 ;
 ANTENNADIFFAREA                          0.160 LAYER ME3 ;
 ANTENNADIFFAREA                          0.160 LAYER ME4 ;
 ANTENNAMAXAREACAR                       21.782 LAYER ME2 ;
 ANTENNAMAXAREACAR                       24.449 LAYER ME3 ;
 ANTENNAMAXAREACAR                       27.116 LAYER ME4 ;
END DI6
PIN DO6
  DIRECTION OUTPUT ;
 PORT
  LAYER ME4 ;
  RECT 28.496 0.000 28.816 0.600 ;
  LAYER ME3 ;
  RECT 28.496 0.000 28.816 0.600 ;
  LAYER ME2 ;
  RECT 28.496 0.000 28.816 0.600 ;
  LAYER ME1 ;
  RECT 28.496 0.000 28.816 0.600 ;
 END
 ANTENNAPARTIALMETALAREA                  5.273 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME3 ;
 ANTENNADIFFAREA                          1.293 LAYER ME4 ;
END DO6
PIN DI5
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 25.054 0.000 25.374 0.600 ;
  LAYER ME3 ;
  RECT 25.054 0.000 25.374 0.600 ;
  LAYER ME2 ;
  RECT 25.054 0.000 25.374 0.600 ;
  LAYER ME1 ;
  RECT 25.054 0.000 25.374 0.600 ;
 END
 ANTENNAPARTIALMETALAREA                  1.058 LAYER ME2 ;
 ANTENNAGATEAREA                          0.072 LAYER ME2 ;
 ANTENNAGATEAREA                          0.072 LAYER ME3 ;
 ANTENNAGATEAREA                          0.072 LAYER ME4 ;
 ANTENNADIFFAREA                          0.160 LAYER ME2 ;
 ANTENNADIFFAREA                          0.160 LAYER ME3 ;
 ANTENNADIFFAREA                          0.160 LAYER ME4 ;
 ANTENNAMAXAREACAR                       21.782 LAYER ME2 ;
 ANTENNAMAXAREACAR                       24.449 LAYER ME3 ;
 ANTENNAMAXAREACAR                       27.116 LAYER ME4 ;
END DI5
PIN DO5
  DIRECTION OUTPUT ;
 PORT
  LAYER ME4 ;
  RECT 24.492 0.000 24.812 0.600 ;
  LAYER ME3 ;
  RECT 24.492 0.000 24.812 0.600 ;
  LAYER ME2 ;
  RECT 24.492 0.000 24.812 0.600 ;
  LAYER ME1 ;
  RECT 24.492 0.000 24.812 0.600 ;
 END
 ANTENNAPARTIALMETALAREA                  5.273 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME3 ;
 ANTENNADIFFAREA                          1.293 LAYER ME4 ;
END DO5
PIN DI4
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 21.050 0.000 21.370 0.600 ;
  LAYER ME3 ;
  RECT 21.050 0.000 21.370 0.600 ;
  LAYER ME2 ;
  RECT 21.050 0.000 21.370 0.600 ;
  LAYER ME1 ;
  RECT 21.050 0.000 21.370 0.600 ;
 END
 ANTENNAPARTIALMETALAREA                  1.058 LAYER ME2 ;
 ANTENNAGATEAREA                          0.072 LAYER ME2 ;
 ANTENNAGATEAREA                          0.072 LAYER ME3 ;
 ANTENNAGATEAREA                          0.072 LAYER ME4 ;
 ANTENNADIFFAREA                          0.160 LAYER ME2 ;
 ANTENNADIFFAREA                          0.160 LAYER ME3 ;
 ANTENNADIFFAREA                          0.160 LAYER ME4 ;
 ANTENNAMAXAREACAR                       21.782 LAYER ME2 ;
 ANTENNAMAXAREACAR                       24.449 LAYER ME3 ;
 ANTENNAMAXAREACAR                       27.116 LAYER ME4 ;
END DI4
PIN DO4
  DIRECTION OUTPUT ;
 PORT
  LAYER ME4 ;
  RECT 20.488 0.000 20.808 0.600 ;
  LAYER ME3 ;
  RECT 20.488 0.000 20.808 0.600 ;
  LAYER ME2 ;
  RECT 20.488 0.000 20.808 0.600 ;
  LAYER ME1 ;
  RECT 20.488 0.000 20.808 0.600 ;
 END
 ANTENNAPARTIALMETALAREA                  5.273 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME3 ;
 ANTENNADIFFAREA                          1.293 LAYER ME4 ;
END DO4
PIN DI3
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 17.046 0.000 17.366 0.600 ;
  LAYER ME3 ;
  RECT 17.046 0.000 17.366 0.600 ;
  LAYER ME2 ;
  RECT 17.046 0.000 17.366 0.600 ;
  LAYER ME1 ;
  RECT 17.046 0.000 17.366 0.600 ;
 END
 ANTENNAPARTIALMETALAREA                  1.058 LAYER ME2 ;
 ANTENNAGATEAREA                          0.072 LAYER ME2 ;
 ANTENNAGATEAREA                          0.072 LAYER ME3 ;
 ANTENNAGATEAREA                          0.072 LAYER ME4 ;
 ANTENNADIFFAREA                          0.160 LAYER ME2 ;
 ANTENNADIFFAREA                          0.160 LAYER ME3 ;
 ANTENNADIFFAREA                          0.160 LAYER ME4 ;
 ANTENNAMAXAREACAR                       21.782 LAYER ME2 ;
 ANTENNAMAXAREACAR                       24.449 LAYER ME3 ;
 ANTENNAMAXAREACAR                       27.116 LAYER ME4 ;
END DI3
PIN DO3
  DIRECTION OUTPUT ;
 PORT
  LAYER ME4 ;
  RECT 16.484 0.000 16.804 0.600 ;
  LAYER ME3 ;
  RECT 16.484 0.000 16.804 0.600 ;
  LAYER ME2 ;
  RECT 16.484 0.000 16.804 0.600 ;
  LAYER ME1 ;
  RECT 16.484 0.000 16.804 0.600 ;
 END
 ANTENNAPARTIALMETALAREA                  5.273 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME3 ;
 ANTENNADIFFAREA                          1.293 LAYER ME4 ;
END DO3
PIN DI2
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 13.042 0.000 13.362 0.600 ;
  LAYER ME3 ;
  RECT 13.042 0.000 13.362 0.600 ;
  LAYER ME2 ;
  RECT 13.042 0.000 13.362 0.600 ;
  LAYER ME1 ;
  RECT 13.042 0.000 13.362 0.600 ;
 END
 ANTENNAPARTIALMETALAREA                  1.058 LAYER ME2 ;
 ANTENNAGATEAREA                          0.072 LAYER ME2 ;
 ANTENNAGATEAREA                          0.072 LAYER ME3 ;
 ANTENNAGATEAREA                          0.072 LAYER ME4 ;
 ANTENNADIFFAREA                          0.160 LAYER ME2 ;
 ANTENNADIFFAREA                          0.160 LAYER ME3 ;
 ANTENNADIFFAREA                          0.160 LAYER ME4 ;
 ANTENNAMAXAREACAR                       21.782 LAYER ME2 ;
 ANTENNAMAXAREACAR                       24.449 LAYER ME3 ;
 ANTENNAMAXAREACAR                       27.116 LAYER ME4 ;
END DI2
PIN DO2
  DIRECTION OUTPUT ;
 PORT
  LAYER ME4 ;
  RECT 12.480 0.000 12.800 0.600 ;
  LAYER ME3 ;
  RECT 12.480 0.000 12.800 0.600 ;
  LAYER ME2 ;
  RECT 12.480 0.000 12.800 0.600 ;
  LAYER ME1 ;
  RECT 12.480 0.000 12.800 0.600 ;
 END
 ANTENNAPARTIALMETALAREA                  5.273 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME3 ;
 ANTENNADIFFAREA                          1.293 LAYER ME4 ;
END DO2
PIN DI1
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 9.038 0.000 9.358 0.600 ;
  LAYER ME3 ;
  RECT 9.038 0.000 9.358 0.600 ;
  LAYER ME2 ;
  RECT 9.038 0.000 9.358 0.600 ;
  LAYER ME1 ;
  RECT 9.038 0.000 9.358 0.600 ;
 END
 ANTENNAPARTIALMETALAREA                  1.058 LAYER ME2 ;
 ANTENNAGATEAREA                          0.072 LAYER ME2 ;
 ANTENNAGATEAREA                          0.072 LAYER ME3 ;
 ANTENNAGATEAREA                          0.072 LAYER ME4 ;
 ANTENNADIFFAREA                          0.160 LAYER ME2 ;
 ANTENNADIFFAREA                          0.160 LAYER ME3 ;
 ANTENNADIFFAREA                          0.160 LAYER ME4 ;
 ANTENNAMAXAREACAR                       21.782 LAYER ME2 ;
 ANTENNAMAXAREACAR                       24.449 LAYER ME3 ;
 ANTENNAMAXAREACAR                       27.116 LAYER ME4 ;
END DI1
PIN DO1
  DIRECTION OUTPUT ;
 PORT
  LAYER ME4 ;
  RECT 8.476 0.000 8.796 0.600 ;
  LAYER ME3 ;
  RECT 8.476 0.000 8.796 0.600 ;
  LAYER ME2 ;
  RECT 8.476 0.000 8.796 0.600 ;
  LAYER ME1 ;
  RECT 8.476 0.000 8.796 0.600 ;
 END
 ANTENNAPARTIALMETALAREA                  5.273 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME3 ;
 ANTENNADIFFAREA                          1.293 LAYER ME4 ;
END DO1
PIN DI0
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 4.472 0.000 4.792 0.600 ;
  LAYER ME3 ;
  RECT 4.472 0.000 4.792 0.600 ;
  LAYER ME2 ;
  RECT 4.472 0.000 4.792 0.600 ;
  LAYER ME1 ;
  RECT 4.472 0.000 4.792 0.600 ;
 END
 ANTENNAPARTIALMETALAREA                  0.346 LAYER ME1 ;
 ANTENNAPARTIALMETALAREA                  1.466 LAYER ME2 ;
 ANTENNAPARTIALMETALAREA                  0.508 LAYER ME3 ;
 ANTENNAGATEAREA                          0.072 LAYER ME3 ;
 ANTENNAGATEAREA                          0.072 LAYER ME4 ;
 ANTENNADIFFAREA                          0.218 LAYER ME1 ;
 ANTENNADIFFAREA                          0.218 LAYER ME2 ;
 ANTENNADIFFAREA                          0.218 LAYER ME3 ;
 ANTENNADIFFAREA                          0.218 LAYER ME4 ;
 ANTENNAMAXAREACAR                       17.267 LAYER ME3 ;
 ANTENNAMAXAREACAR                       19.933 LAYER ME4 ;
END DI0
PIN DO0
  DIRECTION OUTPUT ;
 PORT
  LAYER ME4 ;
  RECT 5.034 0.000 5.354 0.600 ;
  LAYER ME3 ;
  RECT 5.034 0.000 5.354 0.600 ;
  LAYER ME2 ;
  RECT 5.034 0.000 5.354 0.600 ;
  LAYER ME1 ;
  RECT 5.034 0.000 5.354 0.600 ;
 END
 ANTENNAPARTIALMETALAREA                  5.602 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME3 ;
 ANTENNADIFFAREA                          1.293 LAYER ME4 ;
END DO0
PIN WEB0
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 3.032 0.000 3.352 0.600 ;
  LAYER ME3 ;
  RECT 3.032 0.000 3.352 0.600 ;
  LAYER ME2 ;
  RECT 3.032 0.000 3.352 0.600 ;
  LAYER ME1 ;
  RECT 3.032 0.000 3.352 0.600 ;
 END
 ANTENNAPARTIALMETALAREA                  1.036 LAYER ME2 ;
 ANTENNAGATEAREA                          0.288 LAYER ME2 ;
 ANTENNAGATEAREA                          0.288 LAYER ME3 ;
 ANTENNAGATEAREA                          0.288 LAYER ME4 ;
 ANTENNADIFFAREA                          0.206 LAYER ME2 ;
 ANTENNADIFFAREA                          0.206 LAYER ME3 ;
 ANTENNADIFFAREA                          0.206 LAYER ME4 ;
 ANTENNAMAXAREACAR                        5.844 LAYER ME2 ;
 ANTENNAMAXAREACAR                        6.511 LAYER ME3 ;
 ANTENNAMAXAREACAR                        7.178 LAYER ME4 ;
END WEB0
PIN A1
  DIRECTION INPUT ;
 PORT
  LAYER ME3 ;
  RECT 276.736 0.000 277.056 0.720 ;
  LAYER ME2 ;
  RECT 276.736 0.000 277.056 0.720 ;
  LAYER ME1 ;
  RECT 276.736 0.000 277.056 0.720 ;
 END
 ANTENNAPARTIALMETALAREA                  3.547 LAYER ME2 ;
 ANTENNAGATEAREA                          0.144 LAYER ME2 ;
 ANTENNAGATEAREA                          0.144 LAYER ME3 ;
 ANTENNADIFFAREA                          0.218 LAYER ME2 ;
 ANTENNADIFFAREA                          0.218 LAYER ME3 ;
 ANTENNAMAXAREACAR                       27.235 LAYER ME2 ;
 ANTENNAMAXAREACAR                       28.835 LAYER ME3 ;
END A1
PIN A2
  DIRECTION INPUT ;
 PORT
  LAYER ME3 ;
  RECT 277.306 0.000 277.626 0.720 ;
  LAYER ME2 ;
  RECT 277.306 0.000 277.626 0.720 ;
  LAYER ME1 ;
  RECT 277.306 0.000 277.626 0.720 ;
 END
 ANTENNAPARTIALMETALAREA                  3.688 LAYER ME2 ;
 ANTENNAGATEAREA                          0.144 LAYER ME2 ;
 ANTENNAGATEAREA                          0.144 LAYER ME3 ;
 ANTENNADIFFAREA                          0.218 LAYER ME2 ;
 ANTENNADIFFAREA                          0.218 LAYER ME3 ;
 ANTENNAMAXAREACAR                       28.214 LAYER ME2 ;
 ANTENNAMAXAREACAR                       29.814 LAYER ME3 ;
END A2
PIN A3
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 270.488 0.000 270.808 0.720 ;
  LAYER ME3 ;
  RECT 270.488 0.000 270.808 0.720 ;
  LAYER ME2 ;
  RECT 270.488 0.000 270.808 0.720 ;
  LAYER ME1 ;
  RECT 270.488 0.000 270.808 0.720 ;
 END
 ANTENNAPARTIALMETALAREA                  4.391 LAYER ME2 ;
 ANTENNAGATEAREA                          0.180 LAYER ME2 ;
 ANTENNAGATEAREA                          0.180 LAYER ME3 ;
 ANTENNAGATEAREA                          0.180 LAYER ME4 ;
 ANTENNADIFFAREA                          0.218 LAYER ME2 ;
 ANTENNADIFFAREA                          0.218 LAYER ME3 ;
 ANTENNADIFFAREA                          0.218 LAYER ME4 ;
 ANTENNAMAXAREACAR                       27.451 LAYER ME2 ;
 ANTENNAMAXAREACAR                       28.731 LAYER ME3 ;
 ANTENNAMAXAREACAR                       30.011 LAYER ME4 ;
END A3
PIN A4
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 269.808 0.000 270.128 0.720 ;
  LAYER ME3 ;
  RECT 269.808 0.000 270.128 0.720 ;
  LAYER ME2 ;
  RECT 269.808 0.000 270.128 0.720 ;
  LAYER ME1 ;
  RECT 269.808 0.000 270.128 0.720 ;
 END
 ANTENNAPARTIALMETALAREA                  3.928 LAYER ME2 ;
 ANTENNAGATEAREA                          0.180 LAYER ME2 ;
 ANTENNAGATEAREA                          0.180 LAYER ME3 ;
 ANTENNAGATEAREA                          0.180 LAYER ME4 ;
 ANTENNADIFFAREA                          0.218 LAYER ME2 ;
 ANTENNADIFFAREA                          0.218 LAYER ME3 ;
 ANTENNADIFFAREA                          0.218 LAYER ME4 ;
 ANTENNAMAXAREACAR                       26.813 LAYER ME2 ;
 ANTENNAMAXAREACAR                       28.093 LAYER ME3 ;
 ANTENNAMAXAREACAR                       29.373 LAYER ME4 ;
END A4
PIN A5
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 266.328 0.000 266.648 0.720 ;
  LAYER ME3 ;
  RECT 266.328 0.000 266.648 0.720 ;
  LAYER ME2 ;
  RECT 266.328 0.000 266.648 0.720 ;
  LAYER ME1 ;
  RECT 266.328 0.000 266.648 0.720 ;
 END
 ANTENNAPARTIALMETALAREA                  4.391 LAYER ME2 ;
 ANTENNAGATEAREA                          0.180 LAYER ME2 ;
 ANTENNAGATEAREA                          0.180 LAYER ME3 ;
 ANTENNAGATEAREA                          0.180 LAYER ME4 ;
 ANTENNADIFFAREA                          0.218 LAYER ME2 ;
 ANTENNADIFFAREA                          0.218 LAYER ME3 ;
 ANTENNADIFFAREA                          0.218 LAYER ME4 ;
 ANTENNAMAXAREACAR                       27.451 LAYER ME2 ;
 ANTENNAMAXAREACAR                       28.731 LAYER ME3 ;
 ANTENNAMAXAREACAR                       30.011 LAYER ME4 ;
END A5
PIN A6
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 265.648 0.000 265.968 0.720 ;
  LAYER ME3 ;
  RECT 265.648 0.000 265.968 0.720 ;
  LAYER ME2 ;
  RECT 265.648 0.000 265.968 0.720 ;
  LAYER ME1 ;
  RECT 265.648 0.000 265.968 0.720 ;
 END
 ANTENNAPARTIALMETALAREA                  3.928 LAYER ME2 ;
 ANTENNAGATEAREA                          0.180 LAYER ME2 ;
 ANTENNAGATEAREA                          0.180 LAYER ME3 ;
 ANTENNAGATEAREA                          0.180 LAYER ME4 ;
 ANTENNADIFFAREA                          0.218 LAYER ME2 ;
 ANTENNADIFFAREA                          0.218 LAYER ME3 ;
 ANTENNADIFFAREA                          0.218 LAYER ME4 ;
 ANTENNAMAXAREACAR                       26.813 LAYER ME2 ;
 ANTENNAMAXAREACAR                       28.093 LAYER ME3 ;
 ANTENNAMAXAREACAR                       29.373 LAYER ME4 ;
END A6
PIN A7
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 262.168 0.000 262.488 0.720 ;
  LAYER ME3 ;
  RECT 262.168 0.000 262.488 0.720 ;
  LAYER ME2 ;
  RECT 262.168 0.000 262.488 0.720 ;
  LAYER ME1 ;
  RECT 262.168 0.000 262.488 0.720 ;
 END
 ANTENNAPARTIALMETALAREA                  4.391 LAYER ME2 ;
 ANTENNAGATEAREA                          0.180 LAYER ME2 ;
 ANTENNAGATEAREA                          0.180 LAYER ME3 ;
 ANTENNAGATEAREA                          0.180 LAYER ME4 ;
 ANTENNADIFFAREA                          0.218 LAYER ME2 ;
 ANTENNADIFFAREA                          0.218 LAYER ME3 ;
 ANTENNADIFFAREA                          0.218 LAYER ME4 ;
 ANTENNAMAXAREACAR                       27.451 LAYER ME2 ;
 ANTENNAMAXAREACAR                       28.731 LAYER ME3 ;
 ANTENNAMAXAREACAR                       30.011 LAYER ME4 ;
END A7
PIN A8
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 261.488 0.000 261.808 0.720 ;
  LAYER ME3 ;
  RECT 261.488 0.000 261.808 0.720 ;
  LAYER ME2 ;
  RECT 261.488 0.000 261.808 0.720 ;
  LAYER ME1 ;
  RECT 261.488 0.000 261.808 0.720 ;
 END
 ANTENNAPARTIALMETALAREA                  3.928 LAYER ME2 ;
 ANTENNAGATEAREA                          0.180 LAYER ME2 ;
 ANTENNAGATEAREA                          0.180 LAYER ME3 ;
 ANTENNAGATEAREA                          0.180 LAYER ME4 ;
 ANTENNADIFFAREA                          0.218 LAYER ME2 ;
 ANTENNADIFFAREA                          0.218 LAYER ME3 ;
 ANTENNADIFFAREA                          0.218 LAYER ME4 ;
 ANTENNAMAXAREACAR                       26.813 LAYER ME2 ;
 ANTENNAMAXAREACAR                       28.093 LAYER ME3 ;
 ANTENNAMAXAREACAR                       29.373 LAYER ME4 ;
END A8
PIN A0
  DIRECTION INPUT ;
 PORT
  LAYER ME3 ;
  RECT 287.322 0.000 287.642 0.662 ;
  LAYER ME2 ;
  RECT 287.322 0.000 287.642 0.662 ;
  LAYER ME1 ;
  RECT 287.322 0.000 287.642 0.662 ;
 END
 ANTENNAPARTIALMETALAREA                  5.907 LAYER ME2 ;
 ANTENNAGATEAREA                          0.108 LAYER ME2 ;
 ANTENNAGATEAREA                          0.108 LAYER ME3 ;
 ANTENNADIFFAREA                          0.218 LAYER ME2 ;
 ANTENNADIFFAREA                          0.218 LAYER ME3 ;
 ANTENNAMAXAREACAR                       58.521 LAYER ME2 ;
 ANTENNAMAXAREACAR                       60.482 LAYER ME3 ;
END A0
PIN DVSE
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 296.913 0.000 297.233 0.720 ;
  LAYER ME3 ;
  RECT 296.913 0.000 297.233 0.720 ;
  LAYER ME3 ;
  RECT 296.913 0.000 297.233 0.720 ;
  LAYER ME2 ;
  RECT 296.913 0.000 297.233 0.720 ;
  LAYER ME2 ;
  RECT 296.913 0.000 297.233 0.720 ;
  LAYER ME1 ;
  RECT 296.913 0.000 297.233 0.720 ;
  LAYER ME1 ;
  RECT 296.913 0.000 297.233 0.720 ;
 END
 ANTENNAPARTIALMETALAREA                  7.809 LAYER ME2 ;
 ANTENNAGATEAREA                          0.612 LAYER ME2 ;
 ANTENNAGATEAREA                          0.612 LAYER ME3 ;
 ANTENNAGATEAREA                          0.612 LAYER ME4 ;
 ANTENNADIFFAREA                          0.218 LAYER ME2 ;
 ANTENNADIFFAREA                          0.218 LAYER ME3 ;
 ANTENNADIFFAREA                          0.218 LAYER ME4 ;
 ANTENNAMAXAREACAR                       76.330 LAYER ME2 ;
 ANTENNAMAXAREACAR                       78.463 LAYER ME3 ;
 ANTENNAMAXAREACAR                       80.596 LAYER ME4 ;
END DVSE
PIN DVS3
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 296.393 0.000 296.713 0.720 ;
  LAYER ME3 ;
  RECT 296.393 0.000 296.713 0.720 ;
  LAYER ME3 ;
  RECT 296.393 0.000 296.713 0.720 ;
  LAYER ME2 ;
  RECT 296.393 0.000 296.713 0.720 ;
  LAYER ME2 ;
  RECT 296.393 0.000 296.713 0.720 ;
  LAYER ME1 ;
  RECT 296.393 0.000 296.713 0.720 ;
  LAYER ME1 ;
  RECT 296.393 0.000 296.713 0.720 ;
 END
 ANTENNAPARTIALMETALAREA                  6.179 LAYER ME2 ;
 ANTENNAGATEAREA                          0.108 LAYER ME2 ;
 ANTENNAGATEAREA                          0.108 LAYER ME3 ;
 ANTENNAGATEAREA                          0.108 LAYER ME4 ;
 ANTENNADIFFAREA                          0.218 LAYER ME2 ;
 ANTENNADIFFAREA                          0.218 LAYER ME3 ;
 ANTENNADIFFAREA                          0.218 LAYER ME4 ;
 ANTENNAMAXAREACAR                       68.823 LAYER ME2 ;
 ANTENNAMAXAREACAR                       70.956 LAYER ME3 ;
 ANTENNAMAXAREACAR                       73.089 LAYER ME4 ;
END DVS3
PIN DVS2
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 297.433 0.000 297.753 0.720 ;
  LAYER ME3 ;
  RECT 297.433 0.000 297.753 0.720 ;
  LAYER ME3 ;
  RECT 297.433 0.000 297.753 0.720 ;
  LAYER ME2 ;
  RECT 297.433 0.000 297.753 0.720 ;
  LAYER ME2 ;
  RECT 297.433 0.000 297.753 0.720 ;
  LAYER ME1 ;
  RECT 297.433 0.000 297.753 0.720 ;
  LAYER ME1 ;
  RECT 297.433 0.000 297.753 0.720 ;
 END
 ANTENNAPARTIALMETALAREA                  7.876 LAYER ME2 ;
 ANTENNAGATEAREA                          0.108 LAYER ME2 ;
 ANTENNAGATEAREA                          0.108 LAYER ME3 ;
 ANTENNAGATEAREA                          0.108 LAYER ME4 ;
 ANTENNADIFFAREA                          0.218 LAYER ME2 ;
 ANTENNADIFFAREA                          0.218 LAYER ME3 ;
 ANTENNADIFFAREA                          0.218 LAYER ME4 ;
 ANTENNAMAXAREACAR                       83.257 LAYER ME2 ;
 ANTENNAMAXAREACAR                       85.391 LAYER ME3 ;
 ANTENNAMAXAREACAR                       87.524 LAYER ME4 ;
END DVS2
PIN DVS1
  DIRECTION INPUT ;
 PORT
  LAYER ME3 ;
  RECT 293.777 0.000 294.097 0.720 ;
  LAYER ME2 ;
  RECT 293.777 0.000 294.097 0.720 ;
  LAYER ME1 ;
  RECT 293.777 0.000 294.097 0.720 ;
 END
 ANTENNAPARTIALMETALAREA                  6.247 LAYER ME2 ;
 ANTENNAGATEAREA                          0.108 LAYER ME2 ;
 ANTENNAGATEAREA                          0.108 LAYER ME3 ;
 ANTENNADIFFAREA                          0.218 LAYER ME2 ;
 ANTENNADIFFAREA                          0.218 LAYER ME3 ;
 ANTENNAMAXAREACAR                       69.294 LAYER ME2 ;
 ANTENNAMAXAREACAR                       71.427 LAYER ME3 ;
END DVS1
PIN DVS0
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 297.953 0.000 298.273 0.720 ;
  LAYER ME3 ;
  RECT 297.953 0.000 298.273 0.720 ;
  LAYER ME3 ;
  RECT 297.953 0.000 298.273 0.720 ;
  LAYER ME2 ;
  RECT 297.953 0.000 298.273 0.720 ;
  LAYER ME2 ;
  RECT 297.953 0.000 298.273 0.720 ;
  LAYER ME1 ;
  RECT 297.953 0.000 298.273 0.720 ;
  LAYER ME1 ;
  RECT 297.953 0.000 298.273 0.720 ;
 END
 ANTENNAPARTIALMETALAREA                  7.119 LAYER ME2 ;
 ANTENNAGATEAREA                          0.108 LAYER ME2 ;
 ANTENNAGATEAREA                          0.108 LAYER ME3 ;
 ANTENNAGATEAREA                          0.108 LAYER ME4 ;
 ANTENNADIFFAREA                          0.218 LAYER ME2 ;
 ANTENNADIFFAREA                          0.218 LAYER ME3 ;
 ANTENNADIFFAREA                          0.218 LAYER ME4 ;
 ANTENNAMAXAREACAR                       77.987 LAYER ME2 ;
 ANTENNAMAXAREACAR                       80.120 LAYER ME3 ;
 ANTENNAMAXAREACAR                       82.254 LAYER ME4 ;
END DVS0
PIN CK
  DIRECTION INPUT ;
 PORT
  LAYER ME3 ;
  RECT 289.861 0.000 290.181 0.720 ;
  LAYER ME2 ;
  RECT 289.861 0.000 290.181 0.720 ;
  LAYER ME1 ;
  RECT 289.861 0.000 290.181 0.720 ;
 END
 ANTENNAPARTIALMETALAREA                  5.257 LAYER ME2 ;
 ANTENNAPARTIALMETALAREA                  8.004 LAYER ME3 ;
 ANTENNAGATEAREA                          0.072 LAYER ME2 ;
 ANTENNAGATEAREA                          1.296 LAYER ME3 ;
 ANTENNADIFFAREA                          0.218 LAYER ME2 ;
 ANTENNADIFFAREA                          0.218 LAYER ME3 ;
 ANTENNAMAXAREACAR                       86.308 LAYER ME2 ;
 ANTENNAMAXAREACAR                      200.681 LAYER ME3 ;
END CK
PIN CSB
  DIRECTION INPUT ;
 PORT
  LAYER ME3 ;
  RECT 281.247 0.000 281.567 0.720 ;
  LAYER ME2 ;
  RECT 281.247 0.000 281.567 0.720 ;
  LAYER ME1 ;
  RECT 281.247 0.000 281.567 0.720 ;
 END
 ANTENNAPARTIALMETALAREA                  5.788 LAYER ME2 ;
 ANTENNAPARTIALMETALAREA                  8.036 LAYER ME3 ;
 ANTENNAGATEAREA                          2.508 LAYER ME2 ;
 ANTENNAGATEAREA                          3.732 LAYER ME3 ;
 ANTENNADIFFAREA                          0.218 LAYER ME2 ;
 ANTENNADIFFAREA                          0.218 LAYER ME3 ;
 ANTENNAMAXAREACAR                        3.046 LAYER ME2 ;
 ANTENNAMAXAREACAR                       40.545 LAYER ME3 ;
END CSB
PIN DI127
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 552.819 0.000 553.139 0.600 ;
  LAYER ME3 ;
  RECT 552.819 0.000 553.139 0.600 ;
  LAYER ME2 ;
  RECT 552.819 0.000 553.139 0.600 ;
  LAYER ME1 ;
  RECT 552.819 0.000 553.139 0.600 ;
 END
 ANTENNAPARTIALMETALAREA                  1.058 LAYER ME2 ;
 ANTENNAGATEAREA                          0.072 LAYER ME2 ;
 ANTENNAGATEAREA                          0.072 LAYER ME3 ;
 ANTENNAGATEAREA                          0.072 LAYER ME4 ;
 ANTENNADIFFAREA                          0.160 LAYER ME2 ;
 ANTENNADIFFAREA                          0.160 LAYER ME3 ;
 ANTENNADIFFAREA                          0.160 LAYER ME4 ;
 ANTENNAMAXAREACAR                       21.782 LAYER ME2 ;
 ANTENNAMAXAREACAR                       24.449 LAYER ME3 ;
 ANTENNAMAXAREACAR                       27.116 LAYER ME4 ;
END DI127
PIN DO127
  DIRECTION OUTPUT ;
 PORT
  LAYER ME4 ;
  RECT 552.257 0.000 552.577 0.600 ;
  LAYER ME3 ;
  RECT 552.257 0.000 552.577 0.600 ;
  LAYER ME2 ;
  RECT 552.257 0.000 552.577 0.600 ;
  LAYER ME1 ;
  RECT 552.257 0.000 552.577 0.600 ;
 END
 ANTENNAPARTIALMETALAREA                  5.273 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME3 ;
 ANTENNADIFFAREA                          1.293 LAYER ME4 ;
END DO127
PIN DI126
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 548.815 0.000 549.135 0.600 ;
  LAYER ME3 ;
  RECT 548.815 0.000 549.135 0.600 ;
  LAYER ME2 ;
  RECT 548.815 0.000 549.135 0.600 ;
  LAYER ME1 ;
  RECT 548.815 0.000 549.135 0.600 ;
 END
 ANTENNAPARTIALMETALAREA                  1.058 LAYER ME2 ;
 ANTENNAGATEAREA                          0.072 LAYER ME2 ;
 ANTENNAGATEAREA                          0.072 LAYER ME3 ;
 ANTENNAGATEAREA                          0.072 LAYER ME4 ;
 ANTENNADIFFAREA                          0.160 LAYER ME2 ;
 ANTENNADIFFAREA                          0.160 LAYER ME3 ;
 ANTENNADIFFAREA                          0.160 LAYER ME4 ;
 ANTENNAMAXAREACAR                       21.782 LAYER ME2 ;
 ANTENNAMAXAREACAR                       24.449 LAYER ME3 ;
 ANTENNAMAXAREACAR                       27.116 LAYER ME4 ;
END DI126
PIN DO126
  DIRECTION OUTPUT ;
 PORT
  LAYER ME4 ;
  RECT 548.253 0.000 548.573 0.600 ;
  LAYER ME3 ;
  RECT 548.253 0.000 548.573 0.600 ;
  LAYER ME2 ;
  RECT 548.253 0.000 548.573 0.600 ;
  LAYER ME1 ;
  RECT 548.253 0.000 548.573 0.600 ;
 END
 ANTENNAPARTIALMETALAREA                  5.273 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME3 ;
 ANTENNADIFFAREA                          1.293 LAYER ME4 ;
END DO126
PIN DI125
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 544.811 0.000 545.131 0.600 ;
  LAYER ME3 ;
  RECT 544.811 0.000 545.131 0.600 ;
  LAYER ME2 ;
  RECT 544.811 0.000 545.131 0.600 ;
  LAYER ME1 ;
  RECT 544.811 0.000 545.131 0.600 ;
 END
 ANTENNAPARTIALMETALAREA                  1.058 LAYER ME2 ;
 ANTENNAGATEAREA                          0.072 LAYER ME2 ;
 ANTENNAGATEAREA                          0.072 LAYER ME3 ;
 ANTENNAGATEAREA                          0.072 LAYER ME4 ;
 ANTENNADIFFAREA                          0.160 LAYER ME2 ;
 ANTENNADIFFAREA                          0.160 LAYER ME3 ;
 ANTENNADIFFAREA                          0.160 LAYER ME4 ;
 ANTENNAMAXAREACAR                       21.782 LAYER ME2 ;
 ANTENNAMAXAREACAR                       24.449 LAYER ME3 ;
 ANTENNAMAXAREACAR                       27.116 LAYER ME4 ;
END DI125
PIN DO125
  DIRECTION OUTPUT ;
 PORT
  LAYER ME4 ;
  RECT 544.249 0.000 544.569 0.600 ;
  LAYER ME3 ;
  RECT 544.249 0.000 544.569 0.600 ;
  LAYER ME2 ;
  RECT 544.249 0.000 544.569 0.600 ;
  LAYER ME1 ;
  RECT 544.249 0.000 544.569 0.600 ;
 END
 ANTENNAPARTIALMETALAREA                  5.273 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME3 ;
 ANTENNADIFFAREA                          1.293 LAYER ME4 ;
END DO125
PIN DI124
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 540.807 0.000 541.127 0.600 ;
  LAYER ME3 ;
  RECT 540.807 0.000 541.127 0.600 ;
  LAYER ME2 ;
  RECT 540.807 0.000 541.127 0.600 ;
  LAYER ME1 ;
  RECT 540.807 0.000 541.127 0.600 ;
 END
 ANTENNAPARTIALMETALAREA                  1.058 LAYER ME2 ;
 ANTENNAGATEAREA                          0.072 LAYER ME2 ;
 ANTENNAGATEAREA                          0.072 LAYER ME3 ;
 ANTENNAGATEAREA                          0.072 LAYER ME4 ;
 ANTENNADIFFAREA                          0.160 LAYER ME2 ;
 ANTENNADIFFAREA                          0.160 LAYER ME3 ;
 ANTENNADIFFAREA                          0.160 LAYER ME4 ;
 ANTENNAMAXAREACAR                       21.782 LAYER ME2 ;
 ANTENNAMAXAREACAR                       24.449 LAYER ME3 ;
 ANTENNAMAXAREACAR                       27.116 LAYER ME4 ;
END DI124
PIN DO124
  DIRECTION OUTPUT ;
 PORT
  LAYER ME4 ;
  RECT 540.245 0.000 540.565 0.600 ;
  LAYER ME3 ;
  RECT 540.245 0.000 540.565 0.600 ;
  LAYER ME2 ;
  RECT 540.245 0.000 540.565 0.600 ;
  LAYER ME1 ;
  RECT 540.245 0.000 540.565 0.600 ;
 END
 ANTENNAPARTIALMETALAREA                  5.273 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME3 ;
 ANTENNADIFFAREA                          1.293 LAYER ME4 ;
END DO124
PIN DI123
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 536.803 0.000 537.123 0.600 ;
  LAYER ME3 ;
  RECT 536.803 0.000 537.123 0.600 ;
  LAYER ME2 ;
  RECT 536.803 0.000 537.123 0.600 ;
  LAYER ME1 ;
  RECT 536.803 0.000 537.123 0.600 ;
 END
 ANTENNAPARTIALMETALAREA                  1.058 LAYER ME2 ;
 ANTENNAGATEAREA                          0.072 LAYER ME2 ;
 ANTENNAGATEAREA                          0.072 LAYER ME3 ;
 ANTENNAGATEAREA                          0.072 LAYER ME4 ;
 ANTENNADIFFAREA                          0.160 LAYER ME2 ;
 ANTENNADIFFAREA                          0.160 LAYER ME3 ;
 ANTENNADIFFAREA                          0.160 LAYER ME4 ;
 ANTENNAMAXAREACAR                       21.782 LAYER ME2 ;
 ANTENNAMAXAREACAR                       24.449 LAYER ME3 ;
 ANTENNAMAXAREACAR                       27.116 LAYER ME4 ;
END DI123
PIN DO123
  DIRECTION OUTPUT ;
 PORT
  LAYER ME4 ;
  RECT 536.241 0.000 536.561 0.600 ;
  LAYER ME3 ;
  RECT 536.241 0.000 536.561 0.600 ;
  LAYER ME2 ;
  RECT 536.241 0.000 536.561 0.600 ;
  LAYER ME1 ;
  RECT 536.241 0.000 536.561 0.600 ;
 END
 ANTENNAPARTIALMETALAREA                  5.273 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME3 ;
 ANTENNADIFFAREA                          1.293 LAYER ME4 ;
END DO123
PIN DI122
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 532.799 0.000 533.119 0.600 ;
  LAYER ME3 ;
  RECT 532.799 0.000 533.119 0.600 ;
  LAYER ME2 ;
  RECT 532.799 0.000 533.119 0.600 ;
  LAYER ME1 ;
  RECT 532.799 0.000 533.119 0.600 ;
 END
 ANTENNAPARTIALMETALAREA                  1.058 LAYER ME2 ;
 ANTENNAGATEAREA                          0.072 LAYER ME2 ;
 ANTENNAGATEAREA                          0.072 LAYER ME3 ;
 ANTENNAGATEAREA                          0.072 LAYER ME4 ;
 ANTENNADIFFAREA                          0.160 LAYER ME2 ;
 ANTENNADIFFAREA                          0.160 LAYER ME3 ;
 ANTENNADIFFAREA                          0.160 LAYER ME4 ;
 ANTENNAMAXAREACAR                       21.782 LAYER ME2 ;
 ANTENNAMAXAREACAR                       24.449 LAYER ME3 ;
 ANTENNAMAXAREACAR                       27.116 LAYER ME4 ;
END DI122
PIN DO122
  DIRECTION OUTPUT ;
 PORT
  LAYER ME4 ;
  RECT 532.237 0.000 532.557 0.600 ;
  LAYER ME3 ;
  RECT 532.237 0.000 532.557 0.600 ;
  LAYER ME2 ;
  RECT 532.237 0.000 532.557 0.600 ;
  LAYER ME1 ;
  RECT 532.237 0.000 532.557 0.600 ;
 END
 ANTENNAPARTIALMETALAREA                  5.273 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME3 ;
 ANTENNADIFFAREA                          1.293 LAYER ME4 ;
END DO122
PIN DI121
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 528.795 0.000 529.115 0.600 ;
  LAYER ME3 ;
  RECT 528.795 0.000 529.115 0.600 ;
  LAYER ME2 ;
  RECT 528.795 0.000 529.115 0.600 ;
  LAYER ME1 ;
  RECT 528.795 0.000 529.115 0.600 ;
 END
 ANTENNAPARTIALMETALAREA                  1.058 LAYER ME2 ;
 ANTENNAGATEAREA                          0.072 LAYER ME2 ;
 ANTENNAGATEAREA                          0.072 LAYER ME3 ;
 ANTENNAGATEAREA                          0.072 LAYER ME4 ;
 ANTENNADIFFAREA                          0.160 LAYER ME2 ;
 ANTENNADIFFAREA                          0.160 LAYER ME3 ;
 ANTENNADIFFAREA                          0.160 LAYER ME4 ;
 ANTENNAMAXAREACAR                       21.782 LAYER ME2 ;
 ANTENNAMAXAREACAR                       24.449 LAYER ME3 ;
 ANTENNAMAXAREACAR                       27.116 LAYER ME4 ;
END DI121
PIN DO121
  DIRECTION OUTPUT ;
 PORT
  LAYER ME4 ;
  RECT 528.233 0.000 528.553 0.600 ;
  LAYER ME3 ;
  RECT 528.233 0.000 528.553 0.600 ;
  LAYER ME2 ;
  RECT 528.233 0.000 528.553 0.600 ;
  LAYER ME1 ;
  RECT 528.233 0.000 528.553 0.600 ;
 END
 ANTENNAPARTIALMETALAREA                  5.273 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME3 ;
 ANTENNADIFFAREA                          1.293 LAYER ME4 ;
END DO121
PIN DI120
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 524.791 0.000 525.111 0.600 ;
  LAYER ME3 ;
  RECT 524.791 0.000 525.111 0.600 ;
  LAYER ME2 ;
  RECT 524.791 0.000 525.111 0.600 ;
  LAYER ME1 ;
  RECT 524.791 0.000 525.111 0.600 ;
 END
 ANTENNAPARTIALMETALAREA                  1.058 LAYER ME2 ;
 ANTENNAGATEAREA                          0.072 LAYER ME2 ;
 ANTENNAGATEAREA                          0.072 LAYER ME3 ;
 ANTENNAGATEAREA                          0.072 LAYER ME4 ;
 ANTENNADIFFAREA                          0.160 LAYER ME2 ;
 ANTENNADIFFAREA                          0.160 LAYER ME3 ;
 ANTENNADIFFAREA                          0.160 LAYER ME4 ;
 ANTENNAMAXAREACAR                       21.782 LAYER ME2 ;
 ANTENNAMAXAREACAR                       24.449 LAYER ME3 ;
 ANTENNAMAXAREACAR                       27.116 LAYER ME4 ;
END DI120
PIN DO120
  DIRECTION OUTPUT ;
 PORT
  LAYER ME4 ;
  RECT 524.229 0.000 524.549 0.600 ;
  LAYER ME3 ;
  RECT 524.229 0.000 524.549 0.600 ;
  LAYER ME2 ;
  RECT 524.229 0.000 524.549 0.600 ;
  LAYER ME1 ;
  RECT 524.229 0.000 524.549 0.600 ;
 END
 ANTENNAPARTIALMETALAREA                  5.273 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME3 ;
 ANTENNADIFFAREA                          1.293 LAYER ME4 ;
END DO120
PIN DI119
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 520.787 0.000 521.107 0.600 ;
  LAYER ME3 ;
  RECT 520.787 0.000 521.107 0.600 ;
  LAYER ME2 ;
  RECT 520.787 0.000 521.107 0.600 ;
  LAYER ME1 ;
  RECT 520.787 0.000 521.107 0.600 ;
 END
 ANTENNAPARTIALMETALAREA                  1.058 LAYER ME2 ;
 ANTENNAGATEAREA                          0.072 LAYER ME2 ;
 ANTENNAGATEAREA                          0.072 LAYER ME3 ;
 ANTENNAGATEAREA                          0.072 LAYER ME4 ;
 ANTENNADIFFAREA                          0.160 LAYER ME2 ;
 ANTENNADIFFAREA                          0.160 LAYER ME3 ;
 ANTENNADIFFAREA                          0.160 LAYER ME4 ;
 ANTENNAMAXAREACAR                       21.782 LAYER ME2 ;
 ANTENNAMAXAREACAR                       24.449 LAYER ME3 ;
 ANTENNAMAXAREACAR                       27.116 LAYER ME4 ;
END DI119
PIN DO119
  DIRECTION OUTPUT ;
 PORT
  LAYER ME4 ;
  RECT 520.225 0.000 520.545 0.600 ;
  LAYER ME3 ;
  RECT 520.225 0.000 520.545 0.600 ;
  LAYER ME2 ;
  RECT 520.225 0.000 520.545 0.600 ;
  LAYER ME1 ;
  RECT 520.225 0.000 520.545 0.600 ;
 END
 ANTENNAPARTIALMETALAREA                  5.273 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME3 ;
 ANTENNADIFFAREA                          1.293 LAYER ME4 ;
END DO119
PIN DI118
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 516.783 0.000 517.103 0.600 ;
  LAYER ME3 ;
  RECT 516.783 0.000 517.103 0.600 ;
  LAYER ME2 ;
  RECT 516.783 0.000 517.103 0.600 ;
  LAYER ME1 ;
  RECT 516.783 0.000 517.103 0.600 ;
 END
 ANTENNAPARTIALMETALAREA                  1.058 LAYER ME2 ;
 ANTENNAGATEAREA                          0.072 LAYER ME2 ;
 ANTENNAGATEAREA                          0.072 LAYER ME3 ;
 ANTENNAGATEAREA                          0.072 LAYER ME4 ;
 ANTENNADIFFAREA                          0.160 LAYER ME2 ;
 ANTENNADIFFAREA                          0.160 LAYER ME3 ;
 ANTENNADIFFAREA                          0.160 LAYER ME4 ;
 ANTENNAMAXAREACAR                       21.782 LAYER ME2 ;
 ANTENNAMAXAREACAR                       24.449 LAYER ME3 ;
 ANTENNAMAXAREACAR                       27.116 LAYER ME4 ;
END DI118
PIN DO118
  DIRECTION OUTPUT ;
 PORT
  LAYER ME4 ;
  RECT 516.221 0.000 516.541 0.600 ;
  LAYER ME3 ;
  RECT 516.221 0.000 516.541 0.600 ;
  LAYER ME2 ;
  RECT 516.221 0.000 516.541 0.600 ;
  LAYER ME1 ;
  RECT 516.221 0.000 516.541 0.600 ;
 END
 ANTENNAPARTIALMETALAREA                  5.273 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME3 ;
 ANTENNADIFFAREA                          1.293 LAYER ME4 ;
END DO118
PIN DI117
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 512.779 0.000 513.099 0.600 ;
  LAYER ME3 ;
  RECT 512.779 0.000 513.099 0.600 ;
  LAYER ME2 ;
  RECT 512.779 0.000 513.099 0.600 ;
  LAYER ME1 ;
  RECT 512.779 0.000 513.099 0.600 ;
 END
 ANTENNAPARTIALMETALAREA                  1.058 LAYER ME2 ;
 ANTENNAGATEAREA                          0.072 LAYER ME2 ;
 ANTENNAGATEAREA                          0.072 LAYER ME3 ;
 ANTENNAGATEAREA                          0.072 LAYER ME4 ;
 ANTENNADIFFAREA                          0.160 LAYER ME2 ;
 ANTENNADIFFAREA                          0.160 LAYER ME3 ;
 ANTENNADIFFAREA                          0.160 LAYER ME4 ;
 ANTENNAMAXAREACAR                       21.782 LAYER ME2 ;
 ANTENNAMAXAREACAR                       24.449 LAYER ME3 ;
 ANTENNAMAXAREACAR                       27.116 LAYER ME4 ;
END DI117
PIN DO117
  DIRECTION OUTPUT ;
 PORT
  LAYER ME4 ;
  RECT 512.217 0.000 512.537 0.600 ;
  LAYER ME3 ;
  RECT 512.217 0.000 512.537 0.600 ;
  LAYER ME2 ;
  RECT 512.217 0.000 512.537 0.600 ;
  LAYER ME1 ;
  RECT 512.217 0.000 512.537 0.600 ;
 END
 ANTENNAPARTIALMETALAREA                  5.273 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME3 ;
 ANTENNADIFFAREA                          1.293 LAYER ME4 ;
END DO117
PIN DI116
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 508.775 0.000 509.095 0.600 ;
  LAYER ME3 ;
  RECT 508.775 0.000 509.095 0.600 ;
  LAYER ME2 ;
  RECT 508.775 0.000 509.095 0.600 ;
  LAYER ME1 ;
  RECT 508.775 0.000 509.095 0.600 ;
 END
 ANTENNAPARTIALMETALAREA                  1.058 LAYER ME2 ;
 ANTENNAGATEAREA                          0.072 LAYER ME2 ;
 ANTENNAGATEAREA                          0.072 LAYER ME3 ;
 ANTENNAGATEAREA                          0.072 LAYER ME4 ;
 ANTENNADIFFAREA                          0.160 LAYER ME2 ;
 ANTENNADIFFAREA                          0.160 LAYER ME3 ;
 ANTENNADIFFAREA                          0.160 LAYER ME4 ;
 ANTENNAMAXAREACAR                       21.782 LAYER ME2 ;
 ANTENNAMAXAREACAR                       24.449 LAYER ME3 ;
 ANTENNAMAXAREACAR                       27.116 LAYER ME4 ;
END DI116
PIN DO116
  DIRECTION OUTPUT ;
 PORT
  LAYER ME4 ;
  RECT 508.213 0.000 508.533 0.600 ;
  LAYER ME3 ;
  RECT 508.213 0.000 508.533 0.600 ;
  LAYER ME2 ;
  RECT 508.213 0.000 508.533 0.600 ;
  LAYER ME1 ;
  RECT 508.213 0.000 508.533 0.600 ;
 END
 ANTENNAPARTIALMETALAREA                  5.273 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME3 ;
 ANTENNADIFFAREA                          1.293 LAYER ME4 ;
END DO116
PIN DI115
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 504.771 0.000 505.091 0.600 ;
  LAYER ME3 ;
  RECT 504.771 0.000 505.091 0.600 ;
  LAYER ME2 ;
  RECT 504.771 0.000 505.091 0.600 ;
  LAYER ME1 ;
  RECT 504.771 0.000 505.091 0.600 ;
 END
 ANTENNAPARTIALMETALAREA                  1.058 LAYER ME2 ;
 ANTENNAGATEAREA                          0.072 LAYER ME2 ;
 ANTENNAGATEAREA                          0.072 LAYER ME3 ;
 ANTENNAGATEAREA                          0.072 LAYER ME4 ;
 ANTENNADIFFAREA                          0.160 LAYER ME2 ;
 ANTENNADIFFAREA                          0.160 LAYER ME3 ;
 ANTENNADIFFAREA                          0.160 LAYER ME4 ;
 ANTENNAMAXAREACAR                       21.782 LAYER ME2 ;
 ANTENNAMAXAREACAR                       24.449 LAYER ME3 ;
 ANTENNAMAXAREACAR                       27.116 LAYER ME4 ;
END DI115
PIN DO115
  DIRECTION OUTPUT ;
 PORT
  LAYER ME4 ;
  RECT 504.209 0.000 504.529 0.600 ;
  LAYER ME3 ;
  RECT 504.209 0.000 504.529 0.600 ;
  LAYER ME2 ;
  RECT 504.209 0.000 504.529 0.600 ;
  LAYER ME1 ;
  RECT 504.209 0.000 504.529 0.600 ;
 END
 ANTENNAPARTIALMETALAREA                  5.273 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME3 ;
 ANTENNADIFFAREA                          1.293 LAYER ME4 ;
END DO115
PIN DI114
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 500.767 0.000 501.087 0.600 ;
  LAYER ME3 ;
  RECT 500.767 0.000 501.087 0.600 ;
  LAYER ME2 ;
  RECT 500.767 0.000 501.087 0.600 ;
  LAYER ME1 ;
  RECT 500.767 0.000 501.087 0.600 ;
 END
 ANTENNAPARTIALMETALAREA                  1.058 LAYER ME2 ;
 ANTENNAGATEAREA                          0.072 LAYER ME2 ;
 ANTENNAGATEAREA                          0.072 LAYER ME3 ;
 ANTENNAGATEAREA                          0.072 LAYER ME4 ;
 ANTENNADIFFAREA                          0.160 LAYER ME2 ;
 ANTENNADIFFAREA                          0.160 LAYER ME3 ;
 ANTENNADIFFAREA                          0.160 LAYER ME4 ;
 ANTENNAMAXAREACAR                       21.782 LAYER ME2 ;
 ANTENNAMAXAREACAR                       24.449 LAYER ME3 ;
 ANTENNAMAXAREACAR                       27.116 LAYER ME4 ;
END DI114
PIN DO114
  DIRECTION OUTPUT ;
 PORT
  LAYER ME4 ;
  RECT 500.205 0.000 500.525 0.600 ;
  LAYER ME3 ;
  RECT 500.205 0.000 500.525 0.600 ;
  LAYER ME2 ;
  RECT 500.205 0.000 500.525 0.600 ;
  LAYER ME1 ;
  RECT 500.205 0.000 500.525 0.600 ;
 END
 ANTENNAPARTIALMETALAREA                  5.273 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME3 ;
 ANTENNADIFFAREA                          1.293 LAYER ME4 ;
END DO114
PIN DI113
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 496.763 0.000 497.083 0.600 ;
  LAYER ME3 ;
  RECT 496.763 0.000 497.083 0.600 ;
  LAYER ME2 ;
  RECT 496.763 0.000 497.083 0.600 ;
  LAYER ME1 ;
  RECT 496.763 0.000 497.083 0.600 ;
 END
 ANTENNAPARTIALMETALAREA                  1.058 LAYER ME2 ;
 ANTENNAGATEAREA                          0.072 LAYER ME2 ;
 ANTENNAGATEAREA                          0.072 LAYER ME3 ;
 ANTENNAGATEAREA                          0.072 LAYER ME4 ;
 ANTENNADIFFAREA                          0.160 LAYER ME2 ;
 ANTENNADIFFAREA                          0.160 LAYER ME3 ;
 ANTENNADIFFAREA                          0.160 LAYER ME4 ;
 ANTENNAMAXAREACAR                       21.782 LAYER ME2 ;
 ANTENNAMAXAREACAR                       24.449 LAYER ME3 ;
 ANTENNAMAXAREACAR                       27.116 LAYER ME4 ;
END DI113
PIN DO113
  DIRECTION OUTPUT ;
 PORT
  LAYER ME4 ;
  RECT 496.201 0.000 496.521 0.600 ;
  LAYER ME3 ;
  RECT 496.201 0.000 496.521 0.600 ;
  LAYER ME2 ;
  RECT 496.201 0.000 496.521 0.600 ;
  LAYER ME1 ;
  RECT 496.201 0.000 496.521 0.600 ;
 END
 ANTENNAPARTIALMETALAREA                  5.273 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME3 ;
 ANTENNADIFFAREA                          1.293 LAYER ME4 ;
END DO113
PIN DI112
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 492.197 0.000 492.517 0.600 ;
  LAYER ME3 ;
  RECT 492.197 0.000 492.517 0.600 ;
  LAYER ME2 ;
  RECT 492.197 0.000 492.517 0.600 ;
  LAYER ME1 ;
  RECT 492.197 0.000 492.517 0.600 ;
 END
 ANTENNAPARTIALMETALAREA                  0.346 LAYER ME1 ;
 ANTENNAPARTIALMETALAREA                  1.466 LAYER ME2 ;
 ANTENNAPARTIALMETALAREA                  0.508 LAYER ME3 ;
 ANTENNAGATEAREA                          0.072 LAYER ME3 ;
 ANTENNAGATEAREA                          0.072 LAYER ME4 ;
 ANTENNADIFFAREA                          0.218 LAYER ME1 ;
 ANTENNADIFFAREA                          0.218 LAYER ME2 ;
 ANTENNADIFFAREA                          0.218 LAYER ME3 ;
 ANTENNADIFFAREA                          0.218 LAYER ME4 ;
 ANTENNAMAXAREACAR                       17.267 LAYER ME3 ;
 ANTENNAMAXAREACAR                       19.933 LAYER ME4 ;
END DI112
PIN DO112
  DIRECTION OUTPUT ;
 PORT
  LAYER ME4 ;
  RECT 492.759 0.000 493.079 0.600 ;
  LAYER ME3 ;
  RECT 492.759 0.000 493.079 0.600 ;
  LAYER ME2 ;
  RECT 492.759 0.000 493.079 0.600 ;
  LAYER ME1 ;
  RECT 492.759 0.000 493.079 0.600 ;
 END
 ANTENNAPARTIALMETALAREA                  5.602 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME3 ;
 ANTENNADIFFAREA                          1.293 LAYER ME4 ;
END DO112
PIN WEB7
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 490.757 0.000 491.077 0.600 ;
  LAYER ME3 ;
  RECT 490.757 0.000 491.077 0.600 ;
  LAYER ME2 ;
  RECT 490.757 0.000 491.077 0.600 ;
  LAYER ME1 ;
  RECT 490.757 0.000 491.077 0.600 ;
 END
 ANTENNAPARTIALMETALAREA                  1.036 LAYER ME2 ;
 ANTENNAGATEAREA                          0.288 LAYER ME2 ;
 ANTENNAGATEAREA                          0.288 LAYER ME3 ;
 ANTENNAGATEAREA                          0.288 LAYER ME4 ;
 ANTENNADIFFAREA                          0.206 LAYER ME2 ;
 ANTENNADIFFAREA                          0.206 LAYER ME3 ;
 ANTENNADIFFAREA                          0.206 LAYER ME4 ;
 ANTENNAMAXAREACAR                        5.844 LAYER ME2 ;
 ANTENNAMAXAREACAR                        6.511 LAYER ME3 ;
 ANTENNAMAXAREACAR                        7.178 LAYER ME4 ;
END WEB7
PIN DI111
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 488.755 0.000 489.075 0.600 ;
  LAYER ME3 ;
  RECT 488.755 0.000 489.075 0.600 ;
  LAYER ME2 ;
  RECT 488.755 0.000 489.075 0.600 ;
  LAYER ME1 ;
  RECT 488.755 0.000 489.075 0.600 ;
 END
 ANTENNAPARTIALMETALAREA                  1.058 LAYER ME2 ;
 ANTENNAGATEAREA                          0.072 LAYER ME2 ;
 ANTENNAGATEAREA                          0.072 LAYER ME3 ;
 ANTENNAGATEAREA                          0.072 LAYER ME4 ;
 ANTENNADIFFAREA                          0.160 LAYER ME2 ;
 ANTENNADIFFAREA                          0.160 LAYER ME3 ;
 ANTENNADIFFAREA                          0.160 LAYER ME4 ;
 ANTENNAMAXAREACAR                       21.782 LAYER ME2 ;
 ANTENNAMAXAREACAR                       24.449 LAYER ME3 ;
 ANTENNAMAXAREACAR                       27.116 LAYER ME4 ;
END DI111
PIN DO111
  DIRECTION OUTPUT ;
 PORT
  LAYER ME4 ;
  RECT 488.193 0.000 488.513 0.600 ;
  LAYER ME3 ;
  RECT 488.193 0.000 488.513 0.600 ;
  LAYER ME2 ;
  RECT 488.193 0.000 488.513 0.600 ;
  LAYER ME1 ;
  RECT 488.193 0.000 488.513 0.600 ;
 END
 ANTENNAPARTIALMETALAREA                  5.273 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME3 ;
 ANTENNADIFFAREA                          1.293 LAYER ME4 ;
END DO111
PIN DI110
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 484.751 0.000 485.071 0.600 ;
  LAYER ME3 ;
  RECT 484.751 0.000 485.071 0.600 ;
  LAYER ME2 ;
  RECT 484.751 0.000 485.071 0.600 ;
  LAYER ME1 ;
  RECT 484.751 0.000 485.071 0.600 ;
 END
 ANTENNAPARTIALMETALAREA                  1.058 LAYER ME2 ;
 ANTENNAGATEAREA                          0.072 LAYER ME2 ;
 ANTENNAGATEAREA                          0.072 LAYER ME3 ;
 ANTENNAGATEAREA                          0.072 LAYER ME4 ;
 ANTENNADIFFAREA                          0.160 LAYER ME2 ;
 ANTENNADIFFAREA                          0.160 LAYER ME3 ;
 ANTENNADIFFAREA                          0.160 LAYER ME4 ;
 ANTENNAMAXAREACAR                       21.782 LAYER ME2 ;
 ANTENNAMAXAREACAR                       24.449 LAYER ME3 ;
 ANTENNAMAXAREACAR                       27.116 LAYER ME4 ;
END DI110
PIN DO110
  DIRECTION OUTPUT ;
 PORT
  LAYER ME4 ;
  RECT 484.189 0.000 484.509 0.600 ;
  LAYER ME3 ;
  RECT 484.189 0.000 484.509 0.600 ;
  LAYER ME2 ;
  RECT 484.189 0.000 484.509 0.600 ;
  LAYER ME1 ;
  RECT 484.189 0.000 484.509 0.600 ;
 END
 ANTENNAPARTIALMETALAREA                  5.273 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME3 ;
 ANTENNADIFFAREA                          1.293 LAYER ME4 ;
END DO110
PIN DI109
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 480.747 0.000 481.067 0.600 ;
  LAYER ME3 ;
  RECT 480.747 0.000 481.067 0.600 ;
  LAYER ME2 ;
  RECT 480.747 0.000 481.067 0.600 ;
  LAYER ME1 ;
  RECT 480.747 0.000 481.067 0.600 ;
 END
 ANTENNAPARTIALMETALAREA                  1.058 LAYER ME2 ;
 ANTENNAGATEAREA                          0.072 LAYER ME2 ;
 ANTENNAGATEAREA                          0.072 LAYER ME3 ;
 ANTENNAGATEAREA                          0.072 LAYER ME4 ;
 ANTENNADIFFAREA                          0.160 LAYER ME2 ;
 ANTENNADIFFAREA                          0.160 LAYER ME3 ;
 ANTENNADIFFAREA                          0.160 LAYER ME4 ;
 ANTENNAMAXAREACAR                       21.782 LAYER ME2 ;
 ANTENNAMAXAREACAR                       24.449 LAYER ME3 ;
 ANTENNAMAXAREACAR                       27.116 LAYER ME4 ;
END DI109
PIN DO109
  DIRECTION OUTPUT ;
 PORT
  LAYER ME4 ;
  RECT 480.185 0.000 480.505 0.600 ;
  LAYER ME3 ;
  RECT 480.185 0.000 480.505 0.600 ;
  LAYER ME2 ;
  RECT 480.185 0.000 480.505 0.600 ;
  LAYER ME1 ;
  RECT 480.185 0.000 480.505 0.600 ;
 END
 ANTENNAPARTIALMETALAREA                  5.273 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME3 ;
 ANTENNADIFFAREA                          1.293 LAYER ME4 ;
END DO109
PIN DI108
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 476.743 0.000 477.063 0.600 ;
  LAYER ME3 ;
  RECT 476.743 0.000 477.063 0.600 ;
  LAYER ME2 ;
  RECT 476.743 0.000 477.063 0.600 ;
  LAYER ME1 ;
  RECT 476.743 0.000 477.063 0.600 ;
 END
 ANTENNAPARTIALMETALAREA                  1.058 LAYER ME2 ;
 ANTENNAGATEAREA                          0.072 LAYER ME2 ;
 ANTENNAGATEAREA                          0.072 LAYER ME3 ;
 ANTENNAGATEAREA                          0.072 LAYER ME4 ;
 ANTENNADIFFAREA                          0.160 LAYER ME2 ;
 ANTENNADIFFAREA                          0.160 LAYER ME3 ;
 ANTENNADIFFAREA                          0.160 LAYER ME4 ;
 ANTENNAMAXAREACAR                       21.782 LAYER ME2 ;
 ANTENNAMAXAREACAR                       24.449 LAYER ME3 ;
 ANTENNAMAXAREACAR                       27.116 LAYER ME4 ;
END DI108
PIN DO108
  DIRECTION OUTPUT ;
 PORT
  LAYER ME4 ;
  RECT 476.181 0.000 476.501 0.600 ;
  LAYER ME3 ;
  RECT 476.181 0.000 476.501 0.600 ;
  LAYER ME2 ;
  RECT 476.181 0.000 476.501 0.600 ;
  LAYER ME1 ;
  RECT 476.181 0.000 476.501 0.600 ;
 END
 ANTENNAPARTIALMETALAREA                  5.273 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME3 ;
 ANTENNADIFFAREA                          1.293 LAYER ME4 ;
END DO108
PIN DI107
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 472.739 0.000 473.059 0.600 ;
  LAYER ME3 ;
  RECT 472.739 0.000 473.059 0.600 ;
  LAYER ME2 ;
  RECT 472.739 0.000 473.059 0.600 ;
  LAYER ME1 ;
  RECT 472.739 0.000 473.059 0.600 ;
 END
 ANTENNAPARTIALMETALAREA                  1.058 LAYER ME2 ;
 ANTENNAGATEAREA                          0.072 LAYER ME2 ;
 ANTENNAGATEAREA                          0.072 LAYER ME3 ;
 ANTENNAGATEAREA                          0.072 LAYER ME4 ;
 ANTENNADIFFAREA                          0.160 LAYER ME2 ;
 ANTENNADIFFAREA                          0.160 LAYER ME3 ;
 ANTENNADIFFAREA                          0.160 LAYER ME4 ;
 ANTENNAMAXAREACAR                       21.782 LAYER ME2 ;
 ANTENNAMAXAREACAR                       24.449 LAYER ME3 ;
 ANTENNAMAXAREACAR                       27.116 LAYER ME4 ;
END DI107
PIN DO107
  DIRECTION OUTPUT ;
 PORT
  LAYER ME4 ;
  RECT 472.177 0.000 472.497 0.600 ;
  LAYER ME3 ;
  RECT 472.177 0.000 472.497 0.600 ;
  LAYER ME2 ;
  RECT 472.177 0.000 472.497 0.600 ;
  LAYER ME1 ;
  RECT 472.177 0.000 472.497 0.600 ;
 END
 ANTENNAPARTIALMETALAREA                  5.273 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME3 ;
 ANTENNADIFFAREA                          1.293 LAYER ME4 ;
END DO107
PIN DI106
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 468.735 0.000 469.055 0.600 ;
  LAYER ME3 ;
  RECT 468.735 0.000 469.055 0.600 ;
  LAYER ME2 ;
  RECT 468.735 0.000 469.055 0.600 ;
  LAYER ME1 ;
  RECT 468.735 0.000 469.055 0.600 ;
 END
 ANTENNAPARTIALMETALAREA                  1.058 LAYER ME2 ;
 ANTENNAGATEAREA                          0.072 LAYER ME2 ;
 ANTENNAGATEAREA                          0.072 LAYER ME3 ;
 ANTENNAGATEAREA                          0.072 LAYER ME4 ;
 ANTENNADIFFAREA                          0.160 LAYER ME2 ;
 ANTENNADIFFAREA                          0.160 LAYER ME3 ;
 ANTENNADIFFAREA                          0.160 LAYER ME4 ;
 ANTENNAMAXAREACAR                       21.782 LAYER ME2 ;
 ANTENNAMAXAREACAR                       24.449 LAYER ME3 ;
 ANTENNAMAXAREACAR                       27.116 LAYER ME4 ;
END DI106
PIN DO106
  DIRECTION OUTPUT ;
 PORT
  LAYER ME4 ;
  RECT 468.173 0.000 468.493 0.600 ;
  LAYER ME3 ;
  RECT 468.173 0.000 468.493 0.600 ;
  LAYER ME2 ;
  RECT 468.173 0.000 468.493 0.600 ;
  LAYER ME1 ;
  RECT 468.173 0.000 468.493 0.600 ;
 END
 ANTENNAPARTIALMETALAREA                  5.273 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME3 ;
 ANTENNADIFFAREA                          1.293 LAYER ME4 ;
END DO106
PIN DI105
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 464.731 0.000 465.051 0.600 ;
  LAYER ME3 ;
  RECT 464.731 0.000 465.051 0.600 ;
  LAYER ME2 ;
  RECT 464.731 0.000 465.051 0.600 ;
  LAYER ME1 ;
  RECT 464.731 0.000 465.051 0.600 ;
 END
 ANTENNAPARTIALMETALAREA                  1.058 LAYER ME2 ;
 ANTENNAGATEAREA                          0.072 LAYER ME2 ;
 ANTENNAGATEAREA                          0.072 LAYER ME3 ;
 ANTENNAGATEAREA                          0.072 LAYER ME4 ;
 ANTENNADIFFAREA                          0.160 LAYER ME2 ;
 ANTENNADIFFAREA                          0.160 LAYER ME3 ;
 ANTENNADIFFAREA                          0.160 LAYER ME4 ;
 ANTENNAMAXAREACAR                       21.782 LAYER ME2 ;
 ANTENNAMAXAREACAR                       24.449 LAYER ME3 ;
 ANTENNAMAXAREACAR                       27.116 LAYER ME4 ;
END DI105
PIN DO105
  DIRECTION OUTPUT ;
 PORT
  LAYER ME4 ;
  RECT 464.169 0.000 464.489 0.600 ;
  LAYER ME3 ;
  RECT 464.169 0.000 464.489 0.600 ;
  LAYER ME2 ;
  RECT 464.169 0.000 464.489 0.600 ;
  LAYER ME1 ;
  RECT 464.169 0.000 464.489 0.600 ;
 END
 ANTENNAPARTIALMETALAREA                  5.273 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME3 ;
 ANTENNADIFFAREA                          1.293 LAYER ME4 ;
END DO105
PIN DI104
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 460.727 0.000 461.047 0.600 ;
  LAYER ME3 ;
  RECT 460.727 0.000 461.047 0.600 ;
  LAYER ME2 ;
  RECT 460.727 0.000 461.047 0.600 ;
  LAYER ME1 ;
  RECT 460.727 0.000 461.047 0.600 ;
 END
 ANTENNAPARTIALMETALAREA                  1.058 LAYER ME2 ;
 ANTENNAGATEAREA                          0.072 LAYER ME2 ;
 ANTENNAGATEAREA                          0.072 LAYER ME3 ;
 ANTENNAGATEAREA                          0.072 LAYER ME4 ;
 ANTENNADIFFAREA                          0.160 LAYER ME2 ;
 ANTENNADIFFAREA                          0.160 LAYER ME3 ;
 ANTENNADIFFAREA                          0.160 LAYER ME4 ;
 ANTENNAMAXAREACAR                       21.782 LAYER ME2 ;
 ANTENNAMAXAREACAR                       24.449 LAYER ME3 ;
 ANTENNAMAXAREACAR                       27.116 LAYER ME4 ;
END DI104
PIN DO104
  DIRECTION OUTPUT ;
 PORT
  LAYER ME4 ;
  RECT 460.165 0.000 460.485 0.600 ;
  LAYER ME3 ;
  RECT 460.165 0.000 460.485 0.600 ;
  LAYER ME2 ;
  RECT 460.165 0.000 460.485 0.600 ;
  LAYER ME1 ;
  RECT 460.165 0.000 460.485 0.600 ;
 END
 ANTENNAPARTIALMETALAREA                  5.273 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME3 ;
 ANTENNADIFFAREA                          1.293 LAYER ME4 ;
END DO104
PIN DI103
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 456.723 0.000 457.043 0.600 ;
  LAYER ME3 ;
  RECT 456.723 0.000 457.043 0.600 ;
  LAYER ME2 ;
  RECT 456.723 0.000 457.043 0.600 ;
  LAYER ME1 ;
  RECT 456.723 0.000 457.043 0.600 ;
 END
 ANTENNAPARTIALMETALAREA                  1.058 LAYER ME2 ;
 ANTENNAGATEAREA                          0.072 LAYER ME2 ;
 ANTENNAGATEAREA                          0.072 LAYER ME3 ;
 ANTENNAGATEAREA                          0.072 LAYER ME4 ;
 ANTENNADIFFAREA                          0.160 LAYER ME2 ;
 ANTENNADIFFAREA                          0.160 LAYER ME3 ;
 ANTENNADIFFAREA                          0.160 LAYER ME4 ;
 ANTENNAMAXAREACAR                       21.782 LAYER ME2 ;
 ANTENNAMAXAREACAR                       24.449 LAYER ME3 ;
 ANTENNAMAXAREACAR                       27.116 LAYER ME4 ;
END DI103
PIN DO103
  DIRECTION OUTPUT ;
 PORT
  LAYER ME4 ;
  RECT 456.161 0.000 456.481 0.600 ;
  LAYER ME3 ;
  RECT 456.161 0.000 456.481 0.600 ;
  LAYER ME2 ;
  RECT 456.161 0.000 456.481 0.600 ;
  LAYER ME1 ;
  RECT 456.161 0.000 456.481 0.600 ;
 END
 ANTENNAPARTIALMETALAREA                  5.273 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME3 ;
 ANTENNADIFFAREA                          1.293 LAYER ME4 ;
END DO103
PIN DI102
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 452.719 0.000 453.039 0.600 ;
  LAYER ME3 ;
  RECT 452.719 0.000 453.039 0.600 ;
  LAYER ME2 ;
  RECT 452.719 0.000 453.039 0.600 ;
  LAYER ME1 ;
  RECT 452.719 0.000 453.039 0.600 ;
 END
 ANTENNAPARTIALMETALAREA                  1.058 LAYER ME2 ;
 ANTENNAGATEAREA                          0.072 LAYER ME2 ;
 ANTENNAGATEAREA                          0.072 LAYER ME3 ;
 ANTENNAGATEAREA                          0.072 LAYER ME4 ;
 ANTENNADIFFAREA                          0.160 LAYER ME2 ;
 ANTENNADIFFAREA                          0.160 LAYER ME3 ;
 ANTENNADIFFAREA                          0.160 LAYER ME4 ;
 ANTENNAMAXAREACAR                       21.782 LAYER ME2 ;
 ANTENNAMAXAREACAR                       24.449 LAYER ME3 ;
 ANTENNAMAXAREACAR                       27.116 LAYER ME4 ;
END DI102
PIN DO102
  DIRECTION OUTPUT ;
 PORT
  LAYER ME4 ;
  RECT 452.157 0.000 452.477 0.600 ;
  LAYER ME3 ;
  RECT 452.157 0.000 452.477 0.600 ;
  LAYER ME2 ;
  RECT 452.157 0.000 452.477 0.600 ;
  LAYER ME1 ;
  RECT 452.157 0.000 452.477 0.600 ;
 END
 ANTENNAPARTIALMETALAREA                  5.273 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME3 ;
 ANTENNADIFFAREA                          1.293 LAYER ME4 ;
END DO102
PIN DI101
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 448.715 0.000 449.035 0.600 ;
  LAYER ME3 ;
  RECT 448.715 0.000 449.035 0.600 ;
  LAYER ME2 ;
  RECT 448.715 0.000 449.035 0.600 ;
  LAYER ME1 ;
  RECT 448.715 0.000 449.035 0.600 ;
 END
 ANTENNAPARTIALMETALAREA                  1.058 LAYER ME2 ;
 ANTENNAGATEAREA                          0.072 LAYER ME2 ;
 ANTENNAGATEAREA                          0.072 LAYER ME3 ;
 ANTENNAGATEAREA                          0.072 LAYER ME4 ;
 ANTENNADIFFAREA                          0.160 LAYER ME2 ;
 ANTENNADIFFAREA                          0.160 LAYER ME3 ;
 ANTENNADIFFAREA                          0.160 LAYER ME4 ;
 ANTENNAMAXAREACAR                       21.782 LAYER ME2 ;
 ANTENNAMAXAREACAR                       24.449 LAYER ME3 ;
 ANTENNAMAXAREACAR                       27.116 LAYER ME4 ;
END DI101
PIN DO101
  DIRECTION OUTPUT ;
 PORT
  LAYER ME4 ;
  RECT 448.153 0.000 448.473 0.600 ;
  LAYER ME3 ;
  RECT 448.153 0.000 448.473 0.600 ;
  LAYER ME2 ;
  RECT 448.153 0.000 448.473 0.600 ;
  LAYER ME1 ;
  RECT 448.153 0.000 448.473 0.600 ;
 END
 ANTENNAPARTIALMETALAREA                  5.273 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME3 ;
 ANTENNADIFFAREA                          1.293 LAYER ME4 ;
END DO101
PIN DI100
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 444.711 0.000 445.031 0.600 ;
  LAYER ME3 ;
  RECT 444.711 0.000 445.031 0.600 ;
  LAYER ME2 ;
  RECT 444.711 0.000 445.031 0.600 ;
  LAYER ME1 ;
  RECT 444.711 0.000 445.031 0.600 ;
 END
 ANTENNAPARTIALMETALAREA                  1.058 LAYER ME2 ;
 ANTENNAGATEAREA                          0.072 LAYER ME2 ;
 ANTENNAGATEAREA                          0.072 LAYER ME3 ;
 ANTENNAGATEAREA                          0.072 LAYER ME4 ;
 ANTENNADIFFAREA                          0.160 LAYER ME2 ;
 ANTENNADIFFAREA                          0.160 LAYER ME3 ;
 ANTENNADIFFAREA                          0.160 LAYER ME4 ;
 ANTENNAMAXAREACAR                       21.782 LAYER ME2 ;
 ANTENNAMAXAREACAR                       24.449 LAYER ME3 ;
 ANTENNAMAXAREACAR                       27.116 LAYER ME4 ;
END DI100
PIN DO100
  DIRECTION OUTPUT ;
 PORT
  LAYER ME4 ;
  RECT 444.149 0.000 444.469 0.600 ;
  LAYER ME3 ;
  RECT 444.149 0.000 444.469 0.600 ;
  LAYER ME2 ;
  RECT 444.149 0.000 444.469 0.600 ;
  LAYER ME1 ;
  RECT 444.149 0.000 444.469 0.600 ;
 END
 ANTENNAPARTIALMETALAREA                  5.273 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME3 ;
 ANTENNADIFFAREA                          1.293 LAYER ME4 ;
END DO100
PIN DI99
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 440.707 0.000 441.027 0.600 ;
  LAYER ME3 ;
  RECT 440.707 0.000 441.027 0.600 ;
  LAYER ME2 ;
  RECT 440.707 0.000 441.027 0.600 ;
  LAYER ME1 ;
  RECT 440.707 0.000 441.027 0.600 ;
 END
 ANTENNAPARTIALMETALAREA                  1.058 LAYER ME2 ;
 ANTENNAGATEAREA                          0.072 LAYER ME2 ;
 ANTENNAGATEAREA                          0.072 LAYER ME3 ;
 ANTENNAGATEAREA                          0.072 LAYER ME4 ;
 ANTENNADIFFAREA                          0.160 LAYER ME2 ;
 ANTENNADIFFAREA                          0.160 LAYER ME3 ;
 ANTENNADIFFAREA                          0.160 LAYER ME4 ;
 ANTENNAMAXAREACAR                       21.782 LAYER ME2 ;
 ANTENNAMAXAREACAR                       24.449 LAYER ME3 ;
 ANTENNAMAXAREACAR                       27.116 LAYER ME4 ;
END DI99
PIN DO99
  DIRECTION OUTPUT ;
 PORT
  LAYER ME4 ;
  RECT 440.145 0.000 440.465 0.600 ;
  LAYER ME3 ;
  RECT 440.145 0.000 440.465 0.600 ;
  LAYER ME2 ;
  RECT 440.145 0.000 440.465 0.600 ;
  LAYER ME1 ;
  RECT 440.145 0.000 440.465 0.600 ;
 END
 ANTENNAPARTIALMETALAREA                  5.273 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME3 ;
 ANTENNADIFFAREA                          1.293 LAYER ME4 ;
END DO99
PIN DI98
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 436.703 0.000 437.023 0.600 ;
  LAYER ME3 ;
  RECT 436.703 0.000 437.023 0.600 ;
  LAYER ME2 ;
  RECT 436.703 0.000 437.023 0.600 ;
  LAYER ME1 ;
  RECT 436.703 0.000 437.023 0.600 ;
 END
 ANTENNAPARTIALMETALAREA                  1.058 LAYER ME2 ;
 ANTENNAGATEAREA                          0.072 LAYER ME2 ;
 ANTENNAGATEAREA                          0.072 LAYER ME3 ;
 ANTENNAGATEAREA                          0.072 LAYER ME4 ;
 ANTENNADIFFAREA                          0.160 LAYER ME2 ;
 ANTENNADIFFAREA                          0.160 LAYER ME3 ;
 ANTENNADIFFAREA                          0.160 LAYER ME4 ;
 ANTENNAMAXAREACAR                       21.782 LAYER ME2 ;
 ANTENNAMAXAREACAR                       24.449 LAYER ME3 ;
 ANTENNAMAXAREACAR                       27.116 LAYER ME4 ;
END DI98
PIN DO98
  DIRECTION OUTPUT ;
 PORT
  LAYER ME4 ;
  RECT 436.141 0.000 436.461 0.600 ;
  LAYER ME3 ;
  RECT 436.141 0.000 436.461 0.600 ;
  LAYER ME2 ;
  RECT 436.141 0.000 436.461 0.600 ;
  LAYER ME1 ;
  RECT 436.141 0.000 436.461 0.600 ;
 END
 ANTENNAPARTIALMETALAREA                  5.273 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME3 ;
 ANTENNADIFFAREA                          1.293 LAYER ME4 ;
END DO98
PIN DI97
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 432.699 0.000 433.019 0.600 ;
  LAYER ME3 ;
  RECT 432.699 0.000 433.019 0.600 ;
  LAYER ME2 ;
  RECT 432.699 0.000 433.019 0.600 ;
  LAYER ME1 ;
  RECT 432.699 0.000 433.019 0.600 ;
 END
 ANTENNAPARTIALMETALAREA                  1.058 LAYER ME2 ;
 ANTENNAGATEAREA                          0.072 LAYER ME2 ;
 ANTENNAGATEAREA                          0.072 LAYER ME3 ;
 ANTENNAGATEAREA                          0.072 LAYER ME4 ;
 ANTENNADIFFAREA                          0.160 LAYER ME2 ;
 ANTENNADIFFAREA                          0.160 LAYER ME3 ;
 ANTENNADIFFAREA                          0.160 LAYER ME4 ;
 ANTENNAMAXAREACAR                       21.782 LAYER ME2 ;
 ANTENNAMAXAREACAR                       24.449 LAYER ME3 ;
 ANTENNAMAXAREACAR                       27.116 LAYER ME4 ;
END DI97
PIN DO97
  DIRECTION OUTPUT ;
 PORT
  LAYER ME4 ;
  RECT 432.137 0.000 432.457 0.600 ;
  LAYER ME3 ;
  RECT 432.137 0.000 432.457 0.600 ;
  LAYER ME2 ;
  RECT 432.137 0.000 432.457 0.600 ;
  LAYER ME1 ;
  RECT 432.137 0.000 432.457 0.600 ;
 END
 ANTENNAPARTIALMETALAREA                  5.273 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME3 ;
 ANTENNADIFFAREA                          1.293 LAYER ME4 ;
END DO97
PIN DI96
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 428.133 0.000 428.453 0.600 ;
  LAYER ME3 ;
  RECT 428.133 0.000 428.453 0.600 ;
  LAYER ME2 ;
  RECT 428.133 0.000 428.453 0.600 ;
  LAYER ME1 ;
  RECT 428.133 0.000 428.453 0.600 ;
 END
 ANTENNAPARTIALMETALAREA                  0.346 LAYER ME1 ;
 ANTENNAPARTIALMETALAREA                  1.466 LAYER ME2 ;
 ANTENNAPARTIALMETALAREA                  0.508 LAYER ME3 ;
 ANTENNAGATEAREA                          0.072 LAYER ME3 ;
 ANTENNAGATEAREA                          0.072 LAYER ME4 ;
 ANTENNADIFFAREA                          0.218 LAYER ME1 ;
 ANTENNADIFFAREA                          0.218 LAYER ME2 ;
 ANTENNADIFFAREA                          0.218 LAYER ME3 ;
 ANTENNADIFFAREA                          0.218 LAYER ME4 ;
 ANTENNAMAXAREACAR                       17.267 LAYER ME3 ;
 ANTENNAMAXAREACAR                       19.933 LAYER ME4 ;
END DI96
PIN DO96
  DIRECTION OUTPUT ;
 PORT
  LAYER ME4 ;
  RECT 428.695 0.000 429.015 0.600 ;
  LAYER ME3 ;
  RECT 428.695 0.000 429.015 0.600 ;
  LAYER ME2 ;
  RECT 428.695 0.000 429.015 0.600 ;
  LAYER ME1 ;
  RECT 428.695 0.000 429.015 0.600 ;
 END
 ANTENNAPARTIALMETALAREA                  5.602 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME3 ;
 ANTENNADIFFAREA                          1.293 LAYER ME4 ;
END DO96
PIN WEB6
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 426.693 0.000 427.013 0.600 ;
  LAYER ME3 ;
  RECT 426.693 0.000 427.013 0.600 ;
  LAYER ME2 ;
  RECT 426.693 0.000 427.013 0.600 ;
  LAYER ME1 ;
  RECT 426.693 0.000 427.013 0.600 ;
 END
 ANTENNAPARTIALMETALAREA                  1.036 LAYER ME2 ;
 ANTENNAGATEAREA                          0.288 LAYER ME2 ;
 ANTENNAGATEAREA                          0.288 LAYER ME3 ;
 ANTENNAGATEAREA                          0.288 LAYER ME4 ;
 ANTENNADIFFAREA                          0.206 LAYER ME2 ;
 ANTENNADIFFAREA                          0.206 LAYER ME3 ;
 ANTENNADIFFAREA                          0.206 LAYER ME4 ;
 ANTENNAMAXAREACAR                        5.844 LAYER ME2 ;
 ANTENNAMAXAREACAR                        6.511 LAYER ME3 ;
 ANTENNAMAXAREACAR                        7.178 LAYER ME4 ;
END WEB6
PIN DI95
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 424.691 0.000 425.011 0.600 ;
  LAYER ME3 ;
  RECT 424.691 0.000 425.011 0.600 ;
  LAYER ME2 ;
  RECT 424.691 0.000 425.011 0.600 ;
  LAYER ME1 ;
  RECT 424.691 0.000 425.011 0.600 ;
 END
 ANTENNAPARTIALMETALAREA                  1.058 LAYER ME2 ;
 ANTENNAGATEAREA                          0.072 LAYER ME2 ;
 ANTENNAGATEAREA                          0.072 LAYER ME3 ;
 ANTENNAGATEAREA                          0.072 LAYER ME4 ;
 ANTENNADIFFAREA                          0.160 LAYER ME2 ;
 ANTENNADIFFAREA                          0.160 LAYER ME3 ;
 ANTENNADIFFAREA                          0.160 LAYER ME4 ;
 ANTENNAMAXAREACAR                       21.782 LAYER ME2 ;
 ANTENNAMAXAREACAR                       24.449 LAYER ME3 ;
 ANTENNAMAXAREACAR                       27.116 LAYER ME4 ;
END DI95
PIN DO95
  DIRECTION OUTPUT ;
 PORT
  LAYER ME4 ;
  RECT 424.129 0.000 424.449 0.600 ;
  LAYER ME3 ;
  RECT 424.129 0.000 424.449 0.600 ;
  LAYER ME2 ;
  RECT 424.129 0.000 424.449 0.600 ;
  LAYER ME1 ;
  RECT 424.129 0.000 424.449 0.600 ;
 END
 ANTENNAPARTIALMETALAREA                  5.273 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME3 ;
 ANTENNADIFFAREA                          1.293 LAYER ME4 ;
END DO95
PIN DI94
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 420.687 0.000 421.007 0.600 ;
  LAYER ME3 ;
  RECT 420.687 0.000 421.007 0.600 ;
  LAYER ME2 ;
  RECT 420.687 0.000 421.007 0.600 ;
  LAYER ME1 ;
  RECT 420.687 0.000 421.007 0.600 ;
 END
 ANTENNAPARTIALMETALAREA                  1.058 LAYER ME2 ;
 ANTENNAGATEAREA                          0.072 LAYER ME2 ;
 ANTENNAGATEAREA                          0.072 LAYER ME3 ;
 ANTENNAGATEAREA                          0.072 LAYER ME4 ;
 ANTENNADIFFAREA                          0.160 LAYER ME2 ;
 ANTENNADIFFAREA                          0.160 LAYER ME3 ;
 ANTENNADIFFAREA                          0.160 LAYER ME4 ;
 ANTENNAMAXAREACAR                       21.782 LAYER ME2 ;
 ANTENNAMAXAREACAR                       24.449 LAYER ME3 ;
 ANTENNAMAXAREACAR                       27.116 LAYER ME4 ;
END DI94
PIN DO94
  DIRECTION OUTPUT ;
 PORT
  LAYER ME4 ;
  RECT 420.125 0.000 420.445 0.600 ;
  LAYER ME3 ;
  RECT 420.125 0.000 420.445 0.600 ;
  LAYER ME2 ;
  RECT 420.125 0.000 420.445 0.600 ;
  LAYER ME1 ;
  RECT 420.125 0.000 420.445 0.600 ;
 END
 ANTENNAPARTIALMETALAREA                  5.273 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME3 ;
 ANTENNADIFFAREA                          1.293 LAYER ME4 ;
END DO94
PIN DI93
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 416.683 0.000 417.003 0.600 ;
  LAYER ME3 ;
  RECT 416.683 0.000 417.003 0.600 ;
  LAYER ME2 ;
  RECT 416.683 0.000 417.003 0.600 ;
  LAYER ME1 ;
  RECT 416.683 0.000 417.003 0.600 ;
 END
 ANTENNAPARTIALMETALAREA                  1.058 LAYER ME2 ;
 ANTENNAGATEAREA                          0.072 LAYER ME2 ;
 ANTENNAGATEAREA                          0.072 LAYER ME3 ;
 ANTENNAGATEAREA                          0.072 LAYER ME4 ;
 ANTENNADIFFAREA                          0.160 LAYER ME2 ;
 ANTENNADIFFAREA                          0.160 LAYER ME3 ;
 ANTENNADIFFAREA                          0.160 LAYER ME4 ;
 ANTENNAMAXAREACAR                       21.782 LAYER ME2 ;
 ANTENNAMAXAREACAR                       24.449 LAYER ME3 ;
 ANTENNAMAXAREACAR                       27.116 LAYER ME4 ;
END DI93
PIN DO93
  DIRECTION OUTPUT ;
 PORT
  LAYER ME4 ;
  RECT 416.121 0.000 416.441 0.600 ;
  LAYER ME3 ;
  RECT 416.121 0.000 416.441 0.600 ;
  LAYER ME2 ;
  RECT 416.121 0.000 416.441 0.600 ;
  LAYER ME1 ;
  RECT 416.121 0.000 416.441 0.600 ;
 END
 ANTENNAPARTIALMETALAREA                  5.273 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME3 ;
 ANTENNADIFFAREA                          1.293 LAYER ME4 ;
END DO93
PIN DI92
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 412.679 0.000 412.999 0.600 ;
  LAYER ME3 ;
  RECT 412.679 0.000 412.999 0.600 ;
  LAYER ME2 ;
  RECT 412.679 0.000 412.999 0.600 ;
  LAYER ME1 ;
  RECT 412.679 0.000 412.999 0.600 ;
 END
 ANTENNAPARTIALMETALAREA                  1.058 LAYER ME2 ;
 ANTENNAGATEAREA                          0.072 LAYER ME2 ;
 ANTENNAGATEAREA                          0.072 LAYER ME3 ;
 ANTENNAGATEAREA                          0.072 LAYER ME4 ;
 ANTENNADIFFAREA                          0.160 LAYER ME2 ;
 ANTENNADIFFAREA                          0.160 LAYER ME3 ;
 ANTENNADIFFAREA                          0.160 LAYER ME4 ;
 ANTENNAMAXAREACAR                       21.782 LAYER ME2 ;
 ANTENNAMAXAREACAR                       24.449 LAYER ME3 ;
 ANTENNAMAXAREACAR                       27.116 LAYER ME4 ;
END DI92
PIN DO92
  DIRECTION OUTPUT ;
 PORT
  LAYER ME4 ;
  RECT 412.117 0.000 412.437 0.600 ;
  LAYER ME3 ;
  RECT 412.117 0.000 412.437 0.600 ;
  LAYER ME2 ;
  RECT 412.117 0.000 412.437 0.600 ;
  LAYER ME1 ;
  RECT 412.117 0.000 412.437 0.600 ;
 END
 ANTENNAPARTIALMETALAREA                  5.273 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME3 ;
 ANTENNADIFFAREA                          1.293 LAYER ME4 ;
END DO92
PIN DI91
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 408.675 0.000 408.995 0.600 ;
  LAYER ME3 ;
  RECT 408.675 0.000 408.995 0.600 ;
  LAYER ME2 ;
  RECT 408.675 0.000 408.995 0.600 ;
  LAYER ME1 ;
  RECT 408.675 0.000 408.995 0.600 ;
 END
 ANTENNAPARTIALMETALAREA                  1.058 LAYER ME2 ;
 ANTENNAGATEAREA                          0.072 LAYER ME2 ;
 ANTENNAGATEAREA                          0.072 LAYER ME3 ;
 ANTENNAGATEAREA                          0.072 LAYER ME4 ;
 ANTENNADIFFAREA                          0.160 LAYER ME2 ;
 ANTENNADIFFAREA                          0.160 LAYER ME3 ;
 ANTENNADIFFAREA                          0.160 LAYER ME4 ;
 ANTENNAMAXAREACAR                       21.782 LAYER ME2 ;
 ANTENNAMAXAREACAR                       24.449 LAYER ME3 ;
 ANTENNAMAXAREACAR                       27.116 LAYER ME4 ;
END DI91
PIN DO91
  DIRECTION OUTPUT ;
 PORT
  LAYER ME4 ;
  RECT 408.113 0.000 408.433 0.600 ;
  LAYER ME3 ;
  RECT 408.113 0.000 408.433 0.600 ;
  LAYER ME2 ;
  RECT 408.113 0.000 408.433 0.600 ;
  LAYER ME1 ;
  RECT 408.113 0.000 408.433 0.600 ;
 END
 ANTENNAPARTIALMETALAREA                  5.273 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME3 ;
 ANTENNADIFFAREA                          1.293 LAYER ME4 ;
END DO91
PIN DI90
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 404.671 0.000 404.991 0.600 ;
  LAYER ME3 ;
  RECT 404.671 0.000 404.991 0.600 ;
  LAYER ME2 ;
  RECT 404.671 0.000 404.991 0.600 ;
  LAYER ME1 ;
  RECT 404.671 0.000 404.991 0.600 ;
 END
 ANTENNAPARTIALMETALAREA                  1.058 LAYER ME2 ;
 ANTENNAGATEAREA                          0.072 LAYER ME2 ;
 ANTENNAGATEAREA                          0.072 LAYER ME3 ;
 ANTENNAGATEAREA                          0.072 LAYER ME4 ;
 ANTENNADIFFAREA                          0.160 LAYER ME2 ;
 ANTENNADIFFAREA                          0.160 LAYER ME3 ;
 ANTENNADIFFAREA                          0.160 LAYER ME4 ;
 ANTENNAMAXAREACAR                       21.782 LAYER ME2 ;
 ANTENNAMAXAREACAR                       24.449 LAYER ME3 ;
 ANTENNAMAXAREACAR                       27.116 LAYER ME4 ;
END DI90
PIN DO90
  DIRECTION OUTPUT ;
 PORT
  LAYER ME4 ;
  RECT 404.109 0.000 404.429 0.600 ;
  LAYER ME3 ;
  RECT 404.109 0.000 404.429 0.600 ;
  LAYER ME2 ;
  RECT 404.109 0.000 404.429 0.600 ;
  LAYER ME1 ;
  RECT 404.109 0.000 404.429 0.600 ;
 END
 ANTENNAPARTIALMETALAREA                  5.273 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME3 ;
 ANTENNADIFFAREA                          1.293 LAYER ME4 ;
END DO90
PIN DI89
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 400.667 0.000 400.987 0.600 ;
  LAYER ME3 ;
  RECT 400.667 0.000 400.987 0.600 ;
  LAYER ME2 ;
  RECT 400.667 0.000 400.987 0.600 ;
  LAYER ME1 ;
  RECT 400.667 0.000 400.987 0.600 ;
 END
 ANTENNAPARTIALMETALAREA                  1.058 LAYER ME2 ;
 ANTENNAGATEAREA                          0.072 LAYER ME2 ;
 ANTENNAGATEAREA                          0.072 LAYER ME3 ;
 ANTENNAGATEAREA                          0.072 LAYER ME4 ;
 ANTENNADIFFAREA                          0.160 LAYER ME2 ;
 ANTENNADIFFAREA                          0.160 LAYER ME3 ;
 ANTENNADIFFAREA                          0.160 LAYER ME4 ;
 ANTENNAMAXAREACAR                       21.782 LAYER ME2 ;
 ANTENNAMAXAREACAR                       24.449 LAYER ME3 ;
 ANTENNAMAXAREACAR                       27.116 LAYER ME4 ;
END DI89
PIN DO89
  DIRECTION OUTPUT ;
 PORT
  LAYER ME4 ;
  RECT 400.105 0.000 400.425 0.600 ;
  LAYER ME3 ;
  RECT 400.105 0.000 400.425 0.600 ;
  LAYER ME2 ;
  RECT 400.105 0.000 400.425 0.600 ;
  LAYER ME1 ;
  RECT 400.105 0.000 400.425 0.600 ;
 END
 ANTENNAPARTIALMETALAREA                  5.273 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME3 ;
 ANTENNADIFFAREA                          1.293 LAYER ME4 ;
END DO89
PIN DI88
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 396.663 0.000 396.983 0.600 ;
  LAYER ME3 ;
  RECT 396.663 0.000 396.983 0.600 ;
  LAYER ME2 ;
  RECT 396.663 0.000 396.983 0.600 ;
  LAYER ME1 ;
  RECT 396.663 0.000 396.983 0.600 ;
 END
 ANTENNAPARTIALMETALAREA                  1.058 LAYER ME2 ;
 ANTENNAGATEAREA                          0.072 LAYER ME2 ;
 ANTENNAGATEAREA                          0.072 LAYER ME3 ;
 ANTENNAGATEAREA                          0.072 LAYER ME4 ;
 ANTENNADIFFAREA                          0.160 LAYER ME2 ;
 ANTENNADIFFAREA                          0.160 LAYER ME3 ;
 ANTENNADIFFAREA                          0.160 LAYER ME4 ;
 ANTENNAMAXAREACAR                       21.782 LAYER ME2 ;
 ANTENNAMAXAREACAR                       24.449 LAYER ME3 ;
 ANTENNAMAXAREACAR                       27.116 LAYER ME4 ;
END DI88
PIN DO88
  DIRECTION OUTPUT ;
 PORT
  LAYER ME4 ;
  RECT 396.101 0.000 396.421 0.600 ;
  LAYER ME3 ;
  RECT 396.101 0.000 396.421 0.600 ;
  LAYER ME2 ;
  RECT 396.101 0.000 396.421 0.600 ;
  LAYER ME1 ;
  RECT 396.101 0.000 396.421 0.600 ;
 END
 ANTENNAPARTIALMETALAREA                  5.273 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME3 ;
 ANTENNADIFFAREA                          1.293 LAYER ME4 ;
END DO88
PIN DI87
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 392.659 0.000 392.979 0.600 ;
  LAYER ME3 ;
  RECT 392.659 0.000 392.979 0.600 ;
  LAYER ME2 ;
  RECT 392.659 0.000 392.979 0.600 ;
  LAYER ME1 ;
  RECT 392.659 0.000 392.979 0.600 ;
 END
 ANTENNAPARTIALMETALAREA                  1.058 LAYER ME2 ;
 ANTENNAGATEAREA                          0.072 LAYER ME2 ;
 ANTENNAGATEAREA                          0.072 LAYER ME3 ;
 ANTENNAGATEAREA                          0.072 LAYER ME4 ;
 ANTENNADIFFAREA                          0.160 LAYER ME2 ;
 ANTENNADIFFAREA                          0.160 LAYER ME3 ;
 ANTENNADIFFAREA                          0.160 LAYER ME4 ;
 ANTENNAMAXAREACAR                       21.782 LAYER ME2 ;
 ANTENNAMAXAREACAR                       24.449 LAYER ME3 ;
 ANTENNAMAXAREACAR                       27.116 LAYER ME4 ;
END DI87
PIN DO87
  DIRECTION OUTPUT ;
 PORT
  LAYER ME4 ;
  RECT 392.097 0.000 392.417 0.600 ;
  LAYER ME3 ;
  RECT 392.097 0.000 392.417 0.600 ;
  LAYER ME2 ;
  RECT 392.097 0.000 392.417 0.600 ;
  LAYER ME1 ;
  RECT 392.097 0.000 392.417 0.600 ;
 END
 ANTENNAPARTIALMETALAREA                  5.273 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME3 ;
 ANTENNADIFFAREA                          1.293 LAYER ME4 ;
END DO87
PIN DI86
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 388.655 0.000 388.975 0.600 ;
  LAYER ME3 ;
  RECT 388.655 0.000 388.975 0.600 ;
  LAYER ME2 ;
  RECT 388.655 0.000 388.975 0.600 ;
  LAYER ME1 ;
  RECT 388.655 0.000 388.975 0.600 ;
 END
 ANTENNAPARTIALMETALAREA                  1.058 LAYER ME2 ;
 ANTENNAGATEAREA                          0.072 LAYER ME2 ;
 ANTENNAGATEAREA                          0.072 LAYER ME3 ;
 ANTENNAGATEAREA                          0.072 LAYER ME4 ;
 ANTENNADIFFAREA                          0.160 LAYER ME2 ;
 ANTENNADIFFAREA                          0.160 LAYER ME3 ;
 ANTENNADIFFAREA                          0.160 LAYER ME4 ;
 ANTENNAMAXAREACAR                       21.782 LAYER ME2 ;
 ANTENNAMAXAREACAR                       24.449 LAYER ME3 ;
 ANTENNAMAXAREACAR                       27.116 LAYER ME4 ;
END DI86
PIN DO86
  DIRECTION OUTPUT ;
 PORT
  LAYER ME4 ;
  RECT 388.093 0.000 388.413 0.600 ;
  LAYER ME3 ;
  RECT 388.093 0.000 388.413 0.600 ;
  LAYER ME2 ;
  RECT 388.093 0.000 388.413 0.600 ;
  LAYER ME1 ;
  RECT 388.093 0.000 388.413 0.600 ;
 END
 ANTENNAPARTIALMETALAREA                  5.273 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME3 ;
 ANTENNADIFFAREA                          1.293 LAYER ME4 ;
END DO86
PIN DI85
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 384.651 0.000 384.971 0.600 ;
  LAYER ME3 ;
  RECT 384.651 0.000 384.971 0.600 ;
  LAYER ME2 ;
  RECT 384.651 0.000 384.971 0.600 ;
  LAYER ME1 ;
  RECT 384.651 0.000 384.971 0.600 ;
 END
 ANTENNAPARTIALMETALAREA                  1.058 LAYER ME2 ;
 ANTENNAGATEAREA                          0.072 LAYER ME2 ;
 ANTENNAGATEAREA                          0.072 LAYER ME3 ;
 ANTENNAGATEAREA                          0.072 LAYER ME4 ;
 ANTENNADIFFAREA                          0.160 LAYER ME2 ;
 ANTENNADIFFAREA                          0.160 LAYER ME3 ;
 ANTENNADIFFAREA                          0.160 LAYER ME4 ;
 ANTENNAMAXAREACAR                       21.782 LAYER ME2 ;
 ANTENNAMAXAREACAR                       24.449 LAYER ME3 ;
 ANTENNAMAXAREACAR                       27.116 LAYER ME4 ;
END DI85
PIN DO85
  DIRECTION OUTPUT ;
 PORT
  LAYER ME4 ;
  RECT 384.089 0.000 384.409 0.600 ;
  LAYER ME3 ;
  RECT 384.089 0.000 384.409 0.600 ;
  LAYER ME2 ;
  RECT 384.089 0.000 384.409 0.600 ;
  LAYER ME1 ;
  RECT 384.089 0.000 384.409 0.600 ;
 END
 ANTENNAPARTIALMETALAREA                  5.273 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME3 ;
 ANTENNADIFFAREA                          1.293 LAYER ME4 ;
END DO85
PIN DI84
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 380.647 0.000 380.967 0.600 ;
  LAYER ME3 ;
  RECT 380.647 0.000 380.967 0.600 ;
  LAYER ME2 ;
  RECT 380.647 0.000 380.967 0.600 ;
  LAYER ME1 ;
  RECT 380.647 0.000 380.967 0.600 ;
 END
 ANTENNAPARTIALMETALAREA                  1.058 LAYER ME2 ;
 ANTENNAGATEAREA                          0.072 LAYER ME2 ;
 ANTENNAGATEAREA                          0.072 LAYER ME3 ;
 ANTENNAGATEAREA                          0.072 LAYER ME4 ;
 ANTENNADIFFAREA                          0.160 LAYER ME2 ;
 ANTENNADIFFAREA                          0.160 LAYER ME3 ;
 ANTENNADIFFAREA                          0.160 LAYER ME4 ;
 ANTENNAMAXAREACAR                       21.782 LAYER ME2 ;
 ANTENNAMAXAREACAR                       24.449 LAYER ME3 ;
 ANTENNAMAXAREACAR                       27.116 LAYER ME4 ;
END DI84
PIN DO84
  DIRECTION OUTPUT ;
 PORT
  LAYER ME4 ;
  RECT 380.085 0.000 380.405 0.600 ;
  LAYER ME3 ;
  RECT 380.085 0.000 380.405 0.600 ;
  LAYER ME2 ;
  RECT 380.085 0.000 380.405 0.600 ;
  LAYER ME1 ;
  RECT 380.085 0.000 380.405 0.600 ;
 END
 ANTENNAPARTIALMETALAREA                  5.273 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME3 ;
 ANTENNADIFFAREA                          1.293 LAYER ME4 ;
END DO84
PIN DI83
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 376.643 0.000 376.963 0.600 ;
  LAYER ME3 ;
  RECT 376.643 0.000 376.963 0.600 ;
  LAYER ME2 ;
  RECT 376.643 0.000 376.963 0.600 ;
  LAYER ME1 ;
  RECT 376.643 0.000 376.963 0.600 ;
 END
 ANTENNAPARTIALMETALAREA                  1.058 LAYER ME2 ;
 ANTENNAGATEAREA                          0.072 LAYER ME2 ;
 ANTENNAGATEAREA                          0.072 LAYER ME3 ;
 ANTENNAGATEAREA                          0.072 LAYER ME4 ;
 ANTENNADIFFAREA                          0.160 LAYER ME2 ;
 ANTENNADIFFAREA                          0.160 LAYER ME3 ;
 ANTENNADIFFAREA                          0.160 LAYER ME4 ;
 ANTENNAMAXAREACAR                       21.782 LAYER ME2 ;
 ANTENNAMAXAREACAR                       24.449 LAYER ME3 ;
 ANTENNAMAXAREACAR                       27.116 LAYER ME4 ;
END DI83
PIN DO83
  DIRECTION OUTPUT ;
 PORT
  LAYER ME4 ;
  RECT 376.081 0.000 376.401 0.600 ;
  LAYER ME3 ;
  RECT 376.081 0.000 376.401 0.600 ;
  LAYER ME2 ;
  RECT 376.081 0.000 376.401 0.600 ;
  LAYER ME1 ;
  RECT 376.081 0.000 376.401 0.600 ;
 END
 ANTENNAPARTIALMETALAREA                  5.273 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME3 ;
 ANTENNADIFFAREA                          1.293 LAYER ME4 ;
END DO83
PIN DI82
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 372.639 0.000 372.959 0.600 ;
  LAYER ME3 ;
  RECT 372.639 0.000 372.959 0.600 ;
  LAYER ME2 ;
  RECT 372.639 0.000 372.959 0.600 ;
  LAYER ME1 ;
  RECT 372.639 0.000 372.959 0.600 ;
 END
 ANTENNAPARTIALMETALAREA                  1.058 LAYER ME2 ;
 ANTENNAGATEAREA                          0.072 LAYER ME2 ;
 ANTENNAGATEAREA                          0.072 LAYER ME3 ;
 ANTENNAGATEAREA                          0.072 LAYER ME4 ;
 ANTENNADIFFAREA                          0.160 LAYER ME2 ;
 ANTENNADIFFAREA                          0.160 LAYER ME3 ;
 ANTENNADIFFAREA                          0.160 LAYER ME4 ;
 ANTENNAMAXAREACAR                       21.782 LAYER ME2 ;
 ANTENNAMAXAREACAR                       24.449 LAYER ME3 ;
 ANTENNAMAXAREACAR                       27.116 LAYER ME4 ;
END DI82
PIN DO82
  DIRECTION OUTPUT ;
 PORT
  LAYER ME4 ;
  RECT 372.077 0.000 372.397 0.600 ;
  LAYER ME3 ;
  RECT 372.077 0.000 372.397 0.600 ;
  LAYER ME2 ;
  RECT 372.077 0.000 372.397 0.600 ;
  LAYER ME1 ;
  RECT 372.077 0.000 372.397 0.600 ;
 END
 ANTENNAPARTIALMETALAREA                  5.273 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME3 ;
 ANTENNADIFFAREA                          1.293 LAYER ME4 ;
END DO82
PIN DI81
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 368.635 0.000 368.955 0.600 ;
  LAYER ME3 ;
  RECT 368.635 0.000 368.955 0.600 ;
  LAYER ME2 ;
  RECT 368.635 0.000 368.955 0.600 ;
  LAYER ME1 ;
  RECT 368.635 0.000 368.955 0.600 ;
 END
 ANTENNAPARTIALMETALAREA                  1.058 LAYER ME2 ;
 ANTENNAGATEAREA                          0.072 LAYER ME2 ;
 ANTENNAGATEAREA                          0.072 LAYER ME3 ;
 ANTENNAGATEAREA                          0.072 LAYER ME4 ;
 ANTENNADIFFAREA                          0.160 LAYER ME2 ;
 ANTENNADIFFAREA                          0.160 LAYER ME3 ;
 ANTENNADIFFAREA                          0.160 LAYER ME4 ;
 ANTENNAMAXAREACAR                       21.782 LAYER ME2 ;
 ANTENNAMAXAREACAR                       24.449 LAYER ME3 ;
 ANTENNAMAXAREACAR                       27.116 LAYER ME4 ;
END DI81
PIN DO81
  DIRECTION OUTPUT ;
 PORT
  LAYER ME4 ;
  RECT 368.073 0.000 368.393 0.600 ;
  LAYER ME3 ;
  RECT 368.073 0.000 368.393 0.600 ;
  LAYER ME2 ;
  RECT 368.073 0.000 368.393 0.600 ;
  LAYER ME1 ;
  RECT 368.073 0.000 368.393 0.600 ;
 END
 ANTENNAPARTIALMETALAREA                  5.273 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME3 ;
 ANTENNADIFFAREA                          1.293 LAYER ME4 ;
END DO81
PIN DI80
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 364.069 0.000 364.389 0.600 ;
  LAYER ME3 ;
  RECT 364.069 0.000 364.389 0.600 ;
  LAYER ME2 ;
  RECT 364.069 0.000 364.389 0.600 ;
  LAYER ME1 ;
  RECT 364.069 0.000 364.389 0.600 ;
 END
 ANTENNAPARTIALMETALAREA                  0.346 LAYER ME1 ;
 ANTENNAPARTIALMETALAREA                  1.466 LAYER ME2 ;
 ANTENNAPARTIALMETALAREA                  0.508 LAYER ME3 ;
 ANTENNAGATEAREA                          0.072 LAYER ME3 ;
 ANTENNAGATEAREA                          0.072 LAYER ME4 ;
 ANTENNADIFFAREA                          0.218 LAYER ME1 ;
 ANTENNADIFFAREA                          0.218 LAYER ME2 ;
 ANTENNADIFFAREA                          0.218 LAYER ME3 ;
 ANTENNADIFFAREA                          0.218 LAYER ME4 ;
 ANTENNAMAXAREACAR                       17.267 LAYER ME3 ;
 ANTENNAMAXAREACAR                       19.933 LAYER ME4 ;
END DI80
PIN DO80
  DIRECTION OUTPUT ;
 PORT
  LAYER ME4 ;
  RECT 364.631 0.000 364.951 0.600 ;
  LAYER ME3 ;
  RECT 364.631 0.000 364.951 0.600 ;
  LAYER ME2 ;
  RECT 364.631 0.000 364.951 0.600 ;
  LAYER ME1 ;
  RECT 364.631 0.000 364.951 0.600 ;
 END
 ANTENNAPARTIALMETALAREA                  5.602 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME3 ;
 ANTENNADIFFAREA                          1.293 LAYER ME4 ;
END DO80
PIN WEB5
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 362.629 0.000 362.949 0.600 ;
  LAYER ME3 ;
  RECT 362.629 0.000 362.949 0.600 ;
  LAYER ME2 ;
  RECT 362.629 0.000 362.949 0.600 ;
  LAYER ME1 ;
  RECT 362.629 0.000 362.949 0.600 ;
 END
 ANTENNAPARTIALMETALAREA                  1.036 LAYER ME2 ;
 ANTENNAGATEAREA                          0.288 LAYER ME2 ;
 ANTENNAGATEAREA                          0.288 LAYER ME3 ;
 ANTENNAGATEAREA                          0.288 LAYER ME4 ;
 ANTENNADIFFAREA                          0.206 LAYER ME2 ;
 ANTENNADIFFAREA                          0.206 LAYER ME3 ;
 ANTENNADIFFAREA                          0.206 LAYER ME4 ;
 ANTENNAMAXAREACAR                        5.844 LAYER ME2 ;
 ANTENNAMAXAREACAR                        6.511 LAYER ME3 ;
 ANTENNAMAXAREACAR                        7.178 LAYER ME4 ;
END WEB5
PIN DI79
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 360.627 0.000 360.947 0.600 ;
  LAYER ME3 ;
  RECT 360.627 0.000 360.947 0.600 ;
  LAYER ME2 ;
  RECT 360.627 0.000 360.947 0.600 ;
  LAYER ME1 ;
  RECT 360.627 0.000 360.947 0.600 ;
 END
 ANTENNAPARTIALMETALAREA                  1.058 LAYER ME2 ;
 ANTENNAGATEAREA                          0.072 LAYER ME2 ;
 ANTENNAGATEAREA                          0.072 LAYER ME3 ;
 ANTENNAGATEAREA                          0.072 LAYER ME4 ;
 ANTENNADIFFAREA                          0.160 LAYER ME2 ;
 ANTENNADIFFAREA                          0.160 LAYER ME3 ;
 ANTENNADIFFAREA                          0.160 LAYER ME4 ;
 ANTENNAMAXAREACAR                       21.782 LAYER ME2 ;
 ANTENNAMAXAREACAR                       24.449 LAYER ME3 ;
 ANTENNAMAXAREACAR                       27.116 LAYER ME4 ;
END DI79
PIN DO79
  DIRECTION OUTPUT ;
 PORT
  LAYER ME4 ;
  RECT 360.065 0.000 360.385 0.600 ;
  LAYER ME3 ;
  RECT 360.065 0.000 360.385 0.600 ;
  LAYER ME2 ;
  RECT 360.065 0.000 360.385 0.600 ;
  LAYER ME1 ;
  RECT 360.065 0.000 360.385 0.600 ;
 END
 ANTENNAPARTIALMETALAREA                  5.273 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME3 ;
 ANTENNADIFFAREA                          1.293 LAYER ME4 ;
END DO79
PIN DI78
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 356.623 0.000 356.943 0.600 ;
  LAYER ME3 ;
  RECT 356.623 0.000 356.943 0.600 ;
  LAYER ME2 ;
  RECT 356.623 0.000 356.943 0.600 ;
  LAYER ME1 ;
  RECT 356.623 0.000 356.943 0.600 ;
 END
 ANTENNAPARTIALMETALAREA                  1.058 LAYER ME2 ;
 ANTENNAGATEAREA                          0.072 LAYER ME2 ;
 ANTENNAGATEAREA                          0.072 LAYER ME3 ;
 ANTENNAGATEAREA                          0.072 LAYER ME4 ;
 ANTENNADIFFAREA                          0.160 LAYER ME2 ;
 ANTENNADIFFAREA                          0.160 LAYER ME3 ;
 ANTENNADIFFAREA                          0.160 LAYER ME4 ;
 ANTENNAMAXAREACAR                       21.782 LAYER ME2 ;
 ANTENNAMAXAREACAR                       24.449 LAYER ME3 ;
 ANTENNAMAXAREACAR                       27.116 LAYER ME4 ;
END DI78
PIN DO78
  DIRECTION OUTPUT ;
 PORT
  LAYER ME4 ;
  RECT 356.061 0.000 356.381 0.600 ;
  LAYER ME3 ;
  RECT 356.061 0.000 356.381 0.600 ;
  LAYER ME2 ;
  RECT 356.061 0.000 356.381 0.600 ;
  LAYER ME1 ;
  RECT 356.061 0.000 356.381 0.600 ;
 END
 ANTENNAPARTIALMETALAREA                  5.273 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME3 ;
 ANTENNADIFFAREA                          1.293 LAYER ME4 ;
END DO78
PIN DI77
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 352.619 0.000 352.939 0.600 ;
  LAYER ME3 ;
  RECT 352.619 0.000 352.939 0.600 ;
  LAYER ME2 ;
  RECT 352.619 0.000 352.939 0.600 ;
  LAYER ME1 ;
  RECT 352.619 0.000 352.939 0.600 ;
 END
 ANTENNAPARTIALMETALAREA                  1.058 LAYER ME2 ;
 ANTENNAGATEAREA                          0.072 LAYER ME2 ;
 ANTENNAGATEAREA                          0.072 LAYER ME3 ;
 ANTENNAGATEAREA                          0.072 LAYER ME4 ;
 ANTENNADIFFAREA                          0.160 LAYER ME2 ;
 ANTENNADIFFAREA                          0.160 LAYER ME3 ;
 ANTENNADIFFAREA                          0.160 LAYER ME4 ;
 ANTENNAMAXAREACAR                       21.782 LAYER ME2 ;
 ANTENNAMAXAREACAR                       24.449 LAYER ME3 ;
 ANTENNAMAXAREACAR                       27.116 LAYER ME4 ;
END DI77
PIN DO77
  DIRECTION OUTPUT ;
 PORT
  LAYER ME4 ;
  RECT 352.057 0.000 352.377 0.600 ;
  LAYER ME3 ;
  RECT 352.057 0.000 352.377 0.600 ;
  LAYER ME2 ;
  RECT 352.057 0.000 352.377 0.600 ;
  LAYER ME1 ;
  RECT 352.057 0.000 352.377 0.600 ;
 END
 ANTENNAPARTIALMETALAREA                  5.273 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME3 ;
 ANTENNADIFFAREA                          1.293 LAYER ME4 ;
END DO77
PIN DI76
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 348.615 0.000 348.935 0.600 ;
  LAYER ME3 ;
  RECT 348.615 0.000 348.935 0.600 ;
  LAYER ME2 ;
  RECT 348.615 0.000 348.935 0.600 ;
  LAYER ME1 ;
  RECT 348.615 0.000 348.935 0.600 ;
 END
 ANTENNAPARTIALMETALAREA                  1.058 LAYER ME2 ;
 ANTENNAGATEAREA                          0.072 LAYER ME2 ;
 ANTENNAGATEAREA                          0.072 LAYER ME3 ;
 ANTENNAGATEAREA                          0.072 LAYER ME4 ;
 ANTENNADIFFAREA                          0.160 LAYER ME2 ;
 ANTENNADIFFAREA                          0.160 LAYER ME3 ;
 ANTENNADIFFAREA                          0.160 LAYER ME4 ;
 ANTENNAMAXAREACAR                       21.782 LAYER ME2 ;
 ANTENNAMAXAREACAR                       24.449 LAYER ME3 ;
 ANTENNAMAXAREACAR                       27.116 LAYER ME4 ;
END DI76
PIN DO76
  DIRECTION OUTPUT ;
 PORT
  LAYER ME4 ;
  RECT 348.053 0.000 348.373 0.600 ;
  LAYER ME3 ;
  RECT 348.053 0.000 348.373 0.600 ;
  LAYER ME2 ;
  RECT 348.053 0.000 348.373 0.600 ;
  LAYER ME1 ;
  RECT 348.053 0.000 348.373 0.600 ;
 END
 ANTENNAPARTIALMETALAREA                  5.273 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME3 ;
 ANTENNADIFFAREA                          1.293 LAYER ME4 ;
END DO76
PIN DI75
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 344.611 0.000 344.931 0.600 ;
  LAYER ME3 ;
  RECT 344.611 0.000 344.931 0.600 ;
  LAYER ME2 ;
  RECT 344.611 0.000 344.931 0.600 ;
  LAYER ME1 ;
  RECT 344.611 0.000 344.931 0.600 ;
 END
 ANTENNAPARTIALMETALAREA                  1.058 LAYER ME2 ;
 ANTENNAGATEAREA                          0.072 LAYER ME2 ;
 ANTENNAGATEAREA                          0.072 LAYER ME3 ;
 ANTENNAGATEAREA                          0.072 LAYER ME4 ;
 ANTENNADIFFAREA                          0.160 LAYER ME2 ;
 ANTENNADIFFAREA                          0.160 LAYER ME3 ;
 ANTENNADIFFAREA                          0.160 LAYER ME4 ;
 ANTENNAMAXAREACAR                       21.782 LAYER ME2 ;
 ANTENNAMAXAREACAR                       24.449 LAYER ME3 ;
 ANTENNAMAXAREACAR                       27.116 LAYER ME4 ;
END DI75
PIN DO75
  DIRECTION OUTPUT ;
 PORT
  LAYER ME4 ;
  RECT 344.049 0.000 344.369 0.600 ;
  LAYER ME3 ;
  RECT 344.049 0.000 344.369 0.600 ;
  LAYER ME2 ;
  RECT 344.049 0.000 344.369 0.600 ;
  LAYER ME1 ;
  RECT 344.049 0.000 344.369 0.600 ;
 END
 ANTENNAPARTIALMETALAREA                  5.273 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME3 ;
 ANTENNADIFFAREA                          1.293 LAYER ME4 ;
END DO75
PIN DI74
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 340.607 0.000 340.927 0.600 ;
  LAYER ME3 ;
  RECT 340.607 0.000 340.927 0.600 ;
  LAYER ME2 ;
  RECT 340.607 0.000 340.927 0.600 ;
  LAYER ME1 ;
  RECT 340.607 0.000 340.927 0.600 ;
 END
 ANTENNAPARTIALMETALAREA                  1.058 LAYER ME2 ;
 ANTENNAGATEAREA                          0.072 LAYER ME2 ;
 ANTENNAGATEAREA                          0.072 LAYER ME3 ;
 ANTENNAGATEAREA                          0.072 LAYER ME4 ;
 ANTENNADIFFAREA                          0.160 LAYER ME2 ;
 ANTENNADIFFAREA                          0.160 LAYER ME3 ;
 ANTENNADIFFAREA                          0.160 LAYER ME4 ;
 ANTENNAMAXAREACAR                       21.782 LAYER ME2 ;
 ANTENNAMAXAREACAR                       24.449 LAYER ME3 ;
 ANTENNAMAXAREACAR                       27.116 LAYER ME4 ;
END DI74
PIN DO74
  DIRECTION OUTPUT ;
 PORT
  LAYER ME4 ;
  RECT 340.045 0.000 340.365 0.600 ;
  LAYER ME3 ;
  RECT 340.045 0.000 340.365 0.600 ;
  LAYER ME2 ;
  RECT 340.045 0.000 340.365 0.600 ;
  LAYER ME1 ;
  RECT 340.045 0.000 340.365 0.600 ;
 END
 ANTENNAPARTIALMETALAREA                  5.273 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME3 ;
 ANTENNADIFFAREA                          1.293 LAYER ME4 ;
END DO74
PIN DI73
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 336.603 0.000 336.923 0.600 ;
  LAYER ME3 ;
  RECT 336.603 0.000 336.923 0.600 ;
  LAYER ME2 ;
  RECT 336.603 0.000 336.923 0.600 ;
  LAYER ME1 ;
  RECT 336.603 0.000 336.923 0.600 ;
 END
 ANTENNAPARTIALMETALAREA                  1.058 LAYER ME2 ;
 ANTENNAGATEAREA                          0.072 LAYER ME2 ;
 ANTENNAGATEAREA                          0.072 LAYER ME3 ;
 ANTENNAGATEAREA                          0.072 LAYER ME4 ;
 ANTENNADIFFAREA                          0.160 LAYER ME2 ;
 ANTENNADIFFAREA                          0.160 LAYER ME3 ;
 ANTENNADIFFAREA                          0.160 LAYER ME4 ;
 ANTENNAMAXAREACAR                       21.782 LAYER ME2 ;
 ANTENNAMAXAREACAR                       24.449 LAYER ME3 ;
 ANTENNAMAXAREACAR                       27.116 LAYER ME4 ;
END DI73
PIN DO73
  DIRECTION OUTPUT ;
 PORT
  LAYER ME4 ;
  RECT 336.041 0.000 336.361 0.600 ;
  LAYER ME3 ;
  RECT 336.041 0.000 336.361 0.600 ;
  LAYER ME2 ;
  RECT 336.041 0.000 336.361 0.600 ;
  LAYER ME1 ;
  RECT 336.041 0.000 336.361 0.600 ;
 END
 ANTENNAPARTIALMETALAREA                  5.273 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME3 ;
 ANTENNADIFFAREA                          1.293 LAYER ME4 ;
END DO73
PIN DI72
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 332.599 0.000 332.919 0.600 ;
  LAYER ME3 ;
  RECT 332.599 0.000 332.919 0.600 ;
  LAYER ME2 ;
  RECT 332.599 0.000 332.919 0.600 ;
  LAYER ME1 ;
  RECT 332.599 0.000 332.919 0.600 ;
 END
 ANTENNAPARTIALMETALAREA                  1.058 LAYER ME2 ;
 ANTENNAGATEAREA                          0.072 LAYER ME2 ;
 ANTENNAGATEAREA                          0.072 LAYER ME3 ;
 ANTENNAGATEAREA                          0.072 LAYER ME4 ;
 ANTENNADIFFAREA                          0.160 LAYER ME2 ;
 ANTENNADIFFAREA                          0.160 LAYER ME3 ;
 ANTENNADIFFAREA                          0.160 LAYER ME4 ;
 ANTENNAMAXAREACAR                       21.782 LAYER ME2 ;
 ANTENNAMAXAREACAR                       24.449 LAYER ME3 ;
 ANTENNAMAXAREACAR                       27.116 LAYER ME4 ;
END DI72
PIN DO72
  DIRECTION OUTPUT ;
 PORT
  LAYER ME4 ;
  RECT 332.037 0.000 332.357 0.600 ;
  LAYER ME3 ;
  RECT 332.037 0.000 332.357 0.600 ;
  LAYER ME2 ;
  RECT 332.037 0.000 332.357 0.600 ;
  LAYER ME1 ;
  RECT 332.037 0.000 332.357 0.600 ;
 END
 ANTENNAPARTIALMETALAREA                  5.273 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME3 ;
 ANTENNADIFFAREA                          1.293 LAYER ME4 ;
END DO72
PIN DI71
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 328.595 0.000 328.915 0.600 ;
  LAYER ME3 ;
  RECT 328.595 0.000 328.915 0.600 ;
  LAYER ME2 ;
  RECT 328.595 0.000 328.915 0.600 ;
  LAYER ME1 ;
  RECT 328.595 0.000 328.915 0.600 ;
 END
 ANTENNAPARTIALMETALAREA                  1.058 LAYER ME2 ;
 ANTENNAGATEAREA                          0.072 LAYER ME2 ;
 ANTENNAGATEAREA                          0.072 LAYER ME3 ;
 ANTENNAGATEAREA                          0.072 LAYER ME4 ;
 ANTENNADIFFAREA                          0.160 LAYER ME2 ;
 ANTENNADIFFAREA                          0.160 LAYER ME3 ;
 ANTENNADIFFAREA                          0.160 LAYER ME4 ;
 ANTENNAMAXAREACAR                       21.782 LAYER ME2 ;
 ANTENNAMAXAREACAR                       24.449 LAYER ME3 ;
 ANTENNAMAXAREACAR                       27.116 LAYER ME4 ;
END DI71
PIN DO71
  DIRECTION OUTPUT ;
 PORT
  LAYER ME4 ;
  RECT 328.033 0.000 328.353 0.600 ;
  LAYER ME3 ;
  RECT 328.033 0.000 328.353 0.600 ;
  LAYER ME2 ;
  RECT 328.033 0.000 328.353 0.600 ;
  LAYER ME1 ;
  RECT 328.033 0.000 328.353 0.600 ;
 END
 ANTENNAPARTIALMETALAREA                  5.273 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME3 ;
 ANTENNADIFFAREA                          1.293 LAYER ME4 ;
END DO71
PIN DI70
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 324.591 0.000 324.911 0.600 ;
  LAYER ME3 ;
  RECT 324.591 0.000 324.911 0.600 ;
  LAYER ME2 ;
  RECT 324.591 0.000 324.911 0.600 ;
  LAYER ME1 ;
  RECT 324.591 0.000 324.911 0.600 ;
 END
 ANTENNAPARTIALMETALAREA                  1.058 LAYER ME2 ;
 ANTENNAGATEAREA                          0.072 LAYER ME2 ;
 ANTENNAGATEAREA                          0.072 LAYER ME3 ;
 ANTENNAGATEAREA                          0.072 LAYER ME4 ;
 ANTENNADIFFAREA                          0.160 LAYER ME2 ;
 ANTENNADIFFAREA                          0.160 LAYER ME3 ;
 ANTENNADIFFAREA                          0.160 LAYER ME4 ;
 ANTENNAMAXAREACAR                       21.782 LAYER ME2 ;
 ANTENNAMAXAREACAR                       24.449 LAYER ME3 ;
 ANTENNAMAXAREACAR                       27.116 LAYER ME4 ;
END DI70
PIN DO70
  DIRECTION OUTPUT ;
 PORT
  LAYER ME4 ;
  RECT 324.029 0.000 324.349 0.600 ;
  LAYER ME3 ;
  RECT 324.029 0.000 324.349 0.600 ;
  LAYER ME2 ;
  RECT 324.029 0.000 324.349 0.600 ;
  LAYER ME1 ;
  RECT 324.029 0.000 324.349 0.600 ;
 END
 ANTENNAPARTIALMETALAREA                  5.273 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME3 ;
 ANTENNADIFFAREA                          1.293 LAYER ME4 ;
END DO70
PIN DI69
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 320.587 0.000 320.907 0.600 ;
  LAYER ME3 ;
  RECT 320.587 0.000 320.907 0.600 ;
  LAYER ME2 ;
  RECT 320.587 0.000 320.907 0.600 ;
  LAYER ME1 ;
  RECT 320.587 0.000 320.907 0.600 ;
 END
 ANTENNAPARTIALMETALAREA                  1.058 LAYER ME2 ;
 ANTENNAGATEAREA                          0.072 LAYER ME2 ;
 ANTENNAGATEAREA                          0.072 LAYER ME3 ;
 ANTENNAGATEAREA                          0.072 LAYER ME4 ;
 ANTENNADIFFAREA                          0.160 LAYER ME2 ;
 ANTENNADIFFAREA                          0.160 LAYER ME3 ;
 ANTENNADIFFAREA                          0.160 LAYER ME4 ;
 ANTENNAMAXAREACAR                       21.782 LAYER ME2 ;
 ANTENNAMAXAREACAR                       24.449 LAYER ME3 ;
 ANTENNAMAXAREACAR                       27.116 LAYER ME4 ;
END DI69
PIN DO69
  DIRECTION OUTPUT ;
 PORT
  LAYER ME4 ;
  RECT 320.025 0.000 320.345 0.600 ;
  LAYER ME3 ;
  RECT 320.025 0.000 320.345 0.600 ;
  LAYER ME2 ;
  RECT 320.025 0.000 320.345 0.600 ;
  LAYER ME1 ;
  RECT 320.025 0.000 320.345 0.600 ;
 END
 ANTENNAPARTIALMETALAREA                  5.273 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME3 ;
 ANTENNADIFFAREA                          1.293 LAYER ME4 ;
END DO69
PIN DI68
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 316.583 0.000 316.903 0.600 ;
  LAYER ME3 ;
  RECT 316.583 0.000 316.903 0.600 ;
  LAYER ME2 ;
  RECT 316.583 0.000 316.903 0.600 ;
  LAYER ME1 ;
  RECT 316.583 0.000 316.903 0.600 ;
 END
 ANTENNAPARTIALMETALAREA                  1.058 LAYER ME2 ;
 ANTENNAGATEAREA                          0.072 LAYER ME2 ;
 ANTENNAGATEAREA                          0.072 LAYER ME3 ;
 ANTENNAGATEAREA                          0.072 LAYER ME4 ;
 ANTENNADIFFAREA                          0.160 LAYER ME2 ;
 ANTENNADIFFAREA                          0.160 LAYER ME3 ;
 ANTENNADIFFAREA                          0.160 LAYER ME4 ;
 ANTENNAMAXAREACAR                       21.782 LAYER ME2 ;
 ANTENNAMAXAREACAR                       24.449 LAYER ME3 ;
 ANTENNAMAXAREACAR                       27.116 LAYER ME4 ;
END DI68
PIN DO68
  DIRECTION OUTPUT ;
 PORT
  LAYER ME4 ;
  RECT 316.021 0.000 316.341 0.600 ;
  LAYER ME3 ;
  RECT 316.021 0.000 316.341 0.600 ;
  LAYER ME2 ;
  RECT 316.021 0.000 316.341 0.600 ;
  LAYER ME1 ;
  RECT 316.021 0.000 316.341 0.600 ;
 END
 ANTENNAPARTIALMETALAREA                  5.273 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME3 ;
 ANTENNADIFFAREA                          1.293 LAYER ME4 ;
END DO68
PIN DI67
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 312.579 0.000 312.899 0.600 ;
  LAYER ME3 ;
  RECT 312.579 0.000 312.899 0.600 ;
  LAYER ME2 ;
  RECT 312.579 0.000 312.899 0.600 ;
  LAYER ME1 ;
  RECT 312.579 0.000 312.899 0.600 ;
 END
 ANTENNAPARTIALMETALAREA                  1.058 LAYER ME2 ;
 ANTENNAGATEAREA                          0.072 LAYER ME2 ;
 ANTENNAGATEAREA                          0.072 LAYER ME3 ;
 ANTENNAGATEAREA                          0.072 LAYER ME4 ;
 ANTENNADIFFAREA                          0.160 LAYER ME2 ;
 ANTENNADIFFAREA                          0.160 LAYER ME3 ;
 ANTENNADIFFAREA                          0.160 LAYER ME4 ;
 ANTENNAMAXAREACAR                       21.782 LAYER ME2 ;
 ANTENNAMAXAREACAR                       24.449 LAYER ME3 ;
 ANTENNAMAXAREACAR                       27.116 LAYER ME4 ;
END DI67
PIN DO67
  DIRECTION OUTPUT ;
 PORT
  LAYER ME4 ;
  RECT 312.017 0.000 312.337 0.600 ;
  LAYER ME3 ;
  RECT 312.017 0.000 312.337 0.600 ;
  LAYER ME2 ;
  RECT 312.017 0.000 312.337 0.600 ;
  LAYER ME1 ;
  RECT 312.017 0.000 312.337 0.600 ;
 END
 ANTENNAPARTIALMETALAREA                  5.273 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME3 ;
 ANTENNADIFFAREA                          1.293 LAYER ME4 ;
END DO67
PIN DI66
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 308.575 0.000 308.895 0.600 ;
  LAYER ME3 ;
  RECT 308.575 0.000 308.895 0.600 ;
  LAYER ME2 ;
  RECT 308.575 0.000 308.895 0.600 ;
  LAYER ME1 ;
  RECT 308.575 0.000 308.895 0.600 ;
 END
 ANTENNAPARTIALMETALAREA                  1.058 LAYER ME2 ;
 ANTENNAGATEAREA                          0.072 LAYER ME2 ;
 ANTENNAGATEAREA                          0.072 LAYER ME3 ;
 ANTENNAGATEAREA                          0.072 LAYER ME4 ;
 ANTENNADIFFAREA                          0.160 LAYER ME2 ;
 ANTENNADIFFAREA                          0.160 LAYER ME3 ;
 ANTENNADIFFAREA                          0.160 LAYER ME4 ;
 ANTENNAMAXAREACAR                       21.782 LAYER ME2 ;
 ANTENNAMAXAREACAR                       24.449 LAYER ME3 ;
 ANTENNAMAXAREACAR                       27.116 LAYER ME4 ;
END DI66
PIN DO66
  DIRECTION OUTPUT ;
 PORT
  LAYER ME4 ;
  RECT 308.013 0.000 308.333 0.600 ;
  LAYER ME3 ;
  RECT 308.013 0.000 308.333 0.600 ;
  LAYER ME2 ;
  RECT 308.013 0.000 308.333 0.600 ;
  LAYER ME1 ;
  RECT 308.013 0.000 308.333 0.600 ;
 END
 ANTENNAPARTIALMETALAREA                  5.273 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME3 ;
 ANTENNADIFFAREA                          1.293 LAYER ME4 ;
END DO66
PIN DI65
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 304.571 0.000 304.891 0.600 ;
  LAYER ME3 ;
  RECT 304.571 0.000 304.891 0.600 ;
  LAYER ME2 ;
  RECT 304.571 0.000 304.891 0.600 ;
  LAYER ME1 ;
  RECT 304.571 0.000 304.891 0.600 ;
 END
 ANTENNAPARTIALMETALAREA                  1.058 LAYER ME2 ;
 ANTENNAGATEAREA                          0.072 LAYER ME2 ;
 ANTENNAGATEAREA                          0.072 LAYER ME3 ;
 ANTENNAGATEAREA                          0.072 LAYER ME4 ;
 ANTENNADIFFAREA                          0.160 LAYER ME2 ;
 ANTENNADIFFAREA                          0.160 LAYER ME3 ;
 ANTENNADIFFAREA                          0.160 LAYER ME4 ;
 ANTENNAMAXAREACAR                       21.782 LAYER ME2 ;
 ANTENNAMAXAREACAR                       24.449 LAYER ME3 ;
 ANTENNAMAXAREACAR                       27.116 LAYER ME4 ;
END DI65
PIN DO65
  DIRECTION OUTPUT ;
 PORT
  LAYER ME4 ;
  RECT 304.009 0.000 304.329 0.600 ;
  LAYER ME3 ;
  RECT 304.009 0.000 304.329 0.600 ;
  LAYER ME2 ;
  RECT 304.009 0.000 304.329 0.600 ;
  LAYER ME1 ;
  RECT 304.009 0.000 304.329 0.600 ;
 END
 ANTENNAPARTIALMETALAREA                  5.273 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME3 ;
 ANTENNADIFFAREA                          1.293 LAYER ME4 ;
END DO65
PIN DI64
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 300.005 0.000 300.325 0.600 ;
  LAYER ME3 ;
  RECT 300.005 0.000 300.325 0.600 ;
  LAYER ME2 ;
  RECT 300.005 0.000 300.325 0.600 ;
  LAYER ME1 ;
  RECT 300.005 0.000 300.325 0.600 ;
 END
 ANTENNAPARTIALMETALAREA                  0.346 LAYER ME1 ;
 ANTENNAPARTIALMETALAREA                  1.466 LAYER ME2 ;
 ANTENNAPARTIALMETALAREA                  0.508 LAYER ME3 ;
 ANTENNAGATEAREA                          0.072 LAYER ME3 ;
 ANTENNAGATEAREA                          0.072 LAYER ME4 ;
 ANTENNADIFFAREA                          0.218 LAYER ME1 ;
 ANTENNADIFFAREA                          0.218 LAYER ME2 ;
 ANTENNADIFFAREA                          0.218 LAYER ME3 ;
 ANTENNADIFFAREA                          0.218 LAYER ME4 ;
 ANTENNAMAXAREACAR                       17.267 LAYER ME3 ;
 ANTENNAMAXAREACAR                       19.933 LAYER ME4 ;
END DI64
PIN DO64
  DIRECTION OUTPUT ;
 PORT
  LAYER ME4 ;
  RECT 300.567 0.000 300.887 0.600 ;
  LAYER ME3 ;
  RECT 300.567 0.000 300.887 0.600 ;
  LAYER ME2 ;
  RECT 300.567 0.000 300.887 0.600 ;
  LAYER ME1 ;
  RECT 300.567 0.000 300.887 0.600 ;
 END
 ANTENNAPARTIALMETALAREA                  5.602 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME3 ;
 ANTENNADIFFAREA                          1.293 LAYER ME4 ;
END DO64
PIN WEB4
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 298.565 0.000 298.885 0.600 ;
  LAYER ME3 ;
  RECT 298.565 0.000 298.885 0.600 ;
  LAYER ME2 ;
  RECT 298.565 0.000 298.885 0.600 ;
  LAYER ME1 ;
  RECT 298.565 0.000 298.885 0.600 ;
 END
 ANTENNAPARTIALMETALAREA                  1.036 LAYER ME2 ;
 ANTENNAGATEAREA                          0.288 LAYER ME2 ;
 ANTENNAGATEAREA                          0.288 LAYER ME3 ;
 ANTENNAGATEAREA                          0.288 LAYER ME4 ;
 ANTENNADIFFAREA                          0.206 LAYER ME2 ;
 ANTENNADIFFAREA                          0.206 LAYER ME3 ;
 ANTENNADIFFAREA                          0.206 LAYER ME4 ;
 ANTENNAMAXAREACAR                        5.844 LAYER ME2 ;
 ANTENNAMAXAREACAR                        6.511 LAYER ME3 ;
 ANTENNAMAXAREACAR                        7.178 LAYER ME4 ;
END WEB4
OBS
  LAYER ME3 SPACING 0.260 ;
  RECT 0.000 0.000 557.611 293.175 ;
  LAYER ME2 SPACING 0.260 ;
  RECT 0.000 0.000 557.611 293.175 ;
  LAYER ME1 SPACING 0.260 ;
  RECT 0.000 0.000 557.611 293.175 ;
  LAYER ME4 SPACING 0.260 ;
  RECT 0.000 0.000 273.598 293.175 ;
  LAYER ME4 SPACING 0.260 ;
  RECT 275.252 0.000 276.372 293.175 ;
  LAYER ME4 SPACING 0.260 ;
  RECT 277.967 0.000 278.687 293.175 ;
  LAYER ME4 SPACING 0.260 ;
  RECT 279.417 0.000 280.137 293.175 ;
  LAYER ME4 SPACING 0.260 ;
  RECT 282.197 0.000 282.797 293.175 ;
  LAYER ME4 SPACING 0.260 ;
  RECT 285.411 0.000 287.097 293.175 ;
  LAYER ME4 SPACING 0.260 ;
  RECT 288.487 0.000 289.607 293.175 ;
  LAYER ME4 SPACING 0.260 ;
  RECT 290.882 0.000 291.602 293.175 ;
  LAYER ME4 SPACING 0.260 ;
  RECT 292.597 0.000 293.317 293.175 ;
  LAYER ME4 SPACING 0.260 ;
  RECT 294.517 0.000 557.611 293.175 ;
END
END SYKB110_512X16X8CM2
END LIBRARY





