# ________________________________________________________________________________________________
# 
# 
#             Synchronous One-Port Register File Compiler
# 
#                 UMC 0.11um LL AE Logic Process
# 
# ________________________________________________________________________________________________
# 
#               
#         Copyright (C) 2024 Faraday Technology Corporation. All Rights Reserved.       
#                
#         This source code is an unpublished work belongs to Faraday Technology Corporation       
#         It is considered a trade secret and is not to be divulged or       
#         used by parties who have not received written authorization from       
#         Faraday Technology Corporation       
#                
#         Faraday's home page can be found at: http://www.faraday-tech.com/       
#                
# ________________________________________________________________________________________________
# 
#        IP Name            :  FSR0K_B_SY                
#        IP Version         :  1.4.0                     
#        IP Release Status  :  Active                    
#        Word               :  128                       
#        Bit                :  2                         
#        Byte               :  8                         
#        Mux                :  4                         
#        Output Loading     :  0.01                      
#        Clock Input Slew   :  0.016                     
#        Data Input Slew    :  0.016                     
#        Ring Type          :  Ringless Model            
#        Ring Width         :  0                         
#        Bus Format         :  0                         
#        Memaker Path       :  /home/mem/Desktop/memlib  
#        GUI Version        :  m20230904                 
#        Date               :  2024/09/10 14:30:15       
# ________________________________________________________________________________________________
# 

VERSION 5.5 ;
NAMESCASESENSITIVE ON ;
MACRO SYKB110_128X2X8CM4
CLASS BLOCK ;
FOREIGN SYKB110_128X2X8CM4 0.000 0.000 ;
ORIGIN 0.000 0.000 ;
SIZE 171.627 BY 68.179 ;
SYMMETRY x y r90 ;
SITE core ;
PIN VCC
  DIRECTION INOUT ;
  USE POWER ;
 PORT
  LAYER ME4 ;
  RECT 109.297 0.000 110.017 33.870 ;
 END
 PORT
  LAYER ME4 ;
  RECT 105.293 0.000 106.013 33.870 ;
 END
 PORT
  LAYER ME4 ;
  RECT 117.305 0.000 118.025 33.870 ;
 END
 PORT
  LAYER ME4 ;
  RECT 113.301 0.000 114.021 33.870 ;
 END
 PORT
  LAYER ME4 ;
  RECT 125.313 0.000 126.033 33.870 ;
 END
 PORT
  LAYER ME4 ;
  RECT 121.309 0.000 122.029 33.870 ;
 END
 PORT
  LAYER ME4 ;
  RECT 133.321 0.000 134.041 33.870 ;
 END
 PORT
  LAYER ME4 ;
  RECT 129.317 0.000 130.037 33.870 ;
 END
 PORT
  LAYER ME4 ;
  RECT 141.329 0.000 142.049 33.870 ;
 END
 PORT
  LAYER ME4 ;
  RECT 137.325 0.000 138.045 33.870 ;
 END
 PORT
  LAYER ME4 ;
  RECT 149.337 0.000 150.057 33.870 ;
 END
 PORT
  LAYER ME4 ;
  RECT 145.333 0.000 146.053 33.870 ;
 END
 PORT
  LAYER ME4 ;
  RECT 157.345 0.000 158.065 33.870 ;
 END
 PORT
  LAYER ME4 ;
  RECT 153.341 0.000 154.061 33.870 ;
 END
 PORT
  LAYER ME4 ;
  RECT 165.353 0.000 166.073 33.870 ;
 END
 PORT
  LAYER ME4 ;
  RECT 161.349 0.000 162.069 33.870 ;
 END
 PORT
  LAYER ME4 ;
  RECT 170.327 0.000 170.707 68.179 ;
 END
 PORT
  LAYER ME4 ;
  RECT 88.405 0.000 89.005 68.179 ;
 END
 PORT
  LAYER ME4 ;
  RECT 92.585 0.000 93.305 68.179 ;
 END
 PORT
  LAYER ME4 ;
  RECT 94.695 0.000 95.815 68.179 ;
 END
 PORT
  LAYER ME4 ;
  RECT 100.725 0.000 101.445 68.179 ;
 END
 PORT
  LAYER ME4 ;
  RECT 102.661 0.921 103.041 68.179 ;
 END
 PORT
  LAYER ME4 ;
  RECT 81.460 0.000 82.580 68.179 ;
 END
 PORT
  LAYER ME4 ;
  RECT 84.175 0.000 84.895 68.179 ;
 END
 PORT
  LAYER ME4 ;
  RECT 79.086 0.000 79.806 67.420 ;
 END
 PORT
  LAYER ME4 ;
  RECT 77.046 0.921 77.766 68.179 ;
 END
 PORT
  LAYER ME4 ;
  RECT 74.926 0.000 75.646 68.179 ;
 END
 PORT
  LAYER ME4 ;
  RECT 72.886 0.921 73.606 68.179 ;
 END
 PORT
  LAYER ME4 ;
  RECT 0.920 0.000 1.300 68.179 ;
 END
 PORT
  LAYER ME4 ;
  RECT 7.556 0.000 8.276 33.870 ;
 END
 PORT
  LAYER ME4 ;
  RECT 3.552 0.000 4.272 33.870 ;
 END
 PORT
  LAYER ME4 ;
  RECT 15.564 0.000 16.284 33.870 ;
 END
 PORT
  LAYER ME4 ;
  RECT 11.560 0.000 12.280 33.870 ;
 END
 PORT
  LAYER ME4 ;
  RECT 23.572 0.000 24.292 33.870 ;
 END
 PORT
  LAYER ME4 ;
  RECT 19.568 0.000 20.288 33.870 ;
 END
 PORT
  LAYER ME4 ;
  RECT 31.580 0.000 32.300 33.870 ;
 END
 PORT
  LAYER ME4 ;
  RECT 27.576 0.000 28.296 33.870 ;
 END
 PORT
  LAYER ME4 ;
  RECT 39.588 0.000 40.308 33.870 ;
 END
 PORT
  LAYER ME4 ;
  RECT 35.584 0.000 36.304 33.870 ;
 END
 PORT
  LAYER ME4 ;
  RECT 47.596 0.000 48.316 33.870 ;
 END
 PORT
  LAYER ME4 ;
  RECT 43.592 0.000 44.312 33.870 ;
 END
 PORT
  LAYER ME4 ;
  RECT 55.604 0.000 56.324 33.870 ;
 END
 PORT
  LAYER ME4 ;
  RECT 51.600 0.000 52.320 33.870 ;
 END
 PORT
  LAYER ME4 ;
  RECT 63.612 0.000 64.332 33.870 ;
 END
 PORT
  LAYER ME4 ;
  RECT 59.608 0.000 60.328 33.870 ;
 END
 PORT
  LAYER ME4 ;
  RECT 70.766 0.000 71.486 68.179 ;
 END
 PORT
  LAYER ME4 ;
  RECT 68.586 0.000 68.966 68.179 ;
 END
 PORT
  LAYER ME4 ;
  RECT 111.489 35.220 111.829 68.179 ;
 END
 PORT
  LAYER ME4 ;
  RECT 109.487 35.220 109.827 68.179 ;
 END
 PORT
  LAYER ME4 ;
  RECT 107.485 35.220 107.825 68.179 ;
 END
 PORT
  LAYER ME4 ;
  RECT 105.483 35.220 105.823 68.179 ;
 END
 PORT
  LAYER ME4 ;
  RECT 119.497 35.220 119.837 68.179 ;
 END
 PORT
  LAYER ME4 ;
  RECT 117.495 35.220 117.835 68.179 ;
 END
 PORT
  LAYER ME4 ;
  RECT 115.493 35.220 115.833 68.179 ;
 END
 PORT
  LAYER ME4 ;
  RECT 113.491 35.220 113.831 68.179 ;
 END
 PORT
  LAYER ME4 ;
  RECT 127.505 35.220 127.845 68.179 ;
 END
 PORT
  LAYER ME4 ;
  RECT 125.503 35.220 125.843 68.179 ;
 END
 PORT
  LAYER ME4 ;
  RECT 123.501 35.220 123.841 68.179 ;
 END
 PORT
  LAYER ME4 ;
  RECT 121.499 35.220 121.839 68.179 ;
 END
 PORT
  LAYER ME4 ;
  RECT 135.513 35.220 135.853 68.179 ;
 END
 PORT
  LAYER ME4 ;
  RECT 133.511 35.220 133.851 68.179 ;
 END
 PORT
  LAYER ME4 ;
  RECT 131.509 35.220 131.849 68.179 ;
 END
 PORT
  LAYER ME4 ;
  RECT 129.507 35.220 129.847 68.179 ;
 END
 PORT
  LAYER ME4 ;
  RECT 143.521 35.220 143.861 68.179 ;
 END
 PORT
  LAYER ME4 ;
  RECT 141.519 35.220 141.859 68.179 ;
 END
 PORT
  LAYER ME4 ;
  RECT 139.517 35.220 139.857 68.179 ;
 END
 PORT
  LAYER ME4 ;
  RECT 137.515 35.220 137.855 68.179 ;
 END
 PORT
  LAYER ME4 ;
  RECT 151.529 35.220 151.869 68.179 ;
 END
 PORT
  LAYER ME4 ;
  RECT 149.527 35.220 149.867 68.179 ;
 END
 PORT
  LAYER ME4 ;
  RECT 147.525 35.220 147.865 68.179 ;
 END
 PORT
  LAYER ME4 ;
  RECT 145.523 35.220 145.863 68.179 ;
 END
 PORT
  LAYER ME4 ;
  RECT 159.537 35.220 159.877 68.179 ;
 END
 PORT
  LAYER ME4 ;
  RECT 157.535 35.220 157.875 68.179 ;
 END
 PORT
  LAYER ME4 ;
  RECT 155.533 35.220 155.873 68.179 ;
 END
 PORT
  LAYER ME4 ;
  RECT 153.531 35.220 153.871 68.179 ;
 END
 PORT
  LAYER ME4 ;
  RECT 167.545 35.220 167.885 68.179 ;
 END
 PORT
  LAYER ME4 ;
  RECT 165.543 35.220 165.883 68.179 ;
 END
 PORT
  LAYER ME4 ;
  RECT 163.541 35.220 163.881 68.179 ;
 END
 PORT
  LAYER ME4 ;
  RECT 161.539 35.220 161.879 68.179 ;
 END
 PORT
  LAYER ME4 ;
  RECT 9.748 35.220 10.088 68.179 ;
 END
 PORT
  LAYER ME4 ;
  RECT 7.746 35.220 8.086 68.179 ;
 END
 PORT
  LAYER ME4 ;
  RECT 5.744 35.220 6.084 68.179 ;
 END
 PORT
  LAYER ME4 ;
  RECT 3.742 35.220 4.082 68.179 ;
 END
 PORT
  LAYER ME4 ;
  RECT 17.756 35.220 18.096 68.179 ;
 END
 PORT
  LAYER ME4 ;
  RECT 15.754 35.220 16.094 68.179 ;
 END
 PORT
  LAYER ME4 ;
  RECT 13.752 35.220 14.092 68.179 ;
 END
 PORT
  LAYER ME4 ;
  RECT 11.750 35.220 12.090 68.179 ;
 END
 PORT
  LAYER ME4 ;
  RECT 25.764 35.220 26.104 68.179 ;
 END
 PORT
  LAYER ME4 ;
  RECT 23.762 35.220 24.102 68.179 ;
 END
 PORT
  LAYER ME4 ;
  RECT 21.760 35.220 22.100 68.179 ;
 END
 PORT
  LAYER ME4 ;
  RECT 19.758 35.220 20.098 68.179 ;
 END
 PORT
  LAYER ME4 ;
  RECT 33.772 35.220 34.112 68.179 ;
 END
 PORT
  LAYER ME4 ;
  RECT 31.770 35.220 32.110 68.179 ;
 END
 PORT
  LAYER ME4 ;
  RECT 29.768 35.220 30.108 68.179 ;
 END
 PORT
  LAYER ME4 ;
  RECT 27.766 35.220 28.106 68.179 ;
 END
 PORT
  LAYER ME4 ;
  RECT 41.780 35.220 42.120 68.179 ;
 END
 PORT
  LAYER ME4 ;
  RECT 39.778 35.220 40.118 68.179 ;
 END
 PORT
  LAYER ME4 ;
  RECT 37.776 35.220 38.116 68.179 ;
 END
 PORT
  LAYER ME4 ;
  RECT 35.774 35.220 36.114 68.179 ;
 END
 PORT
  LAYER ME4 ;
  RECT 49.788 35.220 50.128 68.179 ;
 END
 PORT
  LAYER ME4 ;
  RECT 47.786 35.220 48.126 68.179 ;
 END
 PORT
  LAYER ME4 ;
  RECT 45.784 35.220 46.124 68.179 ;
 END
 PORT
  LAYER ME4 ;
  RECT 43.782 35.220 44.122 68.179 ;
 END
 PORT
  LAYER ME4 ;
  RECT 57.796 35.220 58.136 68.179 ;
 END
 PORT
  LAYER ME4 ;
  RECT 55.794 35.220 56.134 68.179 ;
 END
 PORT
  LAYER ME4 ;
  RECT 53.792 35.220 54.132 68.179 ;
 END
 PORT
  LAYER ME4 ;
  RECT 51.790 35.220 52.130 68.179 ;
 END
 PORT
  LAYER ME4 ;
  RECT 65.804 35.220 66.144 68.179 ;
 END
 PORT
  LAYER ME4 ;
  RECT 63.802 35.220 64.142 68.179 ;
 END
 PORT
  LAYER ME4 ;
  RECT 61.800 35.220 62.140 68.179 ;
 END
 PORT
  LAYER ME4 ;
  RECT 59.798 35.220 60.138 68.179 ;
 END
END VCC
PIN GND
  DIRECTION INOUT ;
  USE GROUND ;
 PORT
  LAYER ME4 ;
  RECT 104.482 0.921 104.822 68.179 ;
 END
 PORT
  LAYER ME4 ;
  RECT 111.299 0.000 112.019 31.570 ;
 END
 PORT
  LAYER ME4 ;
  RECT 112.490 0.000 112.830 68.179 ;
 END
 PORT
  LAYER ME4 ;
  RECT 106.484 0.000 106.824 68.179 ;
 END
 PORT
  LAYER ME4 ;
  RECT 107.295 0.000 108.015 31.570 ;
 END
 PORT
  LAYER ME4 ;
  RECT 108.486 0.921 108.826 68.179 ;
 END
 PORT
  LAYER ME4 ;
  RECT 110.488 0.921 110.828 68.179 ;
 END
 PORT
  LAYER ME4 ;
  RECT 119.307 0.000 120.027 31.570 ;
 END
 PORT
  LAYER ME4 ;
  RECT 120.498 0.000 120.838 68.179 ;
 END
 PORT
  LAYER ME4 ;
  RECT 114.492 0.000 114.832 68.179 ;
 END
 PORT
  LAYER ME4 ;
  RECT 115.303 0.000 116.023 31.570 ;
 END
 PORT
  LAYER ME4 ;
  RECT 116.494 0.921 116.834 68.179 ;
 END
 PORT
  LAYER ME4 ;
  RECT 118.496 0.921 118.836 68.179 ;
 END
 PORT
  LAYER ME4 ;
  RECT 127.315 0.000 128.035 31.570 ;
 END
 PORT
  LAYER ME4 ;
  RECT 128.506 0.000 128.846 68.179 ;
 END
 PORT
  LAYER ME4 ;
  RECT 122.500 0.000 122.840 68.179 ;
 END
 PORT
  LAYER ME4 ;
  RECT 123.311 0.000 124.031 31.570 ;
 END
 PORT
  LAYER ME4 ;
  RECT 124.502 0.921 124.842 68.179 ;
 END
 PORT
  LAYER ME4 ;
  RECT 126.504 0.921 126.844 68.179 ;
 END
 PORT
  LAYER ME4 ;
  RECT 135.323 0.000 136.043 31.570 ;
 END
 PORT
  LAYER ME4 ;
  RECT 136.514 0.000 136.854 68.179 ;
 END
 PORT
  LAYER ME4 ;
  RECT 130.508 0.000 130.848 68.179 ;
 END
 PORT
  LAYER ME4 ;
  RECT 131.319 0.000 132.039 31.570 ;
 END
 PORT
  LAYER ME4 ;
  RECT 132.510 0.921 132.850 68.179 ;
 END
 PORT
  LAYER ME4 ;
  RECT 134.512 0.921 134.852 68.179 ;
 END
 PORT
  LAYER ME4 ;
  RECT 143.331 0.000 144.051 31.570 ;
 END
 PORT
  LAYER ME4 ;
  RECT 144.522 0.000 144.862 68.179 ;
 END
 PORT
  LAYER ME4 ;
  RECT 138.516 0.000 138.856 68.179 ;
 END
 PORT
  LAYER ME4 ;
  RECT 139.327 0.000 140.047 31.570 ;
 END
 PORT
  LAYER ME4 ;
  RECT 140.518 0.921 140.858 68.179 ;
 END
 PORT
  LAYER ME4 ;
  RECT 142.520 0.921 142.860 68.179 ;
 END
 PORT
  LAYER ME4 ;
  RECT 151.339 0.000 152.059 31.570 ;
 END
 PORT
  LAYER ME4 ;
  RECT 152.530 0.000 152.870 68.179 ;
 END
 PORT
  LAYER ME4 ;
  RECT 146.524 0.000 146.864 68.179 ;
 END
 PORT
  LAYER ME4 ;
  RECT 147.335 0.000 148.055 31.570 ;
 END
 PORT
  LAYER ME4 ;
  RECT 148.526 0.921 148.866 68.179 ;
 END
 PORT
  LAYER ME4 ;
  RECT 150.528 0.921 150.868 68.179 ;
 END
 PORT
  LAYER ME4 ;
  RECT 159.347 0.000 160.067 31.570 ;
 END
 PORT
  LAYER ME4 ;
  RECT 160.538 0.000 160.878 68.179 ;
 END
 PORT
  LAYER ME4 ;
  RECT 154.532 0.000 154.872 68.179 ;
 END
 PORT
  LAYER ME4 ;
  RECT 155.343 0.000 156.063 31.570 ;
 END
 PORT
  LAYER ME4 ;
  RECT 156.534 0.921 156.874 68.179 ;
 END
 PORT
  LAYER ME4 ;
  RECT 158.536 0.921 158.876 68.179 ;
 END
 PORT
  LAYER ME4 ;
  RECT 167.355 0.000 168.075 31.570 ;
 END
 PORT
  LAYER ME4 ;
  RECT 168.546 0.000 168.886 68.179 ;
 END
 PORT
  LAYER ME4 ;
  RECT 162.540 0.000 162.880 68.179 ;
 END
 PORT
  LAYER ME4 ;
  RECT 163.351 0.000 164.071 31.570 ;
 END
 PORT
  LAYER ME4 ;
  RECT 164.542 0.921 164.882 68.179 ;
 END
 PORT
  LAYER ME4 ;
  RECT 166.544 0.921 166.884 68.179 ;
 END
 PORT
  LAYER ME4 ;
  RECT 169.547 0.000 169.887 68.179 ;
 END
 PORT
  LAYER ME4 ;
  RECT 85.625 0.000 86.345 68.179 ;
 END
 PORT
  LAYER ME4 ;
  RECT 91.619 0.000 92.339 68.179 ;
 END
 PORT
  LAYER ME4 ;
  RECT 97.090 0.000 97.810 68.179 ;
 END
 PORT
  LAYER ME4 ;
  RECT 98.805 0.000 99.525 68.179 ;
 END
 PORT
  LAYER ME4 ;
  RECT 101.801 0.000 102.401 68.179 ;
 END
 PORT
  LAYER ME4 ;
  RECT 103.481 0.921 103.821 68.179 ;
 END
 PORT
  LAYER ME4 ;
  RECT 78.066 0.000 78.786 68.179 ;
 END
 PORT
  LAYER ME4 ;
  RECT 76.026 0.921 76.746 67.420 ;
 END
 PORT
  LAYER ME4 ;
  RECT 73.906 0.000 74.626 68.179 ;
 END
 PORT
  LAYER ME4 ;
  RECT 71.866 0.921 72.586 68.179 ;
 END
 PORT
  LAYER ME4 ;
  RECT 1.740 0.000 2.080 68.179 ;
 END
 PORT
  LAYER ME4 ;
  RECT 2.741 0.921 3.081 68.179 ;
 END
 PORT
  LAYER ME4 ;
  RECT 9.558 0.000 10.278 31.570 ;
 END
 PORT
  LAYER ME4 ;
  RECT 10.749 0.000 11.089 68.179 ;
 END
 PORT
  LAYER ME4 ;
  RECT 4.743 0.000 5.083 68.179 ;
 END
 PORT
  LAYER ME4 ;
  RECT 5.554 0.000 6.274 31.570 ;
 END
 PORT
  LAYER ME4 ;
  RECT 6.745 0.921 7.085 68.179 ;
 END
 PORT
  LAYER ME4 ;
  RECT 8.747 0.921 9.087 68.179 ;
 END
 PORT
  LAYER ME4 ;
  RECT 17.566 0.000 18.286 31.570 ;
 END
 PORT
  LAYER ME4 ;
  RECT 18.757 0.000 19.097 68.179 ;
 END
 PORT
  LAYER ME4 ;
  RECT 12.751 0.000 13.091 68.179 ;
 END
 PORT
  LAYER ME4 ;
  RECT 13.562 0.000 14.282 31.570 ;
 END
 PORT
  LAYER ME4 ;
  RECT 14.753 0.921 15.093 68.179 ;
 END
 PORT
  LAYER ME4 ;
  RECT 16.755 0.921 17.095 68.179 ;
 END
 PORT
  LAYER ME4 ;
  RECT 25.574 0.000 26.294 31.570 ;
 END
 PORT
  LAYER ME4 ;
  RECT 26.765 0.000 27.105 68.179 ;
 END
 PORT
  LAYER ME4 ;
  RECT 20.759 0.000 21.099 68.179 ;
 END
 PORT
  LAYER ME4 ;
  RECT 21.570 0.000 22.290 31.570 ;
 END
 PORT
  LAYER ME4 ;
  RECT 22.761 0.921 23.101 68.179 ;
 END
 PORT
  LAYER ME4 ;
  RECT 24.763 0.921 25.103 68.179 ;
 END
 PORT
  LAYER ME4 ;
  RECT 33.582 0.000 34.302 31.570 ;
 END
 PORT
  LAYER ME4 ;
  RECT 34.773 0.000 35.113 68.179 ;
 END
 PORT
  LAYER ME4 ;
  RECT 28.767 0.000 29.107 68.179 ;
 END
 PORT
  LAYER ME4 ;
  RECT 29.578 0.000 30.298 31.570 ;
 END
 PORT
  LAYER ME4 ;
  RECT 30.769 0.921 31.109 68.179 ;
 END
 PORT
  LAYER ME4 ;
  RECT 32.771 0.921 33.111 68.179 ;
 END
 PORT
  LAYER ME4 ;
  RECT 41.590 0.000 42.310 31.570 ;
 END
 PORT
  LAYER ME4 ;
  RECT 42.781 0.000 43.121 68.179 ;
 END
 PORT
  LAYER ME4 ;
  RECT 36.775 0.000 37.115 68.179 ;
 END
 PORT
  LAYER ME4 ;
  RECT 37.586 0.000 38.306 31.570 ;
 END
 PORT
  LAYER ME4 ;
  RECT 38.777 0.921 39.117 68.179 ;
 END
 PORT
  LAYER ME4 ;
  RECT 40.779 0.921 41.119 68.179 ;
 END
 PORT
  LAYER ME4 ;
  RECT 49.598 0.000 50.318 31.570 ;
 END
 PORT
  LAYER ME4 ;
  RECT 50.789 0.000 51.129 68.179 ;
 END
 PORT
  LAYER ME4 ;
  RECT 44.783 0.000 45.123 68.179 ;
 END
 PORT
  LAYER ME4 ;
  RECT 45.594 0.000 46.314 31.570 ;
 END
 PORT
  LAYER ME4 ;
  RECT 46.785 0.921 47.125 68.179 ;
 END
 PORT
  LAYER ME4 ;
  RECT 48.787 0.921 49.127 68.179 ;
 END
 PORT
  LAYER ME4 ;
  RECT 57.606 0.000 58.326 31.570 ;
 END
 PORT
  LAYER ME4 ;
  RECT 58.797 0.000 59.137 68.179 ;
 END
 PORT
  LAYER ME4 ;
  RECT 52.791 0.000 53.131 68.179 ;
 END
 PORT
  LAYER ME4 ;
  RECT 53.602 0.000 54.322 31.570 ;
 END
 PORT
  LAYER ME4 ;
  RECT 54.793 0.921 55.133 68.179 ;
 END
 PORT
  LAYER ME4 ;
  RECT 56.795 0.921 57.135 68.179 ;
 END
 PORT
  LAYER ME4 ;
  RECT 65.614 0.000 66.334 31.570 ;
 END
 PORT
  LAYER ME4 ;
  RECT 66.805 0.000 67.145 68.179 ;
 END
 PORT
  LAYER ME4 ;
  RECT 60.799 0.000 61.139 68.179 ;
 END
 PORT
  LAYER ME4 ;
  RECT 61.610 0.000 62.330 31.570 ;
 END
 PORT
  LAYER ME4 ;
  RECT 62.801 0.921 63.141 68.179 ;
 END
 PORT
  LAYER ME4 ;
  RECT 64.803 0.921 65.143 68.179 ;
 END
 PORT
  LAYER ME4 ;
  RECT 69.746 0.000 70.466 68.179 ;
 END
 PORT
  LAYER ME4 ;
  RECT 67.806 0.000 68.146 68.179 ;
 END
END GND
PIN DI7
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 64.662 0.000 64.942 0.720 ;
  LAYER ME3 ;
  RECT 64.662 0.000 64.942 0.720 ;
  LAYER ME2 ;
  RECT 64.662 0.000 64.942 0.720 ;
  LAYER ME1 ;
  RECT 64.662 0.000 64.942 0.720 ;
 END
 ANTENNAPARTIALMETALAREA                  0.805 LAYER ME1 ;
 ANTENNAGATEAREA                          0.072 LAYER ME1 ;
 ANTENNAGATEAREA                          0.072 LAYER ME2 ;
 ANTENNAGATEAREA                          0.072 LAYER ME3 ;
 ANTENNAGATEAREA                          0.072 LAYER ME4 ;
 ANTENNADIFFAREA                          0.218 LAYER ME1 ;
 ANTENNADIFFAREA                          0.218 LAYER ME2 ;
 ANTENNADIFFAREA                          0.218 LAYER ME3 ;
 ANTENNADIFFAREA                          0.218 LAYER ME4 ;
 ANTENNAMAXAREACAR                       13.984 LAYER ME1 ;
 ANTENNAMAXAREACAR                       16.784 LAYER ME2 ;
 ANTENNAMAXAREACAR                       19.584 LAYER ME3 ;
 ANTENNAMAXAREACAR                       22.384 LAYER ME4 ;
END DI7
PIN DO7
  DIRECTION OUTPUT ;
 PORT
  LAYER ME4 ;
  RECT 62.684 0.000 62.964 0.720 ;
  LAYER ME3 ;
  RECT 62.684 0.000 62.964 0.720 ;
  LAYER ME2 ;
  RECT 62.684 0.000 62.964 0.720 ;
  LAYER ME1 ;
  RECT 62.684 0.000 62.964 0.720 ;
 END
 ANTENNAPARTIALMETALAREA                  2.030 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME3 ;
 ANTENNADIFFAREA                          1.293 LAYER ME4 ;
END DO7
PIN DI6
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 56.654 0.000 56.934 0.720 ;
  LAYER ME3 ;
  RECT 56.654 0.000 56.934 0.720 ;
  LAYER ME2 ;
  RECT 56.654 0.000 56.934 0.720 ;
  LAYER ME1 ;
  RECT 56.654 0.000 56.934 0.720 ;
 END
 ANTENNAPARTIALMETALAREA                  0.522 LAYER ME1 ;
 ANTENNAGATEAREA                          0.072 LAYER ME1 ;
 ANTENNAGATEAREA                          0.072 LAYER ME2 ;
 ANTENNAGATEAREA                          0.072 LAYER ME3 ;
 ANTENNAGATEAREA                          0.072 LAYER ME4 ;
 ANTENNADIFFAREA                          0.218 LAYER ME1 ;
 ANTENNADIFFAREA                          0.218 LAYER ME2 ;
 ANTENNADIFFAREA                          0.218 LAYER ME3 ;
 ANTENNADIFFAREA                          0.218 LAYER ME4 ;
 ANTENNAMAXAREACAR                       10.048 LAYER ME1 ;
 ANTENNAMAXAREACAR                       12.848 LAYER ME2 ;
 ANTENNAMAXAREACAR                       15.648 LAYER ME3 ;
 ANTENNAMAXAREACAR                       18.448 LAYER ME4 ;
END DI6
PIN DO6
  DIRECTION OUTPUT ;
 PORT
  LAYER ME4 ;
  RECT 54.596 0.000 54.876 0.720 ;
  LAYER ME3 ;
  RECT 54.596 0.000 54.876 0.720 ;
  LAYER ME2 ;
  RECT 54.596 0.000 54.876 0.720 ;
  LAYER ME1 ;
  RECT 54.596 0.000 54.876 0.720 ;
 END
 ANTENNAPARTIALMETALAREA                  2.030 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME3 ;
 ANTENNADIFFAREA                          1.293 LAYER ME4 ;
END DO6
PIN WEB3
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 55.076 0.000 55.356 0.720 ;
  LAYER ME3 ;
  RECT 55.076 0.000 55.356 0.720 ;
  LAYER ME2 ;
  RECT 55.076 0.000 55.356 0.720 ;
  LAYER ME1 ;
  RECT 55.076 0.000 55.356 0.720 ;
 END
 ANTENNAPARTIALMETALAREA                  0.436 LAYER ME2 ;
 ANTENNAGATEAREA                          0.288 LAYER ME2 ;
 ANTENNAGATEAREA                          0.288 LAYER ME3 ;
 ANTENNAGATEAREA                          0.288 LAYER ME4 ;
 ANTENNADIFFAREA                          0.218 LAYER ME2 ;
 ANTENNADIFFAREA                          0.218 LAYER ME3 ;
 ANTENNADIFFAREA                          0.218 LAYER ME4 ;
 ANTENNAMAXAREACAR                        4.602 LAYER ME2 ;
 ANTENNAMAXAREACAR                        5.302 LAYER ME3 ;
 ANTENNAMAXAREACAR                        6.002 LAYER ME4 ;
END WEB3
PIN DI5
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 48.646 0.000 48.926 0.720 ;
  LAYER ME3 ;
  RECT 48.646 0.000 48.926 0.720 ;
  LAYER ME2 ;
  RECT 48.646 0.000 48.926 0.720 ;
  LAYER ME1 ;
  RECT 48.646 0.000 48.926 0.720 ;
 END
 ANTENNAPARTIALMETALAREA                  0.805 LAYER ME1 ;
 ANTENNAGATEAREA                          0.072 LAYER ME1 ;
 ANTENNAGATEAREA                          0.072 LAYER ME2 ;
 ANTENNAGATEAREA                          0.072 LAYER ME3 ;
 ANTENNAGATEAREA                          0.072 LAYER ME4 ;
 ANTENNADIFFAREA                          0.218 LAYER ME1 ;
 ANTENNADIFFAREA                          0.218 LAYER ME2 ;
 ANTENNADIFFAREA                          0.218 LAYER ME3 ;
 ANTENNADIFFAREA                          0.218 LAYER ME4 ;
 ANTENNAMAXAREACAR                       13.984 LAYER ME1 ;
 ANTENNAMAXAREACAR                       16.784 LAYER ME2 ;
 ANTENNAMAXAREACAR                       19.584 LAYER ME3 ;
 ANTENNAMAXAREACAR                       22.384 LAYER ME4 ;
END DI5
PIN DO5
  DIRECTION OUTPUT ;
 PORT
  LAYER ME4 ;
  RECT 46.668 0.000 46.948 0.720 ;
  LAYER ME3 ;
  RECT 46.668 0.000 46.948 0.720 ;
  LAYER ME2 ;
  RECT 46.668 0.000 46.948 0.720 ;
  LAYER ME1 ;
  RECT 46.668 0.000 46.948 0.720 ;
 END
 ANTENNAPARTIALMETALAREA                  2.030 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME3 ;
 ANTENNADIFFAREA                          1.293 LAYER ME4 ;
END DO5
PIN DI4
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 40.638 0.000 40.918 0.720 ;
  LAYER ME3 ;
  RECT 40.638 0.000 40.918 0.720 ;
  LAYER ME2 ;
  RECT 40.638 0.000 40.918 0.720 ;
  LAYER ME1 ;
  RECT 40.638 0.000 40.918 0.720 ;
 END
 ANTENNAPARTIALMETALAREA                  0.522 LAYER ME1 ;
 ANTENNAGATEAREA                          0.072 LAYER ME1 ;
 ANTENNAGATEAREA                          0.072 LAYER ME2 ;
 ANTENNAGATEAREA                          0.072 LAYER ME3 ;
 ANTENNAGATEAREA                          0.072 LAYER ME4 ;
 ANTENNADIFFAREA                          0.218 LAYER ME1 ;
 ANTENNADIFFAREA                          0.218 LAYER ME2 ;
 ANTENNADIFFAREA                          0.218 LAYER ME3 ;
 ANTENNADIFFAREA                          0.218 LAYER ME4 ;
 ANTENNAMAXAREACAR                       10.048 LAYER ME1 ;
 ANTENNAMAXAREACAR                       12.848 LAYER ME2 ;
 ANTENNAMAXAREACAR                       15.648 LAYER ME3 ;
 ANTENNAMAXAREACAR                       18.448 LAYER ME4 ;
END DI4
PIN DO4
  DIRECTION OUTPUT ;
 PORT
  LAYER ME4 ;
  RECT 38.580 0.000 38.860 0.720 ;
  LAYER ME3 ;
  RECT 38.580 0.000 38.860 0.720 ;
  LAYER ME2 ;
  RECT 38.580 0.000 38.860 0.720 ;
  LAYER ME1 ;
  RECT 38.580 0.000 38.860 0.720 ;
 END
 ANTENNAPARTIALMETALAREA                  2.030 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME3 ;
 ANTENNADIFFAREA                          1.293 LAYER ME4 ;
END DO4
PIN WEB2
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 39.060 0.000 39.340 0.720 ;
  LAYER ME3 ;
  RECT 39.060 0.000 39.340 0.720 ;
  LAYER ME2 ;
  RECT 39.060 0.000 39.340 0.720 ;
  LAYER ME1 ;
  RECT 39.060 0.000 39.340 0.720 ;
 END
 ANTENNAPARTIALMETALAREA                  0.436 LAYER ME2 ;
 ANTENNAGATEAREA                          0.288 LAYER ME2 ;
 ANTENNAGATEAREA                          0.288 LAYER ME3 ;
 ANTENNAGATEAREA                          0.288 LAYER ME4 ;
 ANTENNADIFFAREA                          0.218 LAYER ME2 ;
 ANTENNADIFFAREA                          0.218 LAYER ME3 ;
 ANTENNADIFFAREA                          0.218 LAYER ME4 ;
 ANTENNAMAXAREACAR                        4.602 LAYER ME2 ;
 ANTENNAMAXAREACAR                        5.302 LAYER ME3 ;
 ANTENNAMAXAREACAR                        6.002 LAYER ME4 ;
END WEB2
PIN DI3
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 32.630 0.000 32.910 0.720 ;
  LAYER ME3 ;
  RECT 32.630 0.000 32.910 0.720 ;
  LAYER ME2 ;
  RECT 32.630 0.000 32.910 0.720 ;
  LAYER ME1 ;
  RECT 32.630 0.000 32.910 0.720 ;
 END
 ANTENNAPARTIALMETALAREA                  0.805 LAYER ME1 ;
 ANTENNAGATEAREA                          0.072 LAYER ME1 ;
 ANTENNAGATEAREA                          0.072 LAYER ME2 ;
 ANTENNAGATEAREA                          0.072 LAYER ME3 ;
 ANTENNAGATEAREA                          0.072 LAYER ME4 ;
 ANTENNADIFFAREA                          0.218 LAYER ME1 ;
 ANTENNADIFFAREA                          0.218 LAYER ME2 ;
 ANTENNADIFFAREA                          0.218 LAYER ME3 ;
 ANTENNADIFFAREA                          0.218 LAYER ME4 ;
 ANTENNAMAXAREACAR                       13.984 LAYER ME1 ;
 ANTENNAMAXAREACAR                       16.784 LAYER ME2 ;
 ANTENNAMAXAREACAR                       19.584 LAYER ME3 ;
 ANTENNAMAXAREACAR                       22.384 LAYER ME4 ;
END DI3
PIN DO3
  DIRECTION OUTPUT ;
 PORT
  LAYER ME4 ;
  RECT 30.652 0.000 30.932 0.720 ;
  LAYER ME3 ;
  RECT 30.652 0.000 30.932 0.720 ;
  LAYER ME2 ;
  RECT 30.652 0.000 30.932 0.720 ;
  LAYER ME1 ;
  RECT 30.652 0.000 30.932 0.720 ;
 END
 ANTENNAPARTIALMETALAREA                  2.030 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME3 ;
 ANTENNADIFFAREA                          1.293 LAYER ME4 ;
END DO3
PIN DI2
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 24.622 0.000 24.902 0.720 ;
  LAYER ME3 ;
  RECT 24.622 0.000 24.902 0.720 ;
  LAYER ME2 ;
  RECT 24.622 0.000 24.902 0.720 ;
  LAYER ME1 ;
  RECT 24.622 0.000 24.902 0.720 ;
 END
 ANTENNAPARTIALMETALAREA                  0.522 LAYER ME1 ;
 ANTENNAGATEAREA                          0.072 LAYER ME1 ;
 ANTENNAGATEAREA                          0.072 LAYER ME2 ;
 ANTENNAGATEAREA                          0.072 LAYER ME3 ;
 ANTENNAGATEAREA                          0.072 LAYER ME4 ;
 ANTENNADIFFAREA                          0.218 LAYER ME1 ;
 ANTENNADIFFAREA                          0.218 LAYER ME2 ;
 ANTENNADIFFAREA                          0.218 LAYER ME3 ;
 ANTENNADIFFAREA                          0.218 LAYER ME4 ;
 ANTENNAMAXAREACAR                       10.048 LAYER ME1 ;
 ANTENNAMAXAREACAR                       12.848 LAYER ME2 ;
 ANTENNAMAXAREACAR                       15.648 LAYER ME3 ;
 ANTENNAMAXAREACAR                       18.448 LAYER ME4 ;
END DI2
PIN DO2
  DIRECTION OUTPUT ;
 PORT
  LAYER ME4 ;
  RECT 22.564 0.000 22.844 0.720 ;
  LAYER ME3 ;
  RECT 22.564 0.000 22.844 0.720 ;
  LAYER ME2 ;
  RECT 22.564 0.000 22.844 0.720 ;
  LAYER ME1 ;
  RECT 22.564 0.000 22.844 0.720 ;
 END
 ANTENNAPARTIALMETALAREA                  2.030 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME3 ;
 ANTENNADIFFAREA                          1.293 LAYER ME4 ;
END DO2
PIN WEB1
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 23.044 0.000 23.324 0.720 ;
  LAYER ME3 ;
  RECT 23.044 0.000 23.324 0.720 ;
  LAYER ME2 ;
  RECT 23.044 0.000 23.324 0.720 ;
  LAYER ME1 ;
  RECT 23.044 0.000 23.324 0.720 ;
 END
 ANTENNAPARTIALMETALAREA                  0.436 LAYER ME2 ;
 ANTENNAGATEAREA                          0.288 LAYER ME2 ;
 ANTENNAGATEAREA                          0.288 LAYER ME3 ;
 ANTENNAGATEAREA                          0.288 LAYER ME4 ;
 ANTENNADIFFAREA                          0.218 LAYER ME2 ;
 ANTENNADIFFAREA                          0.218 LAYER ME3 ;
 ANTENNADIFFAREA                          0.218 LAYER ME4 ;
 ANTENNAMAXAREACAR                        4.602 LAYER ME2 ;
 ANTENNAMAXAREACAR                        5.302 LAYER ME3 ;
 ANTENNAMAXAREACAR                        6.002 LAYER ME4 ;
END WEB1
PIN DI1
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 16.614 0.000 16.894 0.720 ;
  LAYER ME3 ;
  RECT 16.614 0.000 16.894 0.720 ;
  LAYER ME2 ;
  RECT 16.614 0.000 16.894 0.720 ;
  LAYER ME1 ;
  RECT 16.614 0.000 16.894 0.720 ;
 END
 ANTENNAPARTIALMETALAREA                  0.805 LAYER ME1 ;
 ANTENNAGATEAREA                          0.072 LAYER ME1 ;
 ANTENNAGATEAREA                          0.072 LAYER ME2 ;
 ANTENNAGATEAREA                          0.072 LAYER ME3 ;
 ANTENNAGATEAREA                          0.072 LAYER ME4 ;
 ANTENNADIFFAREA                          0.218 LAYER ME1 ;
 ANTENNADIFFAREA                          0.218 LAYER ME2 ;
 ANTENNADIFFAREA                          0.218 LAYER ME3 ;
 ANTENNADIFFAREA                          0.218 LAYER ME4 ;
 ANTENNAMAXAREACAR                       13.984 LAYER ME1 ;
 ANTENNAMAXAREACAR                       16.784 LAYER ME2 ;
 ANTENNAMAXAREACAR                       19.584 LAYER ME3 ;
 ANTENNAMAXAREACAR                       22.384 LAYER ME4 ;
END DI1
PIN DO1
  DIRECTION OUTPUT ;
 PORT
  LAYER ME4 ;
  RECT 14.636 0.000 14.916 0.720 ;
  LAYER ME3 ;
  RECT 14.636 0.000 14.916 0.720 ;
  LAYER ME2 ;
  RECT 14.636 0.000 14.916 0.720 ;
  LAYER ME1 ;
  RECT 14.636 0.000 14.916 0.720 ;
 END
 ANTENNAPARTIALMETALAREA                  2.030 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME3 ;
 ANTENNADIFFAREA                          1.293 LAYER ME4 ;
END DO1
PIN DI0
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 8.606 0.000 8.886 0.720 ;
  LAYER ME3 ;
  RECT 8.606 0.000 8.886 0.720 ;
  LAYER ME2 ;
  RECT 8.606 0.000 8.886 0.720 ;
  LAYER ME1 ;
  RECT 8.606 0.000 8.886 0.720 ;
 END
 ANTENNAPARTIALMETALAREA                  0.522 LAYER ME1 ;
 ANTENNAGATEAREA                          0.072 LAYER ME1 ;
 ANTENNAGATEAREA                          0.072 LAYER ME2 ;
 ANTENNAGATEAREA                          0.072 LAYER ME3 ;
 ANTENNAGATEAREA                          0.072 LAYER ME4 ;
 ANTENNADIFFAREA                          0.218 LAYER ME1 ;
 ANTENNADIFFAREA                          0.218 LAYER ME2 ;
 ANTENNADIFFAREA                          0.218 LAYER ME3 ;
 ANTENNADIFFAREA                          0.218 LAYER ME4 ;
 ANTENNAMAXAREACAR                       10.048 LAYER ME1 ;
 ANTENNAMAXAREACAR                       12.848 LAYER ME2 ;
 ANTENNAMAXAREACAR                       15.648 LAYER ME3 ;
 ANTENNAMAXAREACAR                       18.448 LAYER ME4 ;
END DI0
PIN DO0
  DIRECTION OUTPUT ;
 PORT
  LAYER ME4 ;
  RECT 6.548 0.000 6.828 0.720 ;
  LAYER ME3 ;
  RECT 6.548 0.000 6.828 0.720 ;
  LAYER ME2 ;
  RECT 6.548 0.000 6.828 0.720 ;
  LAYER ME1 ;
  RECT 6.548 0.000 6.828 0.720 ;
 END
 ANTENNAPARTIALMETALAREA                  2.030 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME3 ;
 ANTENNADIFFAREA                          1.293 LAYER ME4 ;
END DO0
PIN WEB0
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 7.028 0.000 7.308 0.720 ;
  LAYER ME3 ;
  RECT 7.028 0.000 7.308 0.720 ;
  LAYER ME2 ;
  RECT 7.028 0.000 7.308 0.720 ;
  LAYER ME1 ;
  RECT 7.028 0.000 7.308 0.720 ;
 END
 ANTENNAPARTIALMETALAREA                  0.436 LAYER ME2 ;
 ANTENNAGATEAREA                          0.288 LAYER ME2 ;
 ANTENNAGATEAREA                          0.288 LAYER ME3 ;
 ANTENNAGATEAREA                          0.288 LAYER ME4 ;
 ANTENNADIFFAREA                          0.218 LAYER ME2 ;
 ANTENNADIFFAREA                          0.218 LAYER ME3 ;
 ANTENNADIFFAREA                          0.218 LAYER ME4 ;
 ANTENNAMAXAREACAR                        4.602 LAYER ME2 ;
 ANTENNAMAXAREACAR                        5.302 LAYER ME3 ;
 ANTENNAMAXAREACAR                        6.002 LAYER ME4 ;
END WEB0
PIN A2
  DIRECTION INPUT ;
 PORT
  LAYER ME3 ;
  RECT 82.948 0.000 83.268 0.600 ;
  LAYER ME2 ;
  RECT 82.948 0.000 83.268 0.600 ;
  LAYER ME1 ;
  RECT 82.948 0.000 83.268 0.600 ;
 END
 ANTENNAPARTIALMETALAREA                  1.067 LAYER ME2 ;
 ANTENNAGATEAREA                          0.144 LAYER ME2 ;
 ANTENNAGATEAREA                          0.144 LAYER ME3 ;
 ANTENNADIFFAREA                          0.218 LAYER ME2 ;
 ANTENNADIFFAREA                          0.218 LAYER ME3 ;
 ANTENNAMAXAREACAR                        9.746 LAYER ME2 ;
 ANTENNAMAXAREACAR                       11.079 LAYER ME3 ;
END A2
PIN A3
  DIRECTION INPUT ;
 PORT
  LAYER ME3 ;
  RECT 83.535 0.000 83.855 0.600 ;
  LAYER ME2 ;
  RECT 83.535 0.000 83.855 0.600 ;
  LAYER ME1 ;
  RECT 83.535 0.000 83.855 0.600 ;
 END
 ANTENNAPARTIALMETALAREA                  1.188 LAYER ME2 ;
 ANTENNAGATEAREA                          0.144 LAYER ME2 ;
 ANTENNAGATEAREA                          0.144 LAYER ME3 ;
 ANTENNADIFFAREA                          0.218 LAYER ME2 ;
 ANTENNADIFFAREA                          0.218 LAYER ME3 ;
 ANTENNAMAXAREACAR                       10.582 LAYER ME2 ;
 ANTENNAMAXAREACAR                       11.915 LAYER ME3 ;
END A3
PIN A4
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 76.696 0.000 77.016 0.600 ;
  LAYER ME3 ;
  RECT 76.696 0.000 77.016 0.600 ;
  LAYER ME2 ;
  RECT 76.696 0.000 77.016 0.600 ;
  LAYER ME1 ;
  RECT 76.696 0.000 77.016 0.600 ;
 END
 ANTENNAPARTIALMETALAREA                  1.910 LAYER ME2 ;
 ANTENNAGATEAREA                          0.180 LAYER ME2 ;
 ANTENNAGATEAREA                          0.180 LAYER ME3 ;
 ANTENNAGATEAREA                          0.180 LAYER ME4 ;
 ANTENNADIFFAREA                          0.218 LAYER ME2 ;
 ANTENNADIFFAREA                          0.218 LAYER ME3 ;
 ANTENNADIFFAREA                          0.218 LAYER ME4 ;
 ANTENNAMAXAREACAR                       13.456 LAYER ME2 ;
 ANTENNAMAXAREACAR                       14.522 LAYER ME3 ;
 ANTENNAMAXAREACAR                       15.589 LAYER ME4 ;
END A4
PIN A5
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 76.076 0.000 76.396 0.600 ;
  LAYER ME3 ;
  RECT 76.076 0.000 76.396 0.600 ;
  LAYER ME2 ;
  RECT 76.076 0.000 76.396 0.600 ;
  LAYER ME1 ;
  RECT 76.076 0.000 76.396 0.600 ;
 END
 ANTENNAPARTIALMETALAREA                  1.447 LAYER ME2 ;
 ANTENNAGATEAREA                          0.180 LAYER ME2 ;
 ANTENNAGATEAREA                          0.180 LAYER ME3 ;
 ANTENNAGATEAREA                          0.180 LAYER ME4 ;
 ANTENNADIFFAREA                          0.218 LAYER ME2 ;
 ANTENNADIFFAREA                          0.218 LAYER ME3 ;
 ANTENNADIFFAREA                          0.218 LAYER ME4 ;
 ANTENNAMAXAREACAR                       12.818 LAYER ME2 ;
 ANTENNAMAXAREACAR                       13.884 LAYER ME3 ;
 ANTENNAMAXAREACAR                       14.951 LAYER ME4 ;
END A5
PIN A6
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 72.596 0.000 72.916 0.600 ;
  LAYER ME3 ;
  RECT 72.596 0.000 72.916 0.600 ;
  LAYER ME2 ;
  RECT 72.596 0.000 72.916 0.600 ;
  LAYER ME1 ;
  RECT 72.596 0.000 72.916 0.600 ;
 END
 ANTENNAPARTIALMETALAREA                  1.910 LAYER ME2 ;
 ANTENNAGATEAREA                          0.180 LAYER ME2 ;
 ANTENNAGATEAREA                          0.180 LAYER ME3 ;
 ANTENNAGATEAREA                          0.180 LAYER ME4 ;
 ANTENNADIFFAREA                          0.218 LAYER ME2 ;
 ANTENNADIFFAREA                          0.218 LAYER ME3 ;
 ANTENNADIFFAREA                          0.218 LAYER ME4 ;
 ANTENNAMAXAREACAR                       13.456 LAYER ME2 ;
 ANTENNAMAXAREACAR                       14.522 LAYER ME3 ;
 ANTENNAMAXAREACAR                       15.589 LAYER ME4 ;
END A6
PIN A1
  DIRECTION INPUT ;
 PORT
  LAYER ME3 ;
  RECT 87.821 0.000 88.141 0.712 ;
  LAYER ME2 ;
  RECT 87.821 0.000 88.141 0.712 ;
  LAYER ME1 ;
  RECT 87.821 0.000 88.141 0.712 ;
 END
 ANTENNAPARTIALMETALAREA                  3.219 LAYER ME2 ;
 ANTENNAGATEAREA                          0.108 LAYER ME2 ;
 ANTENNAGATEAREA                          0.108 LAYER ME3 ;
 ANTENNADIFFAREA                          0.218 LAYER ME2 ;
 ANTENNADIFFAREA                          0.218 LAYER ME3 ;
 ANTENNAMAXAREACAR                       33.245 LAYER ME2 ;
 ANTENNAMAXAREACAR                       35.355 LAYER ME3 ;
END A1
PIN A0
  DIRECTION INPUT ;
 PORT
  LAYER ME3 ;
  RECT 91.050 0.000 91.370 0.712 ;
  LAYER ME2 ;
  RECT 91.050 0.000 91.370 0.712 ;
  LAYER ME1 ;
  RECT 91.050 0.000 91.370 0.712 ;
 END
 ANTENNAPARTIALMETALAREA                  3.457 LAYER ME2 ;
 ANTENNAGATEAREA                          0.108 LAYER ME2 ;
 ANTENNAGATEAREA                          0.108 LAYER ME3 ;
 ANTENNADIFFAREA                          0.218 LAYER ME2 ;
 ANTENNADIFFAREA                          0.218 LAYER ME3 ;
 ANTENNAMAXAREACAR                       35.986 LAYER ME2 ;
 ANTENNAMAXAREACAR                       38.095 LAYER ME3 ;
END A0
PIN DVSE
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 103.641 0.000 103.961 0.717 ;
  LAYER ME3 ;
  RECT 103.641 0.000 103.961 0.717 ;
  LAYER ME3 ;
  RECT 103.641 0.000 103.961 0.717 ;
  LAYER ME2 ;
  RECT 103.641 0.000 103.961 0.717 ;
  LAYER ME2 ;
  RECT 103.641 0.000 103.961 0.717 ;
  LAYER ME1 ;
  RECT 103.641 0.000 103.961 0.717 ;
  LAYER ME1 ;
  RECT 103.641 0.000 103.961 0.717 ;
 END
 ANTENNAPARTIALMETALAREA                  5.305 LAYER ME2 ;
 ANTENNAGATEAREA                          0.612 LAYER ME2 ;
 ANTENNAGATEAREA                          0.612 LAYER ME3 ;
 ANTENNAGATEAREA                          0.612 LAYER ME4 ;
 ANTENNADIFFAREA                          0.218 LAYER ME2 ;
 ANTENNADIFFAREA                          0.218 LAYER ME3 ;
 ANTENNADIFFAREA                          0.218 LAYER ME4 ;
 ANTENNAMAXAREACAR                       53.132 LAYER ME2 ;
 ANTENNAMAXAREACAR                       55.256 LAYER ME3 ;
 ANTENNAMAXAREACAR                       57.381 LAYER ME4 ;
END DVSE
PIN DVS3
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 103.121 0.000 103.441 0.717 ;
  LAYER ME3 ;
  RECT 103.121 0.000 103.441 0.717 ;
  LAYER ME3 ;
  RECT 103.121 0.000 103.441 0.717 ;
  LAYER ME2 ;
  RECT 103.121 0.000 103.441 0.717 ;
  LAYER ME2 ;
  RECT 103.121 0.000 103.441 0.717 ;
  LAYER ME1 ;
  RECT 103.121 0.000 103.441 0.717 ;
  LAYER ME1 ;
  RECT 103.121 0.000 103.441 0.717 ;
 END
 ANTENNAPARTIALMETALAREA                  3.675 LAYER ME2 ;
 ANTENNAGATEAREA                          0.108 LAYER ME2 ;
 ANTENNAGATEAREA                          0.108 LAYER ME3 ;
 ANTENNAGATEAREA                          0.108 LAYER ME4 ;
 ANTENNADIFFAREA                          0.218 LAYER ME2 ;
 ANTENNADIFFAREA                          0.218 LAYER ME3 ;
 ANTENNADIFFAREA                          0.218 LAYER ME4 ;
 ANTENNAMAXAREACAR                       45.625 LAYER ME2 ;
 ANTENNAMAXAREACAR                       47.749 LAYER ME3 ;
 ANTENNAMAXAREACAR                       49.874 LAYER ME4 ;
END DVS3
PIN DVS2
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 104.161 0.000 104.481 0.717 ;
  LAYER ME3 ;
  RECT 104.161 0.000 104.481 0.717 ;
  LAYER ME3 ;
  RECT 104.161 0.000 104.481 0.717 ;
  LAYER ME2 ;
  RECT 104.161 0.000 104.481 0.717 ;
  LAYER ME2 ;
  RECT 104.161 0.000 104.481 0.717 ;
  LAYER ME1 ;
  RECT 104.161 0.000 104.481 0.717 ;
  LAYER ME1 ;
  RECT 104.161 0.000 104.481 0.717 ;
 END
 ANTENNAPARTIALMETALAREA                  5.371 LAYER ME2 ;
 ANTENNAGATEAREA                          0.108 LAYER ME2 ;
 ANTENNAGATEAREA                          0.108 LAYER ME3 ;
 ANTENNAGATEAREA                          0.108 LAYER ME4 ;
 ANTENNADIFFAREA                          0.218 LAYER ME2 ;
 ANTENNADIFFAREA                          0.218 LAYER ME3 ;
 ANTENNADIFFAREA                          0.218 LAYER ME4 ;
 ANTENNAMAXAREACAR                       60.060 LAYER ME2 ;
 ANTENNAMAXAREACAR                       62.184 LAYER ME3 ;
 ANTENNAMAXAREACAR                       64.309 LAYER ME4 ;
END DVS2
PIN DVS1
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 102.601 0.000 102.921 0.717 ;
  LAYER ME3 ;
  RECT 102.601 0.000 102.921 0.717 ;
  LAYER ME3 ;
  RECT 102.601 0.000 102.921 0.717 ;
  LAYER ME2 ;
  RECT 102.601 0.000 102.921 0.717 ;
  LAYER ME2 ;
  RECT 102.601 0.000 102.921 0.717 ;
  LAYER ME1 ;
  RECT 102.601 0.000 102.921 0.717 ;
  LAYER ME1 ;
  RECT 102.601 0.000 102.921 0.717 ;
 END
 ANTENNAPARTIALMETALAREA                  3.307 LAYER ME2 ;
 ANTENNAGATEAREA                          0.108 LAYER ME2 ;
 ANTENNAGATEAREA                          0.108 LAYER ME3 ;
 ANTENNAGATEAREA                          0.108 LAYER ME4 ;
 ANTENNADIFFAREA                          0.218 LAYER ME2 ;
 ANTENNADIFFAREA                          0.218 LAYER ME3 ;
 ANTENNADIFFAREA                          0.218 LAYER ME4 ;
 ANTENNAMAXAREACAR                       42.063 LAYER ME2 ;
 ANTENNAMAXAREACAR                       44.188 LAYER ME3 ;
 ANTENNAMAXAREACAR                       46.312 LAYER ME4 ;
END DVS1
PIN DVS0
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 104.681 0.000 105.001 0.693 ;
  LAYER ME3 ;
  RECT 104.681 0.000 105.001 0.693 ;
  LAYER ME3 ;
  RECT 104.681 0.000 105.001 0.693 ;
  LAYER ME2 ;
  RECT 104.681 0.000 105.001 0.693 ;
  LAYER ME2 ;
  RECT 104.681 0.000 105.001 0.693 ;
  LAYER ME1 ;
  RECT 104.681 0.000 105.001 0.693 ;
  LAYER ME1 ;
  RECT 104.681 0.000 105.001 0.693 ;
 END
 ANTENNAPARTIALMETALAREA                  4.376 LAYER ME2 ;
 ANTENNAGATEAREA                          0.108 LAYER ME2 ;
 ANTENNAGATEAREA                          0.108 LAYER ME3 ;
 ANTENNAGATEAREA                          0.108 LAYER ME4 ;
 ANTENNADIFFAREA                          0.218 LAYER ME2 ;
 ANTENNADIFFAREA                          0.218 LAYER ME3 ;
 ANTENNADIFFAREA                          0.218 LAYER ME4 ;
 ANTENNAMAXAREACAR                       53.260 LAYER ME2 ;
 ANTENNAMAXAREACAR                       55.313 LAYER ME3 ;
 ANTENNAMAXAREACAR                       57.367 LAYER ME4 ;
END DVS0
PIN CK
  DIRECTION INPUT ;
 PORT
  LAYER ME3 ;
  RECT 96.117 0.000 96.437 0.713 ;
  LAYER ME2 ;
  RECT 96.117 0.000 96.437 0.713 ;
  LAYER ME1 ;
  RECT 96.117 0.000 96.437 0.713 ;
 END
 ANTENNAPARTIALMETALAREA                  2.392 LAYER ME2 ;
 ANTENNAPARTIALMETALAREA                  7.363 LAYER ME3 ;
 ANTENNAGATEAREA                          0.072 LAYER ME2 ;
 ANTENNAGATEAREA                          1.260 LAYER ME3 ;
 ANTENNADIFFAREA                          0.218 LAYER ME2 ;
 ANTENNADIFFAREA                          0.218 LAYER ME3 ;
 ANTENNAMAXAREACAR                       46.148 LAYER ME2 ;
 ANTENNAMAXAREACAR                      151.587 LAYER ME3 ;
END CK
PIN CSB
  DIRECTION INPUT ;
 PORT
  LAYER ME3 ;
  RECT 89.329 0.000 89.649 0.712 ;
  LAYER ME2 ;
  RECT 89.329 0.000 89.649 0.712 ;
  LAYER ME1 ;
  RECT 89.329 0.000 89.649 0.712 ;
 END
 ANTENNAPARTIALMETALAREA                  3.350 LAYER ME2 ;
 ANTENNAPARTIALMETALAREA                  7.235 LAYER ME3 ;
 ANTENNAGATEAREA                          2.244 LAYER ME2 ;
 ANTENNAGATEAREA                          3.216 LAYER ME3 ;
 ANTENNADIFFAREA                          0.218 LAYER ME2 ;
 ANTENNADIFFAREA                          0.218 LAYER ME3 ;
 ANTENNAMAXAREACAR                       17.231 LAYER ME2 ;
 ANTENNAMAXAREACAR                       51.784 LAYER ME3 ;
END CSB
PIN DI15
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 166.403 0.000 166.683 0.720 ;
  LAYER ME3 ;
  RECT 166.403 0.000 166.683 0.720 ;
  LAYER ME2 ;
  RECT 166.403 0.000 166.683 0.720 ;
  LAYER ME1 ;
  RECT 166.403 0.000 166.683 0.720 ;
 END
 ANTENNAPARTIALMETALAREA                  0.805 LAYER ME1 ;
 ANTENNAGATEAREA                          0.072 LAYER ME1 ;
 ANTENNAGATEAREA                          0.072 LAYER ME2 ;
 ANTENNAGATEAREA                          0.072 LAYER ME3 ;
 ANTENNAGATEAREA                          0.072 LAYER ME4 ;
 ANTENNADIFFAREA                          0.218 LAYER ME1 ;
 ANTENNADIFFAREA                          0.218 LAYER ME2 ;
 ANTENNADIFFAREA                          0.218 LAYER ME3 ;
 ANTENNADIFFAREA                          0.218 LAYER ME4 ;
 ANTENNAMAXAREACAR                       13.984 LAYER ME1 ;
 ANTENNAMAXAREACAR                       16.784 LAYER ME2 ;
 ANTENNAMAXAREACAR                       19.584 LAYER ME3 ;
 ANTENNAMAXAREACAR                       22.384 LAYER ME4 ;
END DI15
PIN DO15
  DIRECTION OUTPUT ;
 PORT
  LAYER ME4 ;
  RECT 164.425 0.000 164.705 0.720 ;
  LAYER ME3 ;
  RECT 164.425 0.000 164.705 0.720 ;
  LAYER ME2 ;
  RECT 164.425 0.000 164.705 0.720 ;
  LAYER ME1 ;
  RECT 164.425 0.000 164.705 0.720 ;
 END
 ANTENNAPARTIALMETALAREA                  2.030 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME3 ;
 ANTENNADIFFAREA                          1.293 LAYER ME4 ;
END DO15
PIN DI14
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 158.395 0.000 158.675 0.720 ;
  LAYER ME3 ;
  RECT 158.395 0.000 158.675 0.720 ;
  LAYER ME2 ;
  RECT 158.395 0.000 158.675 0.720 ;
  LAYER ME1 ;
  RECT 158.395 0.000 158.675 0.720 ;
 END
 ANTENNAPARTIALMETALAREA                  0.522 LAYER ME1 ;
 ANTENNAGATEAREA                          0.072 LAYER ME1 ;
 ANTENNAGATEAREA                          0.072 LAYER ME2 ;
 ANTENNAGATEAREA                          0.072 LAYER ME3 ;
 ANTENNAGATEAREA                          0.072 LAYER ME4 ;
 ANTENNADIFFAREA                          0.218 LAYER ME1 ;
 ANTENNADIFFAREA                          0.218 LAYER ME2 ;
 ANTENNADIFFAREA                          0.218 LAYER ME3 ;
 ANTENNADIFFAREA                          0.218 LAYER ME4 ;
 ANTENNAMAXAREACAR                       10.048 LAYER ME1 ;
 ANTENNAMAXAREACAR                       12.848 LAYER ME2 ;
 ANTENNAMAXAREACAR                       15.648 LAYER ME3 ;
 ANTENNAMAXAREACAR                       18.448 LAYER ME4 ;
END DI14
PIN DO14
  DIRECTION OUTPUT ;
 PORT
  LAYER ME4 ;
  RECT 156.337 0.000 156.617 0.720 ;
  LAYER ME3 ;
  RECT 156.337 0.000 156.617 0.720 ;
  LAYER ME2 ;
  RECT 156.337 0.000 156.617 0.720 ;
  LAYER ME1 ;
  RECT 156.337 0.000 156.617 0.720 ;
 END
 ANTENNAPARTIALMETALAREA                  2.030 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME3 ;
 ANTENNADIFFAREA                          1.293 LAYER ME4 ;
END DO14
PIN WEB7
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 156.817 0.000 157.097 0.720 ;
  LAYER ME3 ;
  RECT 156.817 0.000 157.097 0.720 ;
  LAYER ME2 ;
  RECT 156.817 0.000 157.097 0.720 ;
  LAYER ME1 ;
  RECT 156.817 0.000 157.097 0.720 ;
 END
 ANTENNAPARTIALMETALAREA                  0.436 LAYER ME2 ;
 ANTENNAGATEAREA                          0.288 LAYER ME2 ;
 ANTENNAGATEAREA                          0.288 LAYER ME3 ;
 ANTENNAGATEAREA                          0.288 LAYER ME4 ;
 ANTENNADIFFAREA                          0.218 LAYER ME2 ;
 ANTENNADIFFAREA                          0.218 LAYER ME3 ;
 ANTENNADIFFAREA                          0.218 LAYER ME4 ;
 ANTENNAMAXAREACAR                        4.602 LAYER ME2 ;
 ANTENNAMAXAREACAR                        5.302 LAYER ME3 ;
 ANTENNAMAXAREACAR                        6.002 LAYER ME4 ;
END WEB7
PIN DI13
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 150.387 0.000 150.667 0.720 ;
  LAYER ME3 ;
  RECT 150.387 0.000 150.667 0.720 ;
  LAYER ME2 ;
  RECT 150.387 0.000 150.667 0.720 ;
  LAYER ME1 ;
  RECT 150.387 0.000 150.667 0.720 ;
 END
 ANTENNAPARTIALMETALAREA                  0.805 LAYER ME1 ;
 ANTENNAGATEAREA                          0.072 LAYER ME1 ;
 ANTENNAGATEAREA                          0.072 LAYER ME2 ;
 ANTENNAGATEAREA                          0.072 LAYER ME3 ;
 ANTENNAGATEAREA                          0.072 LAYER ME4 ;
 ANTENNADIFFAREA                          0.218 LAYER ME1 ;
 ANTENNADIFFAREA                          0.218 LAYER ME2 ;
 ANTENNADIFFAREA                          0.218 LAYER ME3 ;
 ANTENNADIFFAREA                          0.218 LAYER ME4 ;
 ANTENNAMAXAREACAR                       13.984 LAYER ME1 ;
 ANTENNAMAXAREACAR                       16.784 LAYER ME2 ;
 ANTENNAMAXAREACAR                       19.584 LAYER ME3 ;
 ANTENNAMAXAREACAR                       22.384 LAYER ME4 ;
END DI13
PIN DO13
  DIRECTION OUTPUT ;
 PORT
  LAYER ME4 ;
  RECT 148.409 0.000 148.689 0.720 ;
  LAYER ME3 ;
  RECT 148.409 0.000 148.689 0.720 ;
  LAYER ME2 ;
  RECT 148.409 0.000 148.689 0.720 ;
  LAYER ME1 ;
  RECT 148.409 0.000 148.689 0.720 ;
 END
 ANTENNAPARTIALMETALAREA                  2.030 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME3 ;
 ANTENNADIFFAREA                          1.293 LAYER ME4 ;
END DO13
PIN DI12
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 142.379 0.000 142.659 0.720 ;
  LAYER ME3 ;
  RECT 142.379 0.000 142.659 0.720 ;
  LAYER ME2 ;
  RECT 142.379 0.000 142.659 0.720 ;
  LAYER ME1 ;
  RECT 142.379 0.000 142.659 0.720 ;
 END
 ANTENNAPARTIALMETALAREA                  0.522 LAYER ME1 ;
 ANTENNAGATEAREA                          0.072 LAYER ME1 ;
 ANTENNAGATEAREA                          0.072 LAYER ME2 ;
 ANTENNAGATEAREA                          0.072 LAYER ME3 ;
 ANTENNAGATEAREA                          0.072 LAYER ME4 ;
 ANTENNADIFFAREA                          0.218 LAYER ME1 ;
 ANTENNADIFFAREA                          0.218 LAYER ME2 ;
 ANTENNADIFFAREA                          0.218 LAYER ME3 ;
 ANTENNADIFFAREA                          0.218 LAYER ME4 ;
 ANTENNAMAXAREACAR                       10.048 LAYER ME1 ;
 ANTENNAMAXAREACAR                       12.848 LAYER ME2 ;
 ANTENNAMAXAREACAR                       15.648 LAYER ME3 ;
 ANTENNAMAXAREACAR                       18.448 LAYER ME4 ;
END DI12
PIN DO12
  DIRECTION OUTPUT ;
 PORT
  LAYER ME4 ;
  RECT 140.321 0.000 140.601 0.720 ;
  LAYER ME3 ;
  RECT 140.321 0.000 140.601 0.720 ;
  LAYER ME2 ;
  RECT 140.321 0.000 140.601 0.720 ;
  LAYER ME1 ;
  RECT 140.321 0.000 140.601 0.720 ;
 END
 ANTENNAPARTIALMETALAREA                  2.030 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME3 ;
 ANTENNADIFFAREA                          1.293 LAYER ME4 ;
END DO12
PIN WEB6
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 140.801 0.000 141.081 0.720 ;
  LAYER ME3 ;
  RECT 140.801 0.000 141.081 0.720 ;
  LAYER ME2 ;
  RECT 140.801 0.000 141.081 0.720 ;
  LAYER ME1 ;
  RECT 140.801 0.000 141.081 0.720 ;
 END
 ANTENNAPARTIALMETALAREA                  0.436 LAYER ME2 ;
 ANTENNAGATEAREA                          0.288 LAYER ME2 ;
 ANTENNAGATEAREA                          0.288 LAYER ME3 ;
 ANTENNAGATEAREA                          0.288 LAYER ME4 ;
 ANTENNADIFFAREA                          0.218 LAYER ME2 ;
 ANTENNADIFFAREA                          0.218 LAYER ME3 ;
 ANTENNADIFFAREA                          0.218 LAYER ME4 ;
 ANTENNAMAXAREACAR                        4.602 LAYER ME2 ;
 ANTENNAMAXAREACAR                        5.302 LAYER ME3 ;
 ANTENNAMAXAREACAR                        6.002 LAYER ME4 ;
END WEB6
PIN DI11
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 134.371 0.000 134.651 0.720 ;
  LAYER ME3 ;
  RECT 134.371 0.000 134.651 0.720 ;
  LAYER ME2 ;
  RECT 134.371 0.000 134.651 0.720 ;
  LAYER ME1 ;
  RECT 134.371 0.000 134.651 0.720 ;
 END
 ANTENNAPARTIALMETALAREA                  0.805 LAYER ME1 ;
 ANTENNAGATEAREA                          0.072 LAYER ME1 ;
 ANTENNAGATEAREA                          0.072 LAYER ME2 ;
 ANTENNAGATEAREA                          0.072 LAYER ME3 ;
 ANTENNAGATEAREA                          0.072 LAYER ME4 ;
 ANTENNADIFFAREA                          0.218 LAYER ME1 ;
 ANTENNADIFFAREA                          0.218 LAYER ME2 ;
 ANTENNADIFFAREA                          0.218 LAYER ME3 ;
 ANTENNADIFFAREA                          0.218 LAYER ME4 ;
 ANTENNAMAXAREACAR                       13.984 LAYER ME1 ;
 ANTENNAMAXAREACAR                       16.784 LAYER ME2 ;
 ANTENNAMAXAREACAR                       19.584 LAYER ME3 ;
 ANTENNAMAXAREACAR                       22.384 LAYER ME4 ;
END DI11
PIN DO11
  DIRECTION OUTPUT ;
 PORT
  LAYER ME4 ;
  RECT 132.393 0.000 132.673 0.720 ;
  LAYER ME3 ;
  RECT 132.393 0.000 132.673 0.720 ;
  LAYER ME2 ;
  RECT 132.393 0.000 132.673 0.720 ;
  LAYER ME1 ;
  RECT 132.393 0.000 132.673 0.720 ;
 END
 ANTENNAPARTIALMETALAREA                  2.030 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME3 ;
 ANTENNADIFFAREA                          1.293 LAYER ME4 ;
END DO11
PIN DI10
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 126.363 0.000 126.643 0.720 ;
  LAYER ME3 ;
  RECT 126.363 0.000 126.643 0.720 ;
  LAYER ME2 ;
  RECT 126.363 0.000 126.643 0.720 ;
  LAYER ME1 ;
  RECT 126.363 0.000 126.643 0.720 ;
 END
 ANTENNAPARTIALMETALAREA                  0.522 LAYER ME1 ;
 ANTENNAGATEAREA                          0.072 LAYER ME1 ;
 ANTENNAGATEAREA                          0.072 LAYER ME2 ;
 ANTENNAGATEAREA                          0.072 LAYER ME3 ;
 ANTENNAGATEAREA                          0.072 LAYER ME4 ;
 ANTENNADIFFAREA                          0.218 LAYER ME1 ;
 ANTENNADIFFAREA                          0.218 LAYER ME2 ;
 ANTENNADIFFAREA                          0.218 LAYER ME3 ;
 ANTENNADIFFAREA                          0.218 LAYER ME4 ;
 ANTENNAMAXAREACAR                       10.048 LAYER ME1 ;
 ANTENNAMAXAREACAR                       12.848 LAYER ME2 ;
 ANTENNAMAXAREACAR                       15.648 LAYER ME3 ;
 ANTENNAMAXAREACAR                       18.448 LAYER ME4 ;
END DI10
PIN DO10
  DIRECTION OUTPUT ;
 PORT
  LAYER ME4 ;
  RECT 124.305 0.000 124.585 0.720 ;
  LAYER ME3 ;
  RECT 124.305 0.000 124.585 0.720 ;
  LAYER ME2 ;
  RECT 124.305 0.000 124.585 0.720 ;
  LAYER ME1 ;
  RECT 124.305 0.000 124.585 0.720 ;
 END
 ANTENNAPARTIALMETALAREA                  2.030 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME3 ;
 ANTENNADIFFAREA                          1.293 LAYER ME4 ;
END DO10
PIN WEB5
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 124.785 0.000 125.065 0.720 ;
  LAYER ME3 ;
  RECT 124.785 0.000 125.065 0.720 ;
  LAYER ME2 ;
  RECT 124.785 0.000 125.065 0.720 ;
  LAYER ME1 ;
  RECT 124.785 0.000 125.065 0.720 ;
 END
 ANTENNAPARTIALMETALAREA                  0.436 LAYER ME2 ;
 ANTENNAGATEAREA                          0.288 LAYER ME2 ;
 ANTENNAGATEAREA                          0.288 LAYER ME3 ;
 ANTENNAGATEAREA                          0.288 LAYER ME4 ;
 ANTENNADIFFAREA                          0.218 LAYER ME2 ;
 ANTENNADIFFAREA                          0.218 LAYER ME3 ;
 ANTENNADIFFAREA                          0.218 LAYER ME4 ;
 ANTENNAMAXAREACAR                        4.602 LAYER ME2 ;
 ANTENNAMAXAREACAR                        5.302 LAYER ME3 ;
 ANTENNAMAXAREACAR                        6.002 LAYER ME4 ;
END WEB5
PIN DI9
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 118.355 0.000 118.635 0.720 ;
  LAYER ME3 ;
  RECT 118.355 0.000 118.635 0.720 ;
  LAYER ME2 ;
  RECT 118.355 0.000 118.635 0.720 ;
  LAYER ME1 ;
  RECT 118.355 0.000 118.635 0.720 ;
 END
 ANTENNAPARTIALMETALAREA                  0.805 LAYER ME1 ;
 ANTENNAGATEAREA                          0.072 LAYER ME1 ;
 ANTENNAGATEAREA                          0.072 LAYER ME2 ;
 ANTENNAGATEAREA                          0.072 LAYER ME3 ;
 ANTENNAGATEAREA                          0.072 LAYER ME4 ;
 ANTENNADIFFAREA                          0.218 LAYER ME1 ;
 ANTENNADIFFAREA                          0.218 LAYER ME2 ;
 ANTENNADIFFAREA                          0.218 LAYER ME3 ;
 ANTENNADIFFAREA                          0.218 LAYER ME4 ;
 ANTENNAMAXAREACAR                       13.984 LAYER ME1 ;
 ANTENNAMAXAREACAR                       16.784 LAYER ME2 ;
 ANTENNAMAXAREACAR                       19.584 LAYER ME3 ;
 ANTENNAMAXAREACAR                       22.384 LAYER ME4 ;
END DI9
PIN DO9
  DIRECTION OUTPUT ;
 PORT
  LAYER ME4 ;
  RECT 116.377 0.000 116.657 0.720 ;
  LAYER ME3 ;
  RECT 116.377 0.000 116.657 0.720 ;
  LAYER ME2 ;
  RECT 116.377 0.000 116.657 0.720 ;
  LAYER ME1 ;
  RECT 116.377 0.000 116.657 0.720 ;
 END
 ANTENNAPARTIALMETALAREA                  2.030 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME3 ;
 ANTENNADIFFAREA                          1.293 LAYER ME4 ;
END DO9
PIN DI8
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 110.347 0.000 110.627 0.720 ;
  LAYER ME3 ;
  RECT 110.347 0.000 110.627 0.720 ;
  LAYER ME2 ;
  RECT 110.347 0.000 110.627 0.720 ;
  LAYER ME1 ;
  RECT 110.347 0.000 110.627 0.720 ;
 END
 ANTENNAPARTIALMETALAREA                  0.522 LAYER ME1 ;
 ANTENNAGATEAREA                          0.072 LAYER ME1 ;
 ANTENNAGATEAREA                          0.072 LAYER ME2 ;
 ANTENNAGATEAREA                          0.072 LAYER ME3 ;
 ANTENNAGATEAREA                          0.072 LAYER ME4 ;
 ANTENNADIFFAREA                          0.218 LAYER ME1 ;
 ANTENNADIFFAREA                          0.218 LAYER ME2 ;
 ANTENNADIFFAREA                          0.218 LAYER ME3 ;
 ANTENNADIFFAREA                          0.218 LAYER ME4 ;
 ANTENNAMAXAREACAR                       10.048 LAYER ME1 ;
 ANTENNAMAXAREACAR                       12.848 LAYER ME2 ;
 ANTENNAMAXAREACAR                       15.648 LAYER ME3 ;
 ANTENNAMAXAREACAR                       18.448 LAYER ME4 ;
END DI8
PIN DO8
  DIRECTION OUTPUT ;
 PORT
  LAYER ME4 ;
  RECT 108.289 0.000 108.569 0.720 ;
  LAYER ME3 ;
  RECT 108.289 0.000 108.569 0.720 ;
  LAYER ME2 ;
  RECT 108.289 0.000 108.569 0.720 ;
  LAYER ME1 ;
  RECT 108.289 0.000 108.569 0.720 ;
 END
 ANTENNAPARTIALMETALAREA                  2.030 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME2 ;
 ANTENNADIFFAREA                          1.293 LAYER ME3 ;
 ANTENNADIFFAREA                          1.293 LAYER ME4 ;
END DO8
PIN WEB4
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 108.769 0.000 109.049 0.720 ;
  LAYER ME3 ;
  RECT 108.769 0.000 109.049 0.720 ;
  LAYER ME2 ;
  RECT 108.769 0.000 109.049 0.720 ;
  LAYER ME1 ;
  RECT 108.769 0.000 109.049 0.720 ;
 END
 ANTENNAPARTIALMETALAREA                  0.436 LAYER ME2 ;
 ANTENNAGATEAREA                          0.288 LAYER ME2 ;
 ANTENNAGATEAREA                          0.288 LAYER ME3 ;
 ANTENNAGATEAREA                          0.288 LAYER ME4 ;
 ANTENNADIFFAREA                          0.218 LAYER ME2 ;
 ANTENNADIFFAREA                          0.218 LAYER ME3 ;
 ANTENNADIFFAREA                          0.218 LAYER ME4 ;
 ANTENNAMAXAREACAR                        4.602 LAYER ME2 ;
 ANTENNAMAXAREACAR                        5.302 LAYER ME3 ;
 ANTENNAMAXAREACAR                        6.002 LAYER ME4 ;
END WEB4
OBS
  LAYER ME3 ;
  RECT 0.000 0.000 171.627 68.179 ;
  LAYER ME2 ;
  RECT 0.000 0.000 171.627 68.179 ;
  LAYER ME1 ;
  RECT 0.000 0.000 171.627 68.179 ;
  LAYER ME4 ;
  RECT 0.000 0.000 79.806 68.179 ;
  LAYER ME4 ;
  RECT 81.460 0.000 82.580 68.179 ;
  LAYER ME4 ;
  RECT 84.175 0.000 84.895 68.179 ;
  LAYER ME4 ;
  RECT 85.625 0.000 86.345 68.179 ;
  LAYER ME4 ;
  RECT 88.405 0.000 89.005 68.179 ;
  LAYER ME4 ;
  RECT 91.619 0.000 93.305 68.179 ;
  LAYER ME4 ;
  RECT 94.695 0.000 95.815 68.179 ;
  LAYER ME4 ;
  RECT 97.090 0.000 97.810 68.179 ;
  LAYER ME4 ;
  RECT 98.805 0.000 99.525 68.179 ;
  LAYER ME4 ;
  RECT 100.725 0.000 171.627 68.179 ;
END
END SYKB110_128X2X8CM4
END LIBRARY





