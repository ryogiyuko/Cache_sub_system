# ________________________________________________________________________________________________
# 
# 
#             Synchronous High-Density Single-Port SRAM Compiler
# 
#                 UMC 0.11um LL AE Logic Process
# 
# ________________________________________________________________________________________________
# 
#               
#         Copyright (C) 2024 Faraday Technology Corporation. All Rights Reserved.       
#                
#         This source code is an unpublished work belongs to Faraday Technology Corporation       
#         It is considered a trade secret and is not to be divulged or       
#         used by parties who have not received written authorization from       
#         Faraday Technology Corporation       
#                
#         Faraday's home page can be found at: http://www.faraday-tech.com/       
#                
# ________________________________________________________________________________________________
# 
#        IP Name            :  FSR0K_D_SH                
#        IP Version         :  1.3.0                     
#        IP Release Status  :  Active                    
#        Word               :  4096                      
#        Bit                :  8                         
#        Byte               :  8                         
#        Mux                :  1                         
#        Output Loading     :  0.01                      
#        Clock Input Slew   :  0.016                     
#        Data Input Slew    :  0.016                     
#        Ring Type          :  Ring Shape Model          
#        Ring Width         :  2                         
#        Bus Format         :  0                         
#        Memaker Path       :  /home/mem/Desktop/memlib  
#        GUI Version        :  m20230904                 
#        Date               :  2024/10/18 10:29:29       
# ________________________________________________________________________________________________
# 

VERSION 5.5 ;
NAMESCASESENSITIVE ON ;
MACRO SHKD110_4096X8X8BM1
CLASS BLOCK ;
FOREIGN SHKD110_4096X8X8BM1 0.000 0.000 ;
ORIGIN 0.000 0.000 ;
SIZE 1379.500 BY 551.210 ;
SYMMETRY x y r90 ;
SITE core ;
PIN DO63
  DIRECTION OUTPUT ;
 PORT
  LAYER ME4 ;
  RECT 1367.600 0.000 1368.400 1.000 ;
  LAYER ME3 ;
  RECT 1367.600 0.000 1368.400 1.000 ;
  LAYER ME2 ;
  RECT 1367.600 0.000 1368.400 1.000 ;
  LAYER ME1 ;
  RECT 1367.600 0.000 1368.400 1.000 ;
 END
 ANTENNAPARTIALMETALAREA                  4.152 LAYER ME2 ;
 ANTENNADIFFAREA                          5.472 LAYER ME2 ;
 ANTENNADIFFAREA                          5.472 LAYER ME3 ;
 ANTENNADIFFAREA                          5.472 LAYER ME4 ;
END DO63
PIN DI63
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 1352.800 0.000 1353.600 1.000 ;
  LAYER ME3 ;
  RECT 1352.800 0.000 1353.600 1.000 ;
  LAYER ME2 ;
  RECT 1352.800 0.000 1353.600 1.000 ;
  LAYER ME1 ;
  RECT 1352.800 0.000 1353.600 1.000 ;
 END
 ANTENNAPARTIALMETALAREA                  3.138 LAYER ME2 ;
 ANTENNAGATEAREA                          0.086 LAYER ME2 ;
 ANTENNAGATEAREA                          0.086 LAYER ME3 ;
 ANTENNAGATEAREA                          0.086 LAYER ME4 ;
 ANTENNADIFFAREA                          0.160 LAYER ME2 ;
 ANTENNADIFFAREA                          0.160 LAYER ME3 ;
 ANTENNADIFFAREA                          0.160 LAYER ME4 ;
 ANTENNAMAXAREACAR                       48.662 LAYER ME2 ;
 ANTENNAMAXAREACAR                       57.921 LAYER ME3 ;
 ANTENNAMAXAREACAR                       67.181 LAYER ME4 ;
END DI63
PIN DO62
  DIRECTION OUTPUT ;
 PORT
  LAYER ME4 ;
  RECT 1347.600 0.000 1348.400 1.000 ;
  LAYER ME3 ;
  RECT 1347.600 0.000 1348.400 1.000 ;
  LAYER ME2 ;
  RECT 1347.600 0.000 1348.400 1.000 ;
  LAYER ME1 ;
  RECT 1347.600 0.000 1348.400 1.000 ;
 END
 ANTENNAPARTIALMETALAREA                  4.160 LAYER ME2 ;
 ANTENNADIFFAREA                          5.472 LAYER ME2 ;
 ANTENNADIFFAREA                          5.472 LAYER ME3 ;
 ANTENNADIFFAREA                          5.472 LAYER ME4 ;
END DO62
PIN DI62
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 1333.200 0.000 1334.000 1.000 ;
  LAYER ME3 ;
  RECT 1333.200 0.000 1334.000 1.000 ;
  LAYER ME2 ;
  RECT 1333.200 0.000 1334.000 1.000 ;
  LAYER ME1 ;
  RECT 1333.200 0.000 1334.000 1.000 ;
 END
 ANTENNAPARTIALMETALAREA                  3.142 LAYER ME2 ;
 ANTENNAGATEAREA                          0.086 LAYER ME2 ;
 ANTENNAGATEAREA                          0.086 LAYER ME3 ;
 ANTENNAGATEAREA                          0.086 LAYER ME4 ;
 ANTENNADIFFAREA                          0.160 LAYER ME2 ;
 ANTENNADIFFAREA                          0.160 LAYER ME3 ;
 ANTENNADIFFAREA                          0.160 LAYER ME4 ;
 ANTENNAMAXAREACAR                       48.708 LAYER ME2 ;
 ANTENNAMAXAREACAR                       57.968 LAYER ME3 ;
 ANTENNAMAXAREACAR                       67.227 LAYER ME4 ;
END DI62
PIN DO61
  DIRECTION OUTPUT ;
 PORT
  LAYER ME4 ;
  RECT 1326.800 0.000 1327.600 1.000 ;
  LAYER ME3 ;
  RECT 1326.800 0.000 1327.600 1.000 ;
  LAYER ME2 ;
  RECT 1326.800 0.000 1327.600 1.000 ;
  LAYER ME1 ;
  RECT 1326.800 0.000 1327.600 1.000 ;
 END
 ANTENNAPARTIALMETALAREA                  4.176 LAYER ME2 ;
 ANTENNADIFFAREA                          5.472 LAYER ME2 ;
 ANTENNADIFFAREA                          5.472 LAYER ME3 ;
 ANTENNADIFFAREA                          5.472 LAYER ME4 ;
END DO61
PIN DI61
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 1312.000 0.000 1312.800 1.000 ;
  LAYER ME3 ;
  RECT 1312.000 0.000 1312.800 1.000 ;
  LAYER ME2 ;
  RECT 1312.000 0.000 1312.800 1.000 ;
  LAYER ME1 ;
  RECT 1312.000 0.000 1312.800 1.000 ;
 END
 ANTENNAPARTIALMETALAREA                  3.118 LAYER ME2 ;
 ANTENNAGATEAREA                          0.086 LAYER ME2 ;
 ANTENNAGATEAREA                          0.086 LAYER ME3 ;
 ANTENNAGATEAREA                          0.086 LAYER ME4 ;
 ANTENNADIFFAREA                          0.160 LAYER ME2 ;
 ANTENNADIFFAREA                          0.160 LAYER ME3 ;
 ANTENNADIFFAREA                          0.160 LAYER ME4 ;
 ANTENNAMAXAREACAR                       48.431 LAYER ME2 ;
 ANTENNAMAXAREACAR                       57.690 LAYER ME3 ;
 ANTENNAMAXAREACAR                       66.949 LAYER ME4 ;
END DI61
PIN DO60
  DIRECTION OUTPUT ;
 PORT
  LAYER ME4 ;
  RECT 1306.800 0.000 1307.600 1.000 ;
  LAYER ME3 ;
  RECT 1306.800 0.000 1307.600 1.000 ;
  LAYER ME2 ;
  RECT 1306.800 0.000 1307.600 1.000 ;
  LAYER ME1 ;
  RECT 1306.800 0.000 1307.600 1.000 ;
 END
 ANTENNAPARTIALMETALAREA                  4.144 LAYER ME2 ;
 ANTENNADIFFAREA                          5.472 LAYER ME2 ;
 ANTENNADIFFAREA                          5.472 LAYER ME3 ;
 ANTENNADIFFAREA                          5.472 LAYER ME4 ;
END DO60
PIN DI60
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 1292.000 0.000 1292.800 1.000 ;
  LAYER ME3 ;
  RECT 1292.000 0.000 1292.800 1.000 ;
  LAYER ME2 ;
  RECT 1292.000 0.000 1292.800 1.000 ;
  LAYER ME1 ;
  RECT 1292.000 0.000 1292.800 1.000 ;
 END
 ANTENNAPARTIALMETALAREA                  3.146 LAYER ME2 ;
 ANTENNAGATEAREA                          0.086 LAYER ME2 ;
 ANTENNAGATEAREA                          0.086 LAYER ME3 ;
 ANTENNAGATEAREA                          0.086 LAYER ME4 ;
 ANTENNADIFFAREA                          0.160 LAYER ME2 ;
 ANTENNADIFFAREA                          0.160 LAYER ME3 ;
 ANTENNADIFFAREA                          0.160 LAYER ME4 ;
 ANTENNAMAXAREACAR                       48.755 LAYER ME2 ;
 ANTENNAMAXAREACAR                       58.014 LAYER ME3 ;
 ANTENNAMAXAREACAR                       67.273 LAYER ME4 ;
END DI60
PIN DO59
  DIRECTION OUTPUT ;
 PORT
  LAYER ME4 ;
  RECT 1285.600 0.000 1286.400 1.000 ;
  LAYER ME3 ;
  RECT 1285.600 0.000 1286.400 1.000 ;
  LAYER ME2 ;
  RECT 1285.600 0.000 1286.400 1.000 ;
  LAYER ME1 ;
  RECT 1285.600 0.000 1286.400 1.000 ;
 END
 ANTENNAPARTIALMETALAREA                  4.160 LAYER ME2 ;
 ANTENNADIFFAREA                          5.472 LAYER ME2 ;
 ANTENNADIFFAREA                          5.472 LAYER ME3 ;
 ANTENNADIFFAREA                          5.472 LAYER ME4 ;
END DO59
PIN DI59
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 1271.200 0.000 1272.000 1.000 ;
  LAYER ME3 ;
  RECT 1271.200 0.000 1272.000 1.000 ;
  LAYER ME2 ;
  RECT 1271.200 0.000 1272.000 1.000 ;
  LAYER ME1 ;
  RECT 1271.200 0.000 1272.000 1.000 ;
 END
 ANTENNAPARTIALMETALAREA                  3.142 LAYER ME2 ;
 ANTENNAGATEAREA                          0.086 LAYER ME2 ;
 ANTENNAGATEAREA                          0.086 LAYER ME3 ;
 ANTENNAGATEAREA                          0.086 LAYER ME4 ;
 ANTENNADIFFAREA                          0.160 LAYER ME2 ;
 ANTENNADIFFAREA                          0.160 LAYER ME3 ;
 ANTENNADIFFAREA                          0.160 LAYER ME4 ;
 ANTENNAMAXAREACAR                       48.708 LAYER ME2 ;
 ANTENNAMAXAREACAR                       57.968 LAYER ME3 ;
 ANTENNAMAXAREACAR                       67.227 LAYER ME4 ;
END DI59
PIN DO58
  DIRECTION OUTPUT ;
 PORT
  LAYER ME4 ;
  RECT 1266.000 0.000 1266.800 1.000 ;
  LAYER ME3 ;
  RECT 1266.000 0.000 1266.800 1.000 ;
  LAYER ME2 ;
  RECT 1266.000 0.000 1266.800 1.000 ;
  LAYER ME1 ;
  RECT 1266.000 0.000 1266.800 1.000 ;
 END
 ANTENNAPARTIALMETALAREA                  4.168 LAYER ME2 ;
 ANTENNADIFFAREA                          5.472 LAYER ME2 ;
 ANTENNADIFFAREA                          5.472 LAYER ME3 ;
 ANTENNADIFFAREA                          5.472 LAYER ME4 ;
END DO58
PIN DI58
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 1251.200 0.000 1252.000 1.000 ;
  LAYER ME3 ;
  RECT 1251.200 0.000 1252.000 1.000 ;
  LAYER ME2 ;
  RECT 1251.200 0.000 1252.000 1.000 ;
  LAYER ME1 ;
  RECT 1251.200 0.000 1252.000 1.000 ;
 END
 ANTENNAPARTIALMETALAREA                  3.122 LAYER ME2 ;
 ANTENNAGATEAREA                          0.086 LAYER ME2 ;
 ANTENNAGATEAREA                          0.086 LAYER ME3 ;
 ANTENNAGATEAREA                          0.086 LAYER ME4 ;
 ANTENNADIFFAREA                          0.160 LAYER ME2 ;
 ANTENNADIFFAREA                          0.160 LAYER ME3 ;
 ANTENNADIFFAREA                          0.160 LAYER ME4 ;
 ANTENNAMAXAREACAR                       48.477 LAYER ME2 ;
 ANTENNAMAXAREACAR                       57.736 LAYER ME3 ;
 ANTENNAMAXAREACAR                       66.995 LAYER ME4 ;
END DI58
PIN DO57
  DIRECTION OUTPUT ;
 PORT
  LAYER ME4 ;
  RECT 1244.800 0.000 1245.600 1.000 ;
  LAYER ME3 ;
  RECT 1244.800 0.000 1245.600 1.000 ;
  LAYER ME2 ;
  RECT 1244.800 0.000 1245.600 1.000 ;
  LAYER ME1 ;
  RECT 1244.800 0.000 1245.600 1.000 ;
 END
 ANTENNAPARTIALMETALAREA                  4.144 LAYER ME2 ;
 ANTENNADIFFAREA                          5.472 LAYER ME2 ;
 ANTENNADIFFAREA                          5.472 LAYER ME3 ;
 ANTENNADIFFAREA                          5.472 LAYER ME4 ;
END DO57
PIN DI57
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 1230.000 0.000 1230.800 1.000 ;
  LAYER ME3 ;
  RECT 1230.000 0.000 1230.800 1.000 ;
  LAYER ME2 ;
  RECT 1230.000 0.000 1230.800 1.000 ;
  LAYER ME1 ;
  RECT 1230.000 0.000 1230.800 1.000 ;
 END
 ANTENNAPARTIALMETALAREA                  3.146 LAYER ME2 ;
 ANTENNAGATEAREA                          0.086 LAYER ME2 ;
 ANTENNAGATEAREA                          0.086 LAYER ME3 ;
 ANTENNAGATEAREA                          0.086 LAYER ME4 ;
 ANTENNADIFFAREA                          0.160 LAYER ME2 ;
 ANTENNADIFFAREA                          0.160 LAYER ME3 ;
 ANTENNADIFFAREA                          0.160 LAYER ME4 ;
 ANTENNAMAXAREACAR                       48.755 LAYER ME2 ;
 ANTENNAMAXAREACAR                       58.014 LAYER ME3 ;
 ANTENNAMAXAREACAR                       67.273 LAYER ME4 ;
END DI57
PIN DO56
  DIRECTION OUTPUT ;
 PORT
  LAYER ME4 ;
  RECT 1224.800 0.000 1225.600 1.000 ;
  LAYER ME3 ;
  RECT 1224.800 0.000 1225.600 1.000 ;
  LAYER ME2 ;
  RECT 1224.800 0.000 1225.600 1.000 ;
  LAYER ME1 ;
  RECT 1224.800 0.000 1225.600 1.000 ;
 END
 ANTENNAPARTIALMETALAREA                  4.168 LAYER ME2 ;
 ANTENNADIFFAREA                          5.472 LAYER ME2 ;
 ANTENNADIFFAREA                          5.472 LAYER ME3 ;
 ANTENNADIFFAREA                          5.472 LAYER ME4 ;
END DO56
PIN WEB7
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 1212.000 0.000 1212.800 1.000 ;
  LAYER ME3 ;
  RECT 1212.000 0.000 1212.800 1.000 ;
  LAYER ME2 ;
  RECT 1212.000 0.000 1212.800 1.000 ;
  LAYER ME1 ;
  RECT 1212.000 0.000 1212.800 1.000 ;
 END
 ANTENNAPARTIALMETALAREA                  2.836 LAYER ME2 ;
 ANTENNAGATEAREA                          0.072 LAYER ME2 ;
 ANTENNAGATEAREA                          0.072 LAYER ME3 ;
 ANTENNAGATEAREA                          0.072 LAYER ME4 ;
 ANTENNADIFFAREA                          0.160 LAYER ME2 ;
 ANTENNADIFFAREA                          0.160 LAYER ME3 ;
 ANTENNADIFFAREA                          0.160 LAYER ME4 ;
 ANTENNAMAXAREACAR                       54.400 LAYER ME2 ;
 ANTENNAMAXAREACAR                       65.511 LAYER ME3 ;
 ANTENNAMAXAREACAR                       76.622 LAYER ME4 ;
END WEB7
PIN DI56
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 1210.400 0.000 1211.200 1.000 ;
  LAYER ME3 ;
  RECT 1210.400 0.000 1211.200 1.000 ;
  LAYER ME2 ;
  RECT 1210.400 0.000 1211.200 1.000 ;
  LAYER ME1 ;
  RECT 1210.400 0.000 1211.200 1.000 ;
 END
 ANTENNAPARTIALMETALAREA                  3.134 LAYER ME2 ;
 ANTENNAGATEAREA                          0.086 LAYER ME2 ;
 ANTENNAGATEAREA                          0.086 LAYER ME3 ;
 ANTENNAGATEAREA                          0.086 LAYER ME4 ;
 ANTENNADIFFAREA                          0.160 LAYER ME2 ;
 ANTENNADIFFAREA                          0.160 LAYER ME3 ;
 ANTENNADIFFAREA                          0.160 LAYER ME4 ;
 ANTENNAMAXAREACAR                       48.616 LAYER ME2 ;
 ANTENNAMAXAREACAR                       57.875 LAYER ME3 ;
 ANTENNAMAXAREACAR                       67.134 LAYER ME4 ;
END DI56
PIN DO55
  DIRECTION OUTPUT ;
 PORT
  LAYER ME4 ;
  RECT 1204.000 0.000 1204.800 1.000 ;
  LAYER ME3 ;
  RECT 1204.000 0.000 1204.800 1.000 ;
  LAYER ME2 ;
  RECT 1204.000 0.000 1204.800 1.000 ;
  LAYER ME1 ;
  RECT 1204.000 0.000 1204.800 1.000 ;
 END
 ANTENNAPARTIALMETALAREA                  4.168 LAYER ME2 ;
 ANTENNADIFFAREA                          5.472 LAYER ME2 ;
 ANTENNADIFFAREA                          5.472 LAYER ME3 ;
 ANTENNADIFFAREA                          5.472 LAYER ME4 ;
END DO55
PIN DI55
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 1189.200 0.000 1190.000 1.000 ;
  LAYER ME3 ;
  RECT 1189.200 0.000 1190.000 1.000 ;
  LAYER ME2 ;
  RECT 1189.200 0.000 1190.000 1.000 ;
  LAYER ME1 ;
  RECT 1189.200 0.000 1190.000 1.000 ;
 END
 ANTENNAPARTIALMETALAREA                  3.122 LAYER ME2 ;
 ANTENNAGATEAREA                          0.086 LAYER ME2 ;
 ANTENNAGATEAREA                          0.086 LAYER ME3 ;
 ANTENNAGATEAREA                          0.086 LAYER ME4 ;
 ANTENNADIFFAREA                          0.160 LAYER ME2 ;
 ANTENNADIFFAREA                          0.160 LAYER ME3 ;
 ANTENNADIFFAREA                          0.160 LAYER ME4 ;
 ANTENNAMAXAREACAR                       48.477 LAYER ME2 ;
 ANTENNAMAXAREACAR                       57.736 LAYER ME3 ;
 ANTENNAMAXAREACAR                       66.995 LAYER ME4 ;
END DI55
PIN DO54
  DIRECTION OUTPUT ;
 PORT
  LAYER ME4 ;
  RECT 1184.000 0.000 1184.800 1.000 ;
  LAYER ME3 ;
  RECT 1184.000 0.000 1184.800 1.000 ;
  LAYER ME2 ;
  RECT 1184.000 0.000 1184.800 1.000 ;
  LAYER ME1 ;
  RECT 1184.000 0.000 1184.800 1.000 ;
 END
 ANTENNAPARTIALMETALAREA                  4.144 LAYER ME2 ;
 ANTENNADIFFAREA                          5.472 LAYER ME2 ;
 ANTENNADIFFAREA                          5.472 LAYER ME3 ;
 ANTENNADIFFAREA                          5.472 LAYER ME4 ;
END DO54
PIN DI54
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 1169.200 0.000 1170.000 1.000 ;
  LAYER ME3 ;
  RECT 1169.200 0.000 1170.000 1.000 ;
  LAYER ME2 ;
  RECT 1169.200 0.000 1170.000 1.000 ;
  LAYER ME1 ;
  RECT 1169.200 0.000 1170.000 1.000 ;
 END
 ANTENNAPARTIALMETALAREA                  3.154 LAYER ME2 ;
 ANTENNAGATEAREA                          0.086 LAYER ME2 ;
 ANTENNAGATEAREA                          0.086 LAYER ME3 ;
 ANTENNAGATEAREA                          0.086 LAYER ME4 ;
 ANTENNADIFFAREA                          0.160 LAYER ME2 ;
 ANTENNADIFFAREA                          0.160 LAYER ME3 ;
 ANTENNADIFFAREA                          0.160 LAYER ME4 ;
 ANTENNAMAXAREACAR                       48.847 LAYER ME2 ;
 ANTENNAMAXAREACAR                       58.106 LAYER ME3 ;
 ANTENNAMAXAREACAR                       67.366 LAYER ME4 ;
END DI54
PIN DO53
  DIRECTION OUTPUT ;
 PORT
  LAYER ME4 ;
  RECT 1162.800 0.000 1163.600 1.000 ;
  LAYER ME3 ;
  RECT 1162.800 0.000 1163.600 1.000 ;
  LAYER ME2 ;
  RECT 1162.800 0.000 1163.600 1.000 ;
  LAYER ME1 ;
  RECT 1162.800 0.000 1163.600 1.000 ;
 END
 ANTENNAPARTIALMETALAREA                  4.168 LAYER ME2 ;
 ANTENNADIFFAREA                          5.472 LAYER ME2 ;
 ANTENNADIFFAREA                          5.472 LAYER ME3 ;
 ANTENNADIFFAREA                          5.472 LAYER ME4 ;
END DO53
PIN DI53
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 1148.400 0.000 1149.200 1.000 ;
  LAYER ME3 ;
  RECT 1148.400 0.000 1149.200 1.000 ;
  LAYER ME2 ;
  RECT 1148.400 0.000 1149.200 1.000 ;
  LAYER ME1 ;
  RECT 1148.400 0.000 1149.200 1.000 ;
 END
 ANTENNAPARTIALMETALAREA                  3.134 LAYER ME2 ;
 ANTENNAGATEAREA                          0.086 LAYER ME2 ;
 ANTENNAGATEAREA                          0.086 LAYER ME3 ;
 ANTENNAGATEAREA                          0.086 LAYER ME4 ;
 ANTENNADIFFAREA                          0.160 LAYER ME2 ;
 ANTENNADIFFAREA                          0.160 LAYER ME3 ;
 ANTENNADIFFAREA                          0.160 LAYER ME4 ;
 ANTENNAMAXAREACAR                       48.616 LAYER ME2 ;
 ANTENNAMAXAREACAR                       57.875 LAYER ME3 ;
 ANTENNAMAXAREACAR                       67.134 LAYER ME4 ;
END DI53
PIN DO52
  DIRECTION OUTPUT ;
 PORT
  LAYER ME4 ;
  RECT 1143.200 0.000 1144.000 1.000 ;
  LAYER ME3 ;
  RECT 1143.200 0.000 1144.000 1.000 ;
  LAYER ME2 ;
  RECT 1143.200 0.000 1144.000 1.000 ;
  LAYER ME1 ;
  RECT 1143.200 0.000 1144.000 1.000 ;
 END
 ANTENNAPARTIALMETALAREA                  4.160 LAYER ME2 ;
 ANTENNADIFFAREA                          5.472 LAYER ME2 ;
 ANTENNADIFFAREA                          5.472 LAYER ME3 ;
 ANTENNADIFFAREA                          5.472 LAYER ME4 ;
END DO52
PIN DI52
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 1128.400 0.000 1129.200 1.000 ;
  LAYER ME3 ;
  RECT 1128.400 0.000 1129.200 1.000 ;
  LAYER ME2 ;
  RECT 1128.400 0.000 1129.200 1.000 ;
  LAYER ME1 ;
  RECT 1128.400 0.000 1129.200 1.000 ;
 END
 ANTENNAPARTIALMETALAREA                  3.130 LAYER ME2 ;
 ANTENNAGATEAREA                          0.086 LAYER ME2 ;
 ANTENNAGATEAREA                          0.086 LAYER ME3 ;
 ANTENNAGATEAREA                          0.086 LAYER ME4 ;
 ANTENNADIFFAREA                          0.160 LAYER ME2 ;
 ANTENNADIFFAREA                          0.160 LAYER ME3 ;
 ANTENNADIFFAREA                          0.160 LAYER ME4 ;
 ANTENNAMAXAREACAR                       48.569 LAYER ME2 ;
 ANTENNAMAXAREACAR                       57.829 LAYER ME3 ;
 ANTENNAMAXAREACAR                       67.088 LAYER ME4 ;
END DI52
PIN DO51
  DIRECTION OUTPUT ;
 PORT
  LAYER ME4 ;
  RECT 1122.000 0.000 1122.800 1.000 ;
  LAYER ME3 ;
  RECT 1122.000 0.000 1122.800 1.000 ;
  LAYER ME2 ;
  RECT 1122.000 0.000 1122.800 1.000 ;
  LAYER ME1 ;
  RECT 1122.000 0.000 1122.800 1.000 ;
 END
 ANTENNAPARTIALMETALAREA                  4.144 LAYER ME2 ;
 ANTENNADIFFAREA                          5.472 LAYER ME2 ;
 ANTENNADIFFAREA                          5.472 LAYER ME3 ;
 ANTENNADIFFAREA                          5.472 LAYER ME4 ;
END DO51
PIN DI51
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 1107.200 0.000 1108.000 1.000 ;
  LAYER ME3 ;
  RECT 1107.200 0.000 1108.000 1.000 ;
  LAYER ME2 ;
  RECT 1107.200 0.000 1108.000 1.000 ;
  LAYER ME1 ;
  RECT 1107.200 0.000 1108.000 1.000 ;
 END
 ANTENNAPARTIALMETALAREA                  3.154 LAYER ME2 ;
 ANTENNAGATEAREA                          0.086 LAYER ME2 ;
 ANTENNAGATEAREA                          0.086 LAYER ME3 ;
 ANTENNAGATEAREA                          0.086 LAYER ME4 ;
 ANTENNADIFFAREA                          0.160 LAYER ME2 ;
 ANTENNADIFFAREA                          0.160 LAYER ME3 ;
 ANTENNADIFFAREA                          0.160 LAYER ME4 ;
 ANTENNAMAXAREACAR                       48.847 LAYER ME2 ;
 ANTENNAMAXAREACAR                       58.106 LAYER ME3 ;
 ANTENNAMAXAREACAR                       67.366 LAYER ME4 ;
END DI51
PIN DO50
  DIRECTION OUTPUT ;
 PORT
  LAYER ME4 ;
  RECT 1102.000 0.000 1102.800 1.000 ;
  LAYER ME3 ;
  RECT 1102.000 0.000 1102.800 1.000 ;
  LAYER ME2 ;
  RECT 1102.000 0.000 1102.800 1.000 ;
  LAYER ME1 ;
  RECT 1102.000 0.000 1102.800 1.000 ;
 END
 ANTENNAPARTIALMETALAREA                  4.176 LAYER ME2 ;
 ANTENNADIFFAREA                          5.472 LAYER ME2 ;
 ANTENNADIFFAREA                          5.472 LAYER ME3 ;
 ANTENNADIFFAREA                          5.472 LAYER ME4 ;
END DO50
PIN DI50
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 1087.600 0.000 1088.400 1.000 ;
  LAYER ME3 ;
  RECT 1087.600 0.000 1088.400 1.000 ;
  LAYER ME2 ;
  RECT 1087.600 0.000 1088.400 1.000 ;
  LAYER ME1 ;
  RECT 1087.600 0.000 1088.400 1.000 ;
 END
 ANTENNAPARTIALMETALAREA                  3.126 LAYER ME2 ;
 ANTENNAGATEAREA                          0.086 LAYER ME2 ;
 ANTENNAGATEAREA                          0.086 LAYER ME3 ;
 ANTENNAGATEAREA                          0.086 LAYER ME4 ;
 ANTENNADIFFAREA                          0.160 LAYER ME2 ;
 ANTENNADIFFAREA                          0.160 LAYER ME3 ;
 ANTENNADIFFAREA                          0.160 LAYER ME4 ;
 ANTENNAMAXAREACAR                       48.523 LAYER ME2 ;
 ANTENNAMAXAREACAR                       57.782 LAYER ME3 ;
 ANTENNAMAXAREACAR                       67.042 LAYER ME4 ;
END DI50
PIN DO49
  DIRECTION OUTPUT ;
 PORT
  LAYER ME4 ;
  RECT 1081.200 0.000 1082.000 1.000 ;
  LAYER ME3 ;
  RECT 1081.200 0.000 1082.000 1.000 ;
  LAYER ME2 ;
  RECT 1081.200 0.000 1082.000 1.000 ;
  LAYER ME1 ;
  RECT 1081.200 0.000 1082.000 1.000 ;
 END
 ANTENNAPARTIALMETALAREA                  4.160 LAYER ME2 ;
 ANTENNADIFFAREA                          5.472 LAYER ME2 ;
 ANTENNADIFFAREA                          5.472 LAYER ME3 ;
 ANTENNADIFFAREA                          5.472 LAYER ME4 ;
END DO49
PIN DI49
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 1066.400 0.000 1067.200 1.000 ;
  LAYER ME3 ;
  RECT 1066.400 0.000 1067.200 1.000 ;
  LAYER ME2 ;
  RECT 1066.400 0.000 1067.200 1.000 ;
  LAYER ME1 ;
  RECT 1066.400 0.000 1067.200 1.000 ;
 END
 ANTENNAPARTIALMETALAREA                  3.130 LAYER ME2 ;
 ANTENNAGATEAREA                          0.086 LAYER ME2 ;
 ANTENNAGATEAREA                          0.086 LAYER ME3 ;
 ANTENNAGATEAREA                          0.086 LAYER ME4 ;
 ANTENNADIFFAREA                          0.160 LAYER ME2 ;
 ANTENNADIFFAREA                          0.160 LAYER ME3 ;
 ANTENNADIFFAREA                          0.160 LAYER ME4 ;
 ANTENNAMAXAREACAR                       48.569 LAYER ME2 ;
 ANTENNAMAXAREACAR                       57.829 LAYER ME3 ;
 ANTENNAMAXAREACAR                       67.088 LAYER ME4 ;
END DI49
PIN DO48
  DIRECTION OUTPUT ;
 PORT
  LAYER ME4 ;
  RECT 1061.200 0.000 1062.000 1.000 ;
  LAYER ME3 ;
  RECT 1061.200 0.000 1062.000 1.000 ;
  LAYER ME2 ;
  RECT 1061.200 0.000 1062.000 1.000 ;
  LAYER ME1 ;
  RECT 1061.200 0.000 1062.000 1.000 ;
 END
 ANTENNAPARTIALMETALAREA                  4.152 LAYER ME2 ;
 ANTENNADIFFAREA                          5.472 LAYER ME2 ;
 ANTENNADIFFAREA                          5.472 LAYER ME3 ;
 ANTENNADIFFAREA                          5.472 LAYER ME4 ;
END DO48
PIN WEB6
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 1048.400 0.000 1049.200 1.000 ;
  LAYER ME3 ;
  RECT 1048.400 0.000 1049.200 1.000 ;
  LAYER ME2 ;
  RECT 1048.400 0.000 1049.200 1.000 ;
  LAYER ME1 ;
  RECT 1048.400 0.000 1049.200 1.000 ;
 END
 ANTENNAPARTIALMETALAREA                  2.840 LAYER ME2 ;
 ANTENNAGATEAREA                          0.072 LAYER ME2 ;
 ANTENNAGATEAREA                          0.072 LAYER ME3 ;
 ANTENNAGATEAREA                          0.072 LAYER ME4 ;
 ANTENNADIFFAREA                          0.160 LAYER ME2 ;
 ANTENNADIFFAREA                          0.160 LAYER ME3 ;
 ANTENNADIFFAREA                          0.160 LAYER ME4 ;
 ANTENNAMAXAREACAR                       54.456 LAYER ME2 ;
 ANTENNAMAXAREACAR                       65.567 LAYER ME3 ;
 ANTENNAMAXAREACAR                       76.678 LAYER ME4 ;
END WEB6
PIN DI48
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 1046.800 0.000 1047.600 1.000 ;
  LAYER ME3 ;
  RECT 1046.800 0.000 1047.600 1.000 ;
  LAYER ME2 ;
  RECT 1046.800 0.000 1047.600 1.000 ;
  LAYER ME1 ;
  RECT 1046.800 0.000 1047.600 1.000 ;
 END
 ANTENNAPARTIALMETALAREA                  3.150 LAYER ME2 ;
 ANTENNAGATEAREA                          0.086 LAYER ME2 ;
 ANTENNAGATEAREA                          0.086 LAYER ME3 ;
 ANTENNAGATEAREA                          0.086 LAYER ME4 ;
 ANTENNADIFFAREA                          0.160 LAYER ME2 ;
 ANTENNADIFFAREA                          0.160 LAYER ME3 ;
 ANTENNADIFFAREA                          0.160 LAYER ME4 ;
 ANTENNAMAXAREACAR                       48.801 LAYER ME2 ;
 ANTENNAMAXAREACAR                       58.060 LAYER ME3 ;
 ANTENNAMAXAREACAR                       67.319 LAYER ME4 ;
END DI48
PIN DO47
  DIRECTION OUTPUT ;
 PORT
  LAYER ME4 ;
  RECT 1040.000 0.000 1040.800 1.000 ;
  LAYER ME3 ;
  RECT 1040.000 0.000 1040.800 1.000 ;
  LAYER ME2 ;
  RECT 1040.000 0.000 1040.800 1.000 ;
  LAYER ME1 ;
  RECT 1040.000 0.000 1040.800 1.000 ;
 END
 ANTENNAPARTIALMETALAREA                  4.176 LAYER ME2 ;
 ANTENNADIFFAREA                          5.472 LAYER ME2 ;
 ANTENNADIFFAREA                          5.472 LAYER ME3 ;
 ANTENNADIFFAREA                          5.472 LAYER ME4 ;
END DO47
PIN DI47
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 1025.600 0.000 1026.400 1.000 ;
  LAYER ME3 ;
  RECT 1025.600 0.000 1026.400 1.000 ;
  LAYER ME2 ;
  RECT 1025.600 0.000 1026.400 1.000 ;
  LAYER ME1 ;
  RECT 1025.600 0.000 1026.400 1.000 ;
 END
 ANTENNAPARTIALMETALAREA                  3.126 LAYER ME2 ;
 ANTENNAGATEAREA                          0.086 LAYER ME2 ;
 ANTENNAGATEAREA                          0.086 LAYER ME3 ;
 ANTENNAGATEAREA                          0.086 LAYER ME4 ;
 ANTENNADIFFAREA                          0.160 LAYER ME2 ;
 ANTENNADIFFAREA                          0.160 LAYER ME3 ;
 ANTENNADIFFAREA                          0.160 LAYER ME4 ;
 ANTENNAMAXAREACAR                       48.523 LAYER ME2 ;
 ANTENNAMAXAREACAR                       57.782 LAYER ME3 ;
 ANTENNAMAXAREACAR                       67.042 LAYER ME4 ;
END DI47
PIN DO46
  DIRECTION OUTPUT ;
 PORT
  LAYER ME4 ;
  RECT 1020.400 0.000 1021.200 1.000 ;
  LAYER ME3 ;
  RECT 1020.400 0.000 1021.200 1.000 ;
  LAYER ME2 ;
  RECT 1020.400 0.000 1021.200 1.000 ;
  LAYER ME1 ;
  RECT 1020.400 0.000 1021.200 1.000 ;
 END
 ANTENNAPARTIALMETALAREA                  4.152 LAYER ME2 ;
 ANTENNADIFFAREA                          5.472 LAYER ME2 ;
 ANTENNADIFFAREA                          5.472 LAYER ME3 ;
 ANTENNADIFFAREA                          5.472 LAYER ME4 ;
END DO46
PIN DI46
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 1005.600 0.000 1006.400 1.000 ;
  LAYER ME3 ;
  RECT 1005.600 0.000 1006.400 1.000 ;
  LAYER ME2 ;
  RECT 1005.600 0.000 1006.400 1.000 ;
  LAYER ME1 ;
  RECT 1005.600 0.000 1006.400 1.000 ;
 END
 ANTENNAPARTIALMETALAREA                  3.138 LAYER ME2 ;
 ANTENNAGATEAREA                          0.086 LAYER ME2 ;
 ANTENNAGATEAREA                          0.086 LAYER ME3 ;
 ANTENNAGATEAREA                          0.086 LAYER ME4 ;
 ANTENNADIFFAREA                          0.160 LAYER ME2 ;
 ANTENNADIFFAREA                          0.160 LAYER ME3 ;
 ANTENNADIFFAREA                          0.160 LAYER ME4 ;
 ANTENNAMAXAREACAR                       48.662 LAYER ME2 ;
 ANTENNAMAXAREACAR                       57.921 LAYER ME3 ;
 ANTENNAMAXAREACAR                       67.181 LAYER ME4 ;
END DI46
PIN DO45
  DIRECTION OUTPUT ;
 PORT
  LAYER ME4 ;
  RECT 999.200 0.000 1000.000 1.000 ;
  LAYER ME3 ;
  RECT 999.200 0.000 1000.000 1.000 ;
  LAYER ME2 ;
  RECT 999.200 0.000 1000.000 1.000 ;
  LAYER ME1 ;
  RECT 999.200 0.000 1000.000 1.000 ;
 END
 ANTENNAPARTIALMETALAREA                  4.152 LAYER ME2 ;
 ANTENNADIFFAREA                          5.472 LAYER ME2 ;
 ANTENNADIFFAREA                          5.472 LAYER ME3 ;
 ANTENNADIFFAREA                          5.472 LAYER ME4 ;
END DO45
PIN DI45
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 984.800 0.000 985.600 1.000 ;
  LAYER ME3 ;
  RECT 984.800 0.000 985.600 1.000 ;
  LAYER ME2 ;
  RECT 984.800 0.000 985.600 1.000 ;
  LAYER ME1 ;
  RECT 984.800 0.000 985.600 1.000 ;
 END
 ANTENNAPARTIALMETALAREA                  3.150 LAYER ME2 ;
 ANTENNAGATEAREA                          0.086 LAYER ME2 ;
 ANTENNAGATEAREA                          0.086 LAYER ME3 ;
 ANTENNAGATEAREA                          0.086 LAYER ME4 ;
 ANTENNADIFFAREA                          0.160 LAYER ME2 ;
 ANTENNADIFFAREA                          0.160 LAYER ME3 ;
 ANTENNADIFFAREA                          0.160 LAYER ME4 ;
 ANTENNAMAXAREACAR                       48.801 LAYER ME2 ;
 ANTENNAMAXAREACAR                       58.060 LAYER ME3 ;
 ANTENNAMAXAREACAR                       67.319 LAYER ME4 ;
END DI45
PIN DO44
  DIRECTION OUTPUT ;
 PORT
  LAYER ME4 ;
  RECT 979.600 0.000 980.400 1.000 ;
  LAYER ME3 ;
  RECT 979.600 0.000 980.400 1.000 ;
  LAYER ME2 ;
  RECT 979.600 0.000 980.400 1.000 ;
  LAYER ME1 ;
  RECT 979.600 0.000 980.400 1.000 ;
 END
 ANTENNAPARTIALMETALAREA                  4.176 LAYER ME2 ;
 ANTENNADIFFAREA                          5.472 LAYER ME2 ;
 ANTENNADIFFAREA                          5.472 LAYER ME3 ;
 ANTENNADIFFAREA                          5.472 LAYER ME4 ;
END DO44
PIN DI44
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 964.800 0.000 965.600 1.000 ;
  LAYER ME3 ;
  RECT 964.800 0.000 965.600 1.000 ;
  LAYER ME2 ;
  RECT 964.800 0.000 965.600 1.000 ;
  LAYER ME1 ;
  RECT 964.800 0.000 965.600 1.000 ;
 END
 ANTENNAPARTIALMETALAREA                  3.118 LAYER ME2 ;
 ANTENNAGATEAREA                          0.086 LAYER ME2 ;
 ANTENNAGATEAREA                          0.086 LAYER ME3 ;
 ANTENNAGATEAREA                          0.086 LAYER ME4 ;
 ANTENNADIFFAREA                          0.160 LAYER ME2 ;
 ANTENNADIFFAREA                          0.160 LAYER ME3 ;
 ANTENNADIFFAREA                          0.160 LAYER ME4 ;
 ANTENNAMAXAREACAR                       48.431 LAYER ME2 ;
 ANTENNAMAXAREACAR                       57.690 LAYER ME3 ;
 ANTENNAMAXAREACAR                       66.949 LAYER ME4 ;
END DI44
PIN DO43
  DIRECTION OUTPUT ;
 PORT
  LAYER ME4 ;
  RECT 958.400 0.000 959.200 1.000 ;
  LAYER ME3 ;
  RECT 958.400 0.000 959.200 1.000 ;
  LAYER ME2 ;
  RECT 958.400 0.000 959.200 1.000 ;
  LAYER ME1 ;
  RECT 958.400 0.000 959.200 1.000 ;
 END
 ANTENNAPARTIALMETALAREA                  4.152 LAYER ME2 ;
 ANTENNADIFFAREA                          5.472 LAYER ME2 ;
 ANTENNADIFFAREA                          5.472 LAYER ME3 ;
 ANTENNADIFFAREA                          5.472 LAYER ME4 ;
END DO43
PIN DI43
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 943.600 0.000 944.400 1.000 ;
  LAYER ME3 ;
  RECT 943.600 0.000 944.400 1.000 ;
  LAYER ME2 ;
  RECT 943.600 0.000 944.400 1.000 ;
  LAYER ME1 ;
  RECT 943.600 0.000 944.400 1.000 ;
 END
 ANTENNAPARTIALMETALAREA                  3.138 LAYER ME2 ;
 ANTENNAGATEAREA                          0.086 LAYER ME2 ;
 ANTENNAGATEAREA                          0.086 LAYER ME3 ;
 ANTENNAGATEAREA                          0.086 LAYER ME4 ;
 ANTENNADIFFAREA                          0.160 LAYER ME2 ;
 ANTENNADIFFAREA                          0.160 LAYER ME3 ;
 ANTENNADIFFAREA                          0.160 LAYER ME4 ;
 ANTENNAMAXAREACAR                       48.662 LAYER ME2 ;
 ANTENNAMAXAREACAR                       57.921 LAYER ME3 ;
 ANTENNAMAXAREACAR                       67.181 LAYER ME4 ;
END DI43
PIN DO42
  DIRECTION OUTPUT ;
 PORT
  LAYER ME4 ;
  RECT 938.400 0.000 939.200 1.000 ;
  LAYER ME3 ;
  RECT 938.400 0.000 939.200 1.000 ;
  LAYER ME2 ;
  RECT 938.400 0.000 939.200 1.000 ;
  LAYER ME1 ;
  RECT 938.400 0.000 939.200 1.000 ;
 END
 ANTENNAPARTIALMETALAREA                  4.160 LAYER ME2 ;
 ANTENNADIFFAREA                          5.472 LAYER ME2 ;
 ANTENNADIFFAREA                          5.472 LAYER ME3 ;
 ANTENNADIFFAREA                          5.472 LAYER ME4 ;
END DO42
PIN DI42
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 924.000 0.000 924.800 1.000 ;
  LAYER ME3 ;
  RECT 924.000 0.000 924.800 1.000 ;
  LAYER ME2 ;
  RECT 924.000 0.000 924.800 1.000 ;
  LAYER ME1 ;
  RECT 924.000 0.000 924.800 1.000 ;
 END
 ANTENNAPARTIALMETALAREA                  3.142 LAYER ME2 ;
 ANTENNAGATEAREA                          0.086 LAYER ME2 ;
 ANTENNAGATEAREA                          0.086 LAYER ME3 ;
 ANTENNAGATEAREA                          0.086 LAYER ME4 ;
 ANTENNADIFFAREA                          0.160 LAYER ME2 ;
 ANTENNADIFFAREA                          0.160 LAYER ME3 ;
 ANTENNADIFFAREA                          0.160 LAYER ME4 ;
 ANTENNAMAXAREACAR                       48.708 LAYER ME2 ;
 ANTENNAMAXAREACAR                       57.968 LAYER ME3 ;
 ANTENNAMAXAREACAR                       67.227 LAYER ME4 ;
END DI42
PIN DO41
  DIRECTION OUTPUT ;
 PORT
  LAYER ME4 ;
  RECT 917.600 0.000 918.400 1.000 ;
  LAYER ME3 ;
  RECT 917.600 0.000 918.400 1.000 ;
  LAYER ME2 ;
  RECT 917.600 0.000 918.400 1.000 ;
  LAYER ME1 ;
  RECT 917.600 0.000 918.400 1.000 ;
 END
 ANTENNAPARTIALMETALAREA                  4.176 LAYER ME2 ;
 ANTENNADIFFAREA                          5.472 LAYER ME2 ;
 ANTENNADIFFAREA                          5.472 LAYER ME3 ;
 ANTENNADIFFAREA                          5.472 LAYER ME4 ;
END DO41
PIN DI41
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 902.800 0.000 903.600 1.000 ;
  LAYER ME3 ;
  RECT 902.800 0.000 903.600 1.000 ;
  LAYER ME2 ;
  RECT 902.800 0.000 903.600 1.000 ;
  LAYER ME1 ;
  RECT 902.800 0.000 903.600 1.000 ;
 END
 ANTENNAPARTIALMETALAREA                  3.118 LAYER ME2 ;
 ANTENNAGATEAREA                          0.086 LAYER ME2 ;
 ANTENNAGATEAREA                          0.086 LAYER ME3 ;
 ANTENNAGATEAREA                          0.086 LAYER ME4 ;
 ANTENNADIFFAREA                          0.160 LAYER ME2 ;
 ANTENNADIFFAREA                          0.160 LAYER ME3 ;
 ANTENNADIFFAREA                          0.160 LAYER ME4 ;
 ANTENNAMAXAREACAR                       48.431 LAYER ME2 ;
 ANTENNAMAXAREACAR                       57.690 LAYER ME3 ;
 ANTENNAMAXAREACAR                       66.949 LAYER ME4 ;
END DI41
PIN DO40
  DIRECTION OUTPUT ;
 PORT
  LAYER ME4 ;
  RECT 897.600 0.000 898.400 1.000 ;
  LAYER ME3 ;
  RECT 897.600 0.000 898.400 1.000 ;
  LAYER ME2 ;
  RECT 897.600 0.000 898.400 1.000 ;
  LAYER ME1 ;
  RECT 897.600 0.000 898.400 1.000 ;
 END
 ANTENNAPARTIALMETALAREA                  4.144 LAYER ME2 ;
 ANTENNADIFFAREA                          5.472 LAYER ME2 ;
 ANTENNADIFFAREA                          5.472 LAYER ME3 ;
 ANTENNADIFFAREA                          5.472 LAYER ME4 ;
END DO40
PIN WEB5
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 884.800 0.000 885.600 1.000 ;
  LAYER ME3 ;
  RECT 884.800 0.000 885.600 1.000 ;
  LAYER ME2 ;
  RECT 884.800 0.000 885.600 1.000 ;
  LAYER ME1 ;
  RECT 884.800 0.000 885.600 1.000 ;
 END
 ANTENNAPARTIALMETALAREA                  2.856 LAYER ME2 ;
 ANTENNAGATEAREA                          0.072 LAYER ME2 ;
 ANTENNAGATEAREA                          0.072 LAYER ME3 ;
 ANTENNAGATEAREA                          0.072 LAYER ME4 ;
 ANTENNADIFFAREA                          0.160 LAYER ME2 ;
 ANTENNADIFFAREA                          0.160 LAYER ME3 ;
 ANTENNADIFFAREA                          0.160 LAYER ME4 ;
 ANTENNAMAXAREACAR                       54.678 LAYER ME2 ;
 ANTENNAMAXAREACAR                       65.789 LAYER ME3 ;
 ANTENNAMAXAREACAR                       76.900 LAYER ME4 ;
END WEB5
PIN DI40
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 882.800 0.000 883.600 1.000 ;
  LAYER ME3 ;
  RECT 882.800 0.000 883.600 1.000 ;
  LAYER ME2 ;
  RECT 882.800 0.000 883.600 1.000 ;
  LAYER ME1 ;
  RECT 882.800 0.000 883.600 1.000 ;
 END
 ANTENNAPARTIALMETALAREA                  3.146 LAYER ME2 ;
 ANTENNAGATEAREA                          0.086 LAYER ME2 ;
 ANTENNAGATEAREA                          0.086 LAYER ME3 ;
 ANTENNAGATEAREA                          0.086 LAYER ME4 ;
 ANTENNADIFFAREA                          0.160 LAYER ME2 ;
 ANTENNADIFFAREA                          0.160 LAYER ME3 ;
 ANTENNADIFFAREA                          0.160 LAYER ME4 ;
 ANTENNAMAXAREACAR                       48.755 LAYER ME2 ;
 ANTENNAMAXAREACAR                       58.014 LAYER ME3 ;
 ANTENNAMAXAREACAR                       67.273 LAYER ME4 ;
END DI40
PIN DO39
  DIRECTION OUTPUT ;
 PORT
  LAYER ME4 ;
  RECT 876.400 0.000 877.200 1.000 ;
  LAYER ME3 ;
  RECT 876.400 0.000 877.200 1.000 ;
  LAYER ME2 ;
  RECT 876.400 0.000 877.200 1.000 ;
  LAYER ME1 ;
  RECT 876.400 0.000 877.200 1.000 ;
 END
 ANTENNAPARTIALMETALAREA                  4.160 LAYER ME2 ;
 ANTENNADIFFAREA                          5.472 LAYER ME2 ;
 ANTENNADIFFAREA                          5.472 LAYER ME3 ;
 ANTENNADIFFAREA                          5.472 LAYER ME4 ;
END DO39
PIN DI39
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 862.000 0.000 862.800 1.000 ;
  LAYER ME3 ;
  RECT 862.000 0.000 862.800 1.000 ;
  LAYER ME2 ;
  RECT 862.000 0.000 862.800 1.000 ;
  LAYER ME1 ;
  RECT 862.000 0.000 862.800 1.000 ;
 END
 ANTENNAPARTIALMETALAREA                  3.142 LAYER ME2 ;
 ANTENNAGATEAREA                          0.086 LAYER ME2 ;
 ANTENNAGATEAREA                          0.086 LAYER ME3 ;
 ANTENNAGATEAREA                          0.086 LAYER ME4 ;
 ANTENNADIFFAREA                          0.160 LAYER ME2 ;
 ANTENNADIFFAREA                          0.160 LAYER ME3 ;
 ANTENNADIFFAREA                          0.160 LAYER ME4 ;
 ANTENNAMAXAREACAR                       48.708 LAYER ME2 ;
 ANTENNAMAXAREACAR                       57.968 LAYER ME3 ;
 ANTENNAMAXAREACAR                       67.227 LAYER ME4 ;
END DI39
PIN DO38
  DIRECTION OUTPUT ;
 PORT
  LAYER ME4 ;
  RECT 856.800 0.000 857.600 1.000 ;
  LAYER ME3 ;
  RECT 856.800 0.000 857.600 1.000 ;
  LAYER ME2 ;
  RECT 856.800 0.000 857.600 1.000 ;
  LAYER ME1 ;
  RECT 856.800 0.000 857.600 1.000 ;
 END
 ANTENNAPARTIALMETALAREA                  4.168 LAYER ME2 ;
 ANTENNADIFFAREA                          5.472 LAYER ME2 ;
 ANTENNADIFFAREA                          5.472 LAYER ME3 ;
 ANTENNADIFFAREA                          5.472 LAYER ME4 ;
END DO38
PIN DI38
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 842.000 0.000 842.800 1.000 ;
  LAYER ME3 ;
  RECT 842.000 0.000 842.800 1.000 ;
  LAYER ME2 ;
  RECT 842.000 0.000 842.800 1.000 ;
  LAYER ME1 ;
  RECT 842.000 0.000 842.800 1.000 ;
 END
 ANTENNAPARTIALMETALAREA                  3.122 LAYER ME2 ;
 ANTENNAGATEAREA                          0.086 LAYER ME2 ;
 ANTENNAGATEAREA                          0.086 LAYER ME3 ;
 ANTENNAGATEAREA                          0.086 LAYER ME4 ;
 ANTENNADIFFAREA                          0.160 LAYER ME2 ;
 ANTENNADIFFAREA                          0.160 LAYER ME3 ;
 ANTENNADIFFAREA                          0.160 LAYER ME4 ;
 ANTENNAMAXAREACAR                       48.477 LAYER ME2 ;
 ANTENNAMAXAREACAR                       57.736 LAYER ME3 ;
 ANTENNAMAXAREACAR                       66.995 LAYER ME4 ;
END DI38
PIN DO37
  DIRECTION OUTPUT ;
 PORT
  LAYER ME4 ;
  RECT 835.600 0.000 836.400 1.000 ;
  LAYER ME3 ;
  RECT 835.600 0.000 836.400 1.000 ;
  LAYER ME2 ;
  RECT 835.600 0.000 836.400 1.000 ;
  LAYER ME1 ;
  RECT 835.600 0.000 836.400 1.000 ;
 END
 ANTENNAPARTIALMETALAREA                  4.144 LAYER ME2 ;
 ANTENNADIFFAREA                          5.472 LAYER ME2 ;
 ANTENNADIFFAREA                          5.472 LAYER ME3 ;
 ANTENNADIFFAREA                          5.472 LAYER ME4 ;
END DO37
PIN DI37
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 820.800 0.000 821.600 1.000 ;
  LAYER ME3 ;
  RECT 820.800 0.000 821.600 1.000 ;
  LAYER ME2 ;
  RECT 820.800 0.000 821.600 1.000 ;
  LAYER ME1 ;
  RECT 820.800 0.000 821.600 1.000 ;
 END
 ANTENNAPARTIALMETALAREA                  3.146 LAYER ME2 ;
 ANTENNAGATEAREA                          0.086 LAYER ME2 ;
 ANTENNAGATEAREA                          0.086 LAYER ME3 ;
 ANTENNAGATEAREA                          0.086 LAYER ME4 ;
 ANTENNADIFFAREA                          0.160 LAYER ME2 ;
 ANTENNADIFFAREA                          0.160 LAYER ME3 ;
 ANTENNADIFFAREA                          0.160 LAYER ME4 ;
 ANTENNAMAXAREACAR                       48.755 LAYER ME2 ;
 ANTENNAMAXAREACAR                       58.014 LAYER ME3 ;
 ANTENNAMAXAREACAR                       67.273 LAYER ME4 ;
END DI37
PIN DO36
  DIRECTION OUTPUT ;
 PORT
  LAYER ME4 ;
  RECT 815.600 0.000 816.400 1.000 ;
  LAYER ME3 ;
  RECT 815.600 0.000 816.400 1.000 ;
  LAYER ME2 ;
  RECT 815.600 0.000 816.400 1.000 ;
  LAYER ME1 ;
  RECT 815.600 0.000 816.400 1.000 ;
 END
 ANTENNAPARTIALMETALAREA                  4.168 LAYER ME2 ;
 ANTENNADIFFAREA                          5.472 LAYER ME2 ;
 ANTENNADIFFAREA                          5.472 LAYER ME3 ;
 ANTENNADIFFAREA                          5.472 LAYER ME4 ;
END DO36
PIN DI36
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 801.200 0.000 802.000 1.000 ;
  LAYER ME3 ;
  RECT 801.200 0.000 802.000 1.000 ;
  LAYER ME2 ;
  RECT 801.200 0.000 802.000 1.000 ;
  LAYER ME1 ;
  RECT 801.200 0.000 802.000 1.000 ;
 END
 ANTENNAPARTIALMETALAREA                  3.134 LAYER ME2 ;
 ANTENNAGATEAREA                          0.086 LAYER ME2 ;
 ANTENNAGATEAREA                          0.086 LAYER ME3 ;
 ANTENNAGATEAREA                          0.086 LAYER ME4 ;
 ANTENNADIFFAREA                          0.160 LAYER ME2 ;
 ANTENNADIFFAREA                          0.160 LAYER ME3 ;
 ANTENNADIFFAREA                          0.160 LAYER ME4 ;
 ANTENNAMAXAREACAR                       48.616 LAYER ME2 ;
 ANTENNAMAXAREACAR                       57.875 LAYER ME3 ;
 ANTENNAMAXAREACAR                       67.134 LAYER ME4 ;
END DI36
PIN DO35
  DIRECTION OUTPUT ;
 PORT
  LAYER ME4 ;
  RECT 794.800 0.000 795.600 1.000 ;
  LAYER ME3 ;
  RECT 794.800 0.000 795.600 1.000 ;
  LAYER ME2 ;
  RECT 794.800 0.000 795.600 1.000 ;
  LAYER ME1 ;
  RECT 794.800 0.000 795.600 1.000 ;
 END
 ANTENNAPARTIALMETALAREA                  4.168 LAYER ME2 ;
 ANTENNADIFFAREA                          5.472 LAYER ME2 ;
 ANTENNADIFFAREA                          5.472 LAYER ME3 ;
 ANTENNADIFFAREA                          5.472 LAYER ME4 ;
END DO35
PIN DI35
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 780.000 0.000 780.800 1.000 ;
  LAYER ME3 ;
  RECT 780.000 0.000 780.800 1.000 ;
  LAYER ME2 ;
  RECT 780.000 0.000 780.800 1.000 ;
  LAYER ME1 ;
  RECT 780.000 0.000 780.800 1.000 ;
 END
 ANTENNAPARTIALMETALAREA                  3.122 LAYER ME2 ;
 ANTENNAGATEAREA                          0.086 LAYER ME2 ;
 ANTENNAGATEAREA                          0.086 LAYER ME3 ;
 ANTENNAGATEAREA                          0.086 LAYER ME4 ;
 ANTENNADIFFAREA                          0.160 LAYER ME2 ;
 ANTENNADIFFAREA                          0.160 LAYER ME3 ;
 ANTENNADIFFAREA                          0.160 LAYER ME4 ;
 ANTENNAMAXAREACAR                       48.477 LAYER ME2 ;
 ANTENNAMAXAREACAR                       57.736 LAYER ME3 ;
 ANTENNAMAXAREACAR                       66.995 LAYER ME4 ;
END DI35
PIN DO34
  DIRECTION OUTPUT ;
 PORT
  LAYER ME4 ;
  RECT 774.800 0.000 775.600 1.000 ;
  LAYER ME3 ;
  RECT 774.800 0.000 775.600 1.000 ;
  LAYER ME2 ;
  RECT 774.800 0.000 775.600 1.000 ;
  LAYER ME1 ;
  RECT 774.800 0.000 775.600 1.000 ;
 END
 ANTENNAPARTIALMETALAREA                  4.144 LAYER ME2 ;
 ANTENNADIFFAREA                          5.472 LAYER ME2 ;
 ANTENNADIFFAREA                          5.472 LAYER ME3 ;
 ANTENNADIFFAREA                          5.472 LAYER ME4 ;
END DO34
PIN DI34
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 760.000 0.000 760.800 1.000 ;
  LAYER ME3 ;
  RECT 760.000 0.000 760.800 1.000 ;
  LAYER ME2 ;
  RECT 760.000 0.000 760.800 1.000 ;
  LAYER ME1 ;
  RECT 760.000 0.000 760.800 1.000 ;
 END
 ANTENNAPARTIALMETALAREA                  3.154 LAYER ME2 ;
 ANTENNAGATEAREA                          0.086 LAYER ME2 ;
 ANTENNAGATEAREA                          0.086 LAYER ME3 ;
 ANTENNAGATEAREA                          0.086 LAYER ME4 ;
 ANTENNADIFFAREA                          0.160 LAYER ME2 ;
 ANTENNADIFFAREA                          0.160 LAYER ME3 ;
 ANTENNADIFFAREA                          0.160 LAYER ME4 ;
 ANTENNAMAXAREACAR                       48.847 LAYER ME2 ;
 ANTENNAMAXAREACAR                       58.106 LAYER ME3 ;
 ANTENNAMAXAREACAR                       67.366 LAYER ME4 ;
END DI34
PIN DO33
  DIRECTION OUTPUT ;
 PORT
  LAYER ME4 ;
  RECT 753.600 0.000 754.400 1.000 ;
  LAYER ME3 ;
  RECT 753.600 0.000 754.400 1.000 ;
  LAYER ME2 ;
  RECT 753.600 0.000 754.400 1.000 ;
  LAYER ME1 ;
  RECT 753.600 0.000 754.400 1.000 ;
 END
 ANTENNAPARTIALMETALAREA                  4.168 LAYER ME2 ;
 ANTENNADIFFAREA                          5.472 LAYER ME2 ;
 ANTENNADIFFAREA                          5.472 LAYER ME3 ;
 ANTENNADIFFAREA                          5.472 LAYER ME4 ;
END DO33
PIN DI33
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 739.200 0.000 740.000 1.000 ;
  LAYER ME3 ;
  RECT 739.200 0.000 740.000 1.000 ;
  LAYER ME2 ;
  RECT 739.200 0.000 740.000 1.000 ;
  LAYER ME1 ;
  RECT 739.200 0.000 740.000 1.000 ;
 END
 ANTENNAPARTIALMETALAREA                  3.134 LAYER ME2 ;
 ANTENNAGATEAREA                          0.086 LAYER ME2 ;
 ANTENNAGATEAREA                          0.086 LAYER ME3 ;
 ANTENNAGATEAREA                          0.086 LAYER ME4 ;
 ANTENNADIFFAREA                          0.160 LAYER ME2 ;
 ANTENNADIFFAREA                          0.160 LAYER ME3 ;
 ANTENNADIFFAREA                          0.160 LAYER ME4 ;
 ANTENNAMAXAREACAR                       48.616 LAYER ME2 ;
 ANTENNAMAXAREACAR                       57.875 LAYER ME3 ;
 ANTENNAMAXAREACAR                       67.134 LAYER ME4 ;
END DI33
PIN DO32
  DIRECTION OUTPUT ;
 PORT
  LAYER ME4 ;
  RECT 734.000 0.000 734.800 1.000 ;
  LAYER ME3 ;
  RECT 734.000 0.000 734.800 1.000 ;
  LAYER ME2 ;
  RECT 734.000 0.000 734.800 1.000 ;
  LAYER ME1 ;
  RECT 734.000 0.000 734.800 1.000 ;
 END
 ANTENNAPARTIALMETALAREA                  4.160 LAYER ME2 ;
 ANTENNADIFFAREA                          5.472 LAYER ME2 ;
 ANTENNADIFFAREA                          5.472 LAYER ME3 ;
 ANTENNADIFFAREA                          5.472 LAYER ME4 ;
END DO32
PIN WEB4
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 720.800 0.000 721.600 1.000 ;
  LAYER ME3 ;
  RECT 720.800 0.000 721.600 1.000 ;
  LAYER ME2 ;
  RECT 720.800 0.000 721.600 1.000 ;
  LAYER ME1 ;
  RECT 720.800 0.000 721.600 1.000 ;
 END
 ANTENNAPARTIALMETALAREA                  2.868 LAYER ME2 ;
 ANTENNAGATEAREA                          0.072 LAYER ME2 ;
 ANTENNAGATEAREA                          0.072 LAYER ME3 ;
 ANTENNAGATEAREA                          0.072 LAYER ME4 ;
 ANTENNADIFFAREA                          0.160 LAYER ME2 ;
 ANTENNADIFFAREA                          0.160 LAYER ME3 ;
 ANTENNADIFFAREA                          0.160 LAYER ME4 ;
 ANTENNAMAXAREACAR                       54.844 LAYER ME2 ;
 ANTENNAMAXAREACAR                       65.956 LAYER ME3 ;
 ANTENNAMAXAREACAR                       77.067 LAYER ME4 ;
END WEB4
PIN DI32
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 719.200 0.000 720.000 1.000 ;
  LAYER ME3 ;
  RECT 719.200 0.000 720.000 1.000 ;
  LAYER ME2 ;
  RECT 719.200 0.000 720.000 1.000 ;
  LAYER ME1 ;
  RECT 719.200 0.000 720.000 1.000 ;
 END
 ANTENNAPARTIALMETALAREA                  3.130 LAYER ME2 ;
 ANTENNAGATEAREA                          0.086 LAYER ME2 ;
 ANTENNAGATEAREA                          0.086 LAYER ME3 ;
 ANTENNAGATEAREA                          0.086 LAYER ME4 ;
 ANTENNADIFFAREA                          0.160 LAYER ME2 ;
 ANTENNADIFFAREA                          0.160 LAYER ME3 ;
 ANTENNADIFFAREA                          0.160 LAYER ME4 ;
 ANTENNAMAXAREACAR                       48.569 LAYER ME2 ;
 ANTENNAMAXAREACAR                       57.829 LAYER ME3 ;
 ANTENNAMAXAREACAR                       67.088 LAYER ME4 ;
END DI32
PIN A3
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 698.400 0.000 699.200 1.000 ;
  LAYER ME3 ;
  RECT 698.400 0.000 699.200 1.000 ;
  LAYER ME2 ;
  RECT 698.400 0.000 699.200 1.000 ;
  LAYER ME1 ;
  RECT 698.400 0.000 699.200 1.000 ;
 END
 ANTENNAPARTIALMETALAREA                  2.044 LAYER ME2 ;
 ANTENNAGATEAREA                          0.180 LAYER ME2 ;
 ANTENNAGATEAREA                          0.180 LAYER ME3 ;
 ANTENNAGATEAREA                          0.180 LAYER ME4 ;
 ANTENNADIFFAREA                          0.160 LAYER ME2 ;
 ANTENNADIFFAREA                          0.160 LAYER ME3 ;
 ANTENNADIFFAREA                          0.160 LAYER ME4 ;
 ANTENNAMAXAREACAR                       17.204 LAYER ME2 ;
 ANTENNAMAXAREACAR                       21.649 LAYER ME3 ;
 ANTENNAMAXAREACAR                       26.093 LAYER ME4 ;
END A3
PIN A1
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 697.200 0.000 698.000 1.000 ;
  LAYER ME3 ;
  RECT 697.200 0.000 698.000 1.000 ;
  LAYER ME2 ;
  RECT 697.200 0.000 698.000 1.000 ;
  LAYER ME1 ;
  RECT 697.200 0.000 698.000 1.000 ;
 END
 ANTENNAPARTIALMETALAREA                  7.314 LAYER ME2 ;
 ANTENNAGATEAREA                          0.192 LAYER ME2 ;
 ANTENNAGATEAREA                          0.192 LAYER ME3 ;
 ANTENNAGATEAREA                          0.192 LAYER ME4 ;
 ANTENNADIFFAREA                          0.160 LAYER ME2 ;
 ANTENNADIFFAREA                          0.160 LAYER ME3 ;
 ANTENNADIFFAREA                          0.160 LAYER ME4 ;
 ANTENNAMAXAREACAR                       43.535 LAYER ME2 ;
 ANTENNAMAXAREACAR                       47.702 LAYER ME3 ;
 ANTENNAMAXAREACAR                       51.869 LAYER ME4 ;
END A1
PIN OE
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 696.000 0.000 696.800 1.000 ;
  LAYER ME3 ;
  RECT 696.000 0.000 696.800 1.000 ;
  LAYER ME2 ;
  RECT 696.000 0.000 696.800 1.000 ;
  LAYER ME1 ;
  RECT 696.000 0.000 696.800 1.000 ;
 END
 ANTENNAPARTIALMETALAREA                  3.386 LAYER ME2 ;
 ANTENNAGATEAREA                          0.840 LAYER ME2 ;
 ANTENNAGATEAREA                          0.840 LAYER ME3 ;
 ANTENNAGATEAREA                          0.840 LAYER ME4 ;
 ANTENNADIFFAREA                          0.160 LAYER ME2 ;
 ANTENNADIFFAREA                          0.160 LAYER ME3 ;
 ANTENNADIFFAREA                          0.160 LAYER ME4 ;
 ANTENNAMAXAREACAR                        5.355 LAYER ME2 ;
 ANTENNAMAXAREACAR                        6.307 LAYER ME3 ;
 ANTENNAMAXAREACAR                        7.260 LAYER ME4 ;
END OE
PIN CS
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 694.800 0.000 695.600 1.000 ;
  LAYER ME3 ;
  RECT 694.800 0.000 695.600 1.000 ;
  LAYER ME2 ;
  RECT 694.800 0.000 695.600 1.000 ;
  LAYER ME1 ;
  RECT 694.800 0.000 695.600 1.000 ;
 END
 ANTENNAPARTIALMETALAREA                  5.092 LAYER ME2 ;
 ANTENNAGATEAREA                          1.680 LAYER ME2 ;
 ANTENNAGATEAREA                          1.680 LAYER ME3 ;
 ANTENNAGATEAREA                          1.680 LAYER ME4 ;
 ANTENNADIFFAREA                          0.160 LAYER ME2 ;
 ANTENNADIFFAREA                          0.160 LAYER ME3 ;
 ANTENNADIFFAREA                          0.160 LAYER ME4 ;
 ANTENNAMAXAREACAR                        3.658 LAYER ME2 ;
 ANTENNAMAXAREACAR                        4.134 LAYER ME3 ;
 ANTENNAMAXAREACAR                        4.610 LAYER ME4 ;
END CS
PIN A2
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 693.600 0.000 694.400 1.000 ;
  LAYER ME3 ;
  RECT 693.600 0.000 694.400 1.000 ;
  LAYER ME2 ;
  RECT 693.600 0.000 694.400 1.000 ;
  LAYER ME1 ;
  RECT 693.600 0.000 694.400 1.000 ;
 END
 ANTENNAPARTIALMETALAREA                  7.382 LAYER ME2 ;
 ANTENNAGATEAREA                          0.192 LAYER ME2 ;
 ANTENNAGATEAREA                          0.192 LAYER ME3 ;
 ANTENNAGATEAREA                          0.192 LAYER ME4 ;
 ANTENNADIFFAREA                          0.160 LAYER ME2 ;
 ANTENNADIFFAREA                          0.160 LAYER ME3 ;
 ANTENNADIFFAREA                          0.160 LAYER ME4 ;
 ANTENNAMAXAREACAR                       43.890 LAYER ME2 ;
 ANTENNAMAXAREACAR                       48.056 LAYER ME3 ;
 ANTENNAMAXAREACAR                       52.223 LAYER ME4 ;
END A2
PIN A0
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 692.400 0.000 693.200 1.000 ;
  LAYER ME3 ;
  RECT 692.400 0.000 693.200 1.000 ;
  LAYER ME2 ;
  RECT 692.400 0.000 693.200 1.000 ;
  LAYER ME1 ;
  RECT 692.400 0.000 693.200 1.000 ;
 END
 ANTENNAPARTIALMETALAREA                  7.414 LAYER ME2 ;
 ANTENNAGATEAREA                          0.192 LAYER ME2 ;
 ANTENNAGATEAREA                          0.192 LAYER ME3 ;
 ANTENNAGATEAREA                          0.192 LAYER ME4 ;
 ANTENNADIFFAREA                          0.160 LAYER ME2 ;
 ANTENNADIFFAREA                          0.160 LAYER ME3 ;
 ANTENNADIFFAREA                          0.160 LAYER ME4 ;
 ANTENNAMAXAREACAR                       44.056 LAYER ME2 ;
 ANTENNAMAXAREACAR                       48.223 LAYER ME3 ;
 ANTENNAMAXAREACAR                       52.390 LAYER ME4 ;
END A0
PIN CK
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 686.400 0.000 687.200 1.000 ;
  LAYER ME3 ;
  RECT 686.400 0.000 687.200 1.000 ;
  LAYER ME2 ;
  RECT 686.400 0.000 687.200 1.000 ;
  LAYER ME1 ;
  RECT 686.400 0.000 687.200 1.000 ;
 END
 ANTENNAPARTIALMETALAREA                  5.514 LAYER ME2 ;
 ANTENNAGATEAREA                          1.908 LAYER ME2 ;
 ANTENNAGATEAREA                          1.908 LAYER ME3 ;
 ANTENNAGATEAREA                          1.908 LAYER ME4 ;
 ANTENNADIFFAREA                          0.160 LAYER ME2 ;
 ANTENNADIFFAREA                          0.160 LAYER ME3 ;
 ANTENNADIFFAREA                          0.160 LAYER ME4 ;
 ANTENNAMAXAREACAR                       59.411 LAYER ME2 ;
 ANTENNAMAXAREACAR                       66.819 LAYER ME3 ;
 ANTENNAMAXAREACAR                       74.226 LAYER ME4 ;
END CK
PIN A4
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 679.200 0.000 680.000 1.000 ;
  LAYER ME3 ;
  RECT 679.200 0.000 680.000 1.000 ;
  LAYER ME2 ;
  RECT 679.200 0.000 680.000 1.000 ;
  LAYER ME1 ;
  RECT 679.200 0.000 680.000 1.000 ;
 END
 ANTENNAPARTIALMETALAREA                  2.196 LAYER ME2 ;
 ANTENNAGATEAREA                          0.180 LAYER ME2 ;
 ANTENNAGATEAREA                          0.180 LAYER ME3 ;
 ANTENNAGATEAREA                          0.180 LAYER ME4 ;
 ANTENNADIFFAREA                          0.160 LAYER ME2 ;
 ANTENNADIFFAREA                          0.160 LAYER ME3 ;
 ANTENNADIFFAREA                          0.160 LAYER ME4 ;
 ANTENNAMAXAREACAR                       18.092 LAYER ME2 ;
 ANTENNAMAXAREACAR                       22.537 LAYER ME3 ;
 ANTENNAMAXAREACAR                       26.981 LAYER ME4 ;
END A4
PIN A5
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 676.800 0.000 677.600 1.000 ;
  LAYER ME3 ;
  RECT 676.800 0.000 677.600 1.000 ;
  LAYER ME2 ;
  RECT 676.800 0.000 677.600 1.000 ;
  LAYER ME1 ;
  RECT 676.800 0.000 677.600 1.000 ;
 END
 ANTENNAPARTIALMETALAREA                  2.390 LAYER ME2 ;
 ANTENNAGATEAREA                          0.180 LAYER ME2 ;
 ANTENNAGATEAREA                          0.180 LAYER ME3 ;
 ANTENNAGATEAREA                          0.180 LAYER ME4 ;
 ANTENNADIFFAREA                          0.160 LAYER ME2 ;
 ANTENNADIFFAREA                          0.160 LAYER ME3 ;
 ANTENNADIFFAREA                          0.160 LAYER ME4 ;
 ANTENNAMAXAREACAR                       19.230 LAYER ME2 ;
 ANTENNAMAXAREACAR                       23.674 LAYER ME3 ;
 ANTENNAMAXAREACAR                       28.119 LAYER ME4 ;
END A5
PIN A6
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 674.000 0.000 674.800 1.000 ;
  LAYER ME3 ;
  RECT 674.000 0.000 674.800 1.000 ;
  LAYER ME2 ;
  RECT 674.000 0.000 674.800 1.000 ;
  LAYER ME1 ;
  RECT 674.000 0.000 674.800 1.000 ;
 END
 ANTENNAPARTIALMETALAREA                  2.402 LAYER ME2 ;
 ANTENNAGATEAREA                          0.180 LAYER ME2 ;
 ANTENNAGATEAREA                          0.180 LAYER ME3 ;
 ANTENNAGATEAREA                          0.180 LAYER ME4 ;
 ANTENNADIFFAREA                          0.160 LAYER ME2 ;
 ANTENNADIFFAREA                          0.160 LAYER ME3 ;
 ANTENNADIFFAREA                          0.160 LAYER ME4 ;
 ANTENNAMAXAREACAR                       19.200 LAYER ME2 ;
 ANTENNAMAXAREACAR                       23.644 LAYER ME3 ;
 ANTENNAMAXAREACAR                       28.089 LAYER ME4 ;
END A6
PIN A7
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 671.200 0.000 672.000 1.000 ;
  LAYER ME3 ;
  RECT 671.200 0.000 672.000 1.000 ;
  LAYER ME2 ;
  RECT 671.200 0.000 672.000 1.000 ;
  LAYER ME1 ;
  RECT 671.200 0.000 672.000 1.000 ;
 END
 ANTENNAPARTIALMETALAREA                  2.394 LAYER ME2 ;
 ANTENNAGATEAREA                          0.180 LAYER ME2 ;
 ANTENNAGATEAREA                          0.180 LAYER ME3 ;
 ANTENNAGATEAREA                          0.180 LAYER ME4 ;
 ANTENNADIFFAREA                          0.160 LAYER ME2 ;
 ANTENNADIFFAREA                          0.160 LAYER ME3 ;
 ANTENNADIFFAREA                          0.160 LAYER ME4 ;
 ANTENNAMAXAREACAR                       19.156 LAYER ME2 ;
 ANTENNAMAXAREACAR                       23.600 LAYER ME3 ;
 ANTENNAMAXAREACAR                       28.044 LAYER ME4 ;
END A7
PIN A8
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 670.000 0.000 670.800 1.000 ;
  LAYER ME3 ;
  RECT 670.000 0.000 670.800 1.000 ;
  LAYER ME2 ;
  RECT 670.000 0.000 670.800 1.000 ;
  LAYER ME1 ;
  RECT 670.000 0.000 670.800 1.000 ;
 END
 ANTENNAPARTIALMETALAREA                  2.402 LAYER ME2 ;
 ANTENNAGATEAREA                          0.180 LAYER ME2 ;
 ANTENNAGATEAREA                          0.180 LAYER ME3 ;
 ANTENNAGATEAREA                          0.180 LAYER ME4 ;
 ANTENNADIFFAREA                          0.160 LAYER ME2 ;
 ANTENNADIFFAREA                          0.160 LAYER ME3 ;
 ANTENNADIFFAREA                          0.160 LAYER ME4 ;
 ANTENNAMAXAREACAR                       19.200 LAYER ME2 ;
 ANTENNAMAXAREACAR                       23.644 LAYER ME3 ;
 ANTENNAMAXAREACAR                       28.089 LAYER ME4 ;
END A8
PIN A9
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 667.200 0.000 668.000 1.000 ;
  LAYER ME3 ;
  RECT 667.200 0.000 668.000 1.000 ;
  LAYER ME2 ;
  RECT 667.200 0.000 668.000 1.000 ;
  LAYER ME1 ;
  RECT 667.200 0.000 668.000 1.000 ;
 END
 ANTENNAPARTIALMETALAREA                  2.394 LAYER ME2 ;
 ANTENNAGATEAREA                          0.180 LAYER ME2 ;
 ANTENNAGATEAREA                          0.180 LAYER ME3 ;
 ANTENNAGATEAREA                          0.180 LAYER ME4 ;
 ANTENNADIFFAREA                          0.160 LAYER ME2 ;
 ANTENNADIFFAREA                          0.160 LAYER ME3 ;
 ANTENNADIFFAREA                          0.160 LAYER ME4 ;
 ANTENNAMAXAREACAR                       19.156 LAYER ME2 ;
 ANTENNAMAXAREACAR                       23.600 LAYER ME3 ;
 ANTENNAMAXAREACAR                       28.044 LAYER ME4 ;
END A9
PIN A10
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 666.000 0.000 666.800 1.000 ;
  LAYER ME3 ;
  RECT 666.000 0.000 666.800 1.000 ;
  LAYER ME2 ;
  RECT 666.000 0.000 666.800 1.000 ;
  LAYER ME1 ;
  RECT 666.000 0.000 666.800 1.000 ;
 END
 ANTENNAPARTIALMETALAREA                  2.402 LAYER ME2 ;
 ANTENNAGATEAREA                          0.180 LAYER ME2 ;
 ANTENNAGATEAREA                          0.180 LAYER ME3 ;
 ANTENNAGATEAREA                          0.180 LAYER ME4 ;
 ANTENNADIFFAREA                          0.160 LAYER ME2 ;
 ANTENNADIFFAREA                          0.160 LAYER ME3 ;
 ANTENNADIFFAREA                          0.160 LAYER ME4 ;
 ANTENNAMAXAREACAR                       19.200 LAYER ME2 ;
 ANTENNAMAXAREACAR                       23.644 LAYER ME3 ;
 ANTENNAMAXAREACAR                       28.089 LAYER ME4 ;
END A10
PIN A11
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 663.200 0.000 664.000 1.000 ;
  LAYER ME3 ;
  RECT 663.200 0.000 664.000 1.000 ;
  LAYER ME2 ;
  RECT 663.200 0.000 664.000 1.000 ;
  LAYER ME1 ;
  RECT 663.200 0.000 664.000 1.000 ;
 END
 ANTENNAPARTIALMETALAREA                  2.394 LAYER ME2 ;
 ANTENNAGATEAREA                          0.180 LAYER ME2 ;
 ANTENNAGATEAREA                          0.180 LAYER ME3 ;
 ANTENNAGATEAREA                          0.180 LAYER ME4 ;
 ANTENNADIFFAREA                          0.160 LAYER ME2 ;
 ANTENNADIFFAREA                          0.160 LAYER ME3 ;
 ANTENNADIFFAREA                          0.160 LAYER ME4 ;
 ANTENNAMAXAREACAR                       19.156 LAYER ME2 ;
 ANTENNAMAXAREACAR                       23.600 LAYER ME3 ;
 ANTENNAMAXAREACAR                       28.044 LAYER ME4 ;
END A11
PIN DO31
  DIRECTION OUTPUT ;
 PORT
  LAYER ME4 ;
  RECT 656.400 0.000 657.200 1.000 ;
  LAYER ME3 ;
  RECT 656.400 0.000 657.200 1.000 ;
  LAYER ME2 ;
  RECT 656.400 0.000 657.200 1.000 ;
  LAYER ME1 ;
  RECT 656.400 0.000 657.200 1.000 ;
 END
 ANTENNAPARTIALMETALAREA                  4.148 LAYER ME2 ;
 ANTENNADIFFAREA                          5.472 LAYER ME2 ;
 ANTENNADIFFAREA                          5.472 LAYER ME3 ;
 ANTENNADIFFAREA                          5.472 LAYER ME4 ;
END DO31
PIN DI31
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 642.000 0.000 642.800 1.000 ;
  LAYER ME3 ;
  RECT 642.000 0.000 642.800 1.000 ;
  LAYER ME2 ;
  RECT 642.000 0.000 642.800 1.000 ;
  LAYER ME1 ;
  RECT 642.000 0.000 642.800 1.000 ;
 END
 ANTENNAPARTIALMETALAREA                  3.154 LAYER ME2 ;
 ANTENNAGATEAREA                          0.086 LAYER ME2 ;
 ANTENNAGATEAREA                          0.086 LAYER ME3 ;
 ANTENNAGATEAREA                          0.086 LAYER ME4 ;
 ANTENNADIFFAREA                          0.160 LAYER ME2 ;
 ANTENNADIFFAREA                          0.160 LAYER ME3 ;
 ANTENNADIFFAREA                          0.160 LAYER ME4 ;
 ANTENNAMAXAREACAR                       48.847 LAYER ME2 ;
 ANTENNAMAXAREACAR                       58.106 LAYER ME3 ;
 ANTENNAMAXAREACAR                       67.366 LAYER ME4 ;
END DI31
PIN DO30
  DIRECTION OUTPUT ;
 PORT
  LAYER ME4 ;
  RECT 636.400 0.000 637.200 1.000 ;
  LAYER ME3 ;
  RECT 636.400 0.000 637.200 1.000 ;
  LAYER ME2 ;
  RECT 636.400 0.000 637.200 1.000 ;
  LAYER ME1 ;
  RECT 636.400 0.000 637.200 1.000 ;
 END
 ANTENNAPARTIALMETALAREA                  4.180 LAYER ME2 ;
 ANTENNADIFFAREA                          5.472 LAYER ME2 ;
 ANTENNADIFFAREA                          5.472 LAYER ME3 ;
 ANTENNADIFFAREA                          5.472 LAYER ME4 ;
END DO30
PIN DI30
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 622.000 0.000 622.800 1.000 ;
  LAYER ME3 ;
  RECT 622.000 0.000 622.800 1.000 ;
  LAYER ME2 ;
  RECT 622.000 0.000 622.800 1.000 ;
  LAYER ME1 ;
  RECT 622.000 0.000 622.800 1.000 ;
 END
 ANTENNAPARTIALMETALAREA                  3.122 LAYER ME2 ;
 ANTENNAGATEAREA                          0.086 LAYER ME2 ;
 ANTENNAGATEAREA                          0.086 LAYER ME3 ;
 ANTENNAGATEAREA                          0.086 LAYER ME4 ;
 ANTENNADIFFAREA                          0.160 LAYER ME2 ;
 ANTENNADIFFAREA                          0.160 LAYER ME3 ;
 ANTENNADIFFAREA                          0.160 LAYER ME4 ;
 ANTENNAMAXAREACAR                       48.477 LAYER ME2 ;
 ANTENNAMAXAREACAR                       57.736 LAYER ME3 ;
 ANTENNAMAXAREACAR                       66.995 LAYER ME4 ;
END DI30
PIN DO29
  DIRECTION OUTPUT ;
 PORT
  LAYER ME4 ;
  RECT 615.600 0.000 616.400 1.000 ;
  LAYER ME3 ;
  RECT 615.600 0.000 616.400 1.000 ;
  LAYER ME2 ;
  RECT 615.600 0.000 616.400 1.000 ;
  LAYER ME1 ;
  RECT 615.600 0.000 616.400 1.000 ;
 END
 ANTENNAPARTIALMETALAREA                  4.156 LAYER ME2 ;
 ANTENNADIFFAREA                          5.472 LAYER ME2 ;
 ANTENNADIFFAREA                          5.472 LAYER ME3 ;
 ANTENNADIFFAREA                          5.472 LAYER ME4 ;
END DO29
PIN DI29
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 600.800 0.000 601.600 1.000 ;
  LAYER ME3 ;
  RECT 600.800 0.000 601.600 1.000 ;
  LAYER ME2 ;
  RECT 600.800 0.000 601.600 1.000 ;
  LAYER ME1 ;
  RECT 600.800 0.000 601.600 1.000 ;
 END
 ANTENNAPARTIALMETALAREA                  3.134 LAYER ME2 ;
 ANTENNAGATEAREA                          0.086 LAYER ME2 ;
 ANTENNAGATEAREA                          0.086 LAYER ME3 ;
 ANTENNAGATEAREA                          0.086 LAYER ME4 ;
 ANTENNADIFFAREA                          0.160 LAYER ME2 ;
 ANTENNADIFFAREA                          0.160 LAYER ME3 ;
 ANTENNADIFFAREA                          0.160 LAYER ME4 ;
 ANTENNAMAXAREACAR                       48.616 LAYER ME2 ;
 ANTENNAMAXAREACAR                       57.875 LAYER ME3 ;
 ANTENNAMAXAREACAR                       67.134 LAYER ME4 ;
END DI29
PIN DO28
  DIRECTION OUTPUT ;
 PORT
  LAYER ME4 ;
  RECT 595.600 0.000 596.400 1.000 ;
  LAYER ME3 ;
  RECT 595.600 0.000 596.400 1.000 ;
  LAYER ME2 ;
  RECT 595.600 0.000 596.400 1.000 ;
  LAYER ME1 ;
  RECT 595.600 0.000 596.400 1.000 ;
 END
 ANTENNAPARTIALMETALAREA                  4.156 LAYER ME2 ;
 ANTENNADIFFAREA                          5.472 LAYER ME2 ;
 ANTENNADIFFAREA                          5.472 LAYER ME3 ;
 ANTENNADIFFAREA                          5.472 LAYER ME4 ;
END DO28
PIN DI28
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 581.200 0.000 582.000 1.000 ;
  LAYER ME3 ;
  RECT 581.200 0.000 582.000 1.000 ;
  LAYER ME2 ;
  RECT 581.200 0.000 582.000 1.000 ;
  LAYER ME1 ;
  RECT 581.200 0.000 582.000 1.000 ;
 END
 ANTENNAPARTIALMETALAREA                  3.146 LAYER ME2 ;
 ANTENNAGATEAREA                          0.086 LAYER ME2 ;
 ANTENNAGATEAREA                          0.086 LAYER ME3 ;
 ANTENNAGATEAREA                          0.086 LAYER ME4 ;
 ANTENNADIFFAREA                          0.160 LAYER ME2 ;
 ANTENNADIFFAREA                          0.160 LAYER ME3 ;
 ANTENNADIFFAREA                          0.160 LAYER ME4 ;
 ANTENNAMAXAREACAR                       48.755 LAYER ME2 ;
 ANTENNAMAXAREACAR                       58.014 LAYER ME3 ;
 ANTENNAMAXAREACAR                       67.273 LAYER ME4 ;
END DI28
PIN DO27
  DIRECTION OUTPUT ;
 PORT
  LAYER ME4 ;
  RECT 574.400 0.000 575.200 1.000 ;
  LAYER ME3 ;
  RECT 574.400 0.000 575.200 1.000 ;
  LAYER ME2 ;
  RECT 574.400 0.000 575.200 1.000 ;
  LAYER ME1 ;
  RECT 574.400 0.000 575.200 1.000 ;
 END
 ANTENNAPARTIALMETALAREA                  4.180 LAYER ME2 ;
 ANTENNADIFFAREA                          5.472 LAYER ME2 ;
 ANTENNADIFFAREA                          5.472 LAYER ME3 ;
 ANTENNADIFFAREA                          5.472 LAYER ME4 ;
END DO27
PIN DI27
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 560.000 0.000 560.800 1.000 ;
  LAYER ME3 ;
  RECT 560.000 0.000 560.800 1.000 ;
  LAYER ME2 ;
  RECT 560.000 0.000 560.800 1.000 ;
  LAYER ME1 ;
  RECT 560.000 0.000 560.800 1.000 ;
 END
 ANTENNAPARTIALMETALAREA                  3.122 LAYER ME2 ;
 ANTENNAGATEAREA                          0.086 LAYER ME2 ;
 ANTENNAGATEAREA                          0.086 LAYER ME3 ;
 ANTENNAGATEAREA                          0.086 LAYER ME4 ;
 ANTENNADIFFAREA                          0.160 LAYER ME2 ;
 ANTENNADIFFAREA                          0.160 LAYER ME3 ;
 ANTENNADIFFAREA                          0.160 LAYER ME4 ;
 ANTENNAMAXAREACAR                       48.477 LAYER ME2 ;
 ANTENNAMAXAREACAR                       57.736 LAYER ME3 ;
 ANTENNAMAXAREACAR                       66.995 LAYER ME4 ;
END DI27
PIN DO26
  DIRECTION OUTPUT ;
 PORT
  LAYER ME4 ;
  RECT 554.800 0.000 555.600 1.000 ;
  LAYER ME3 ;
  RECT 554.800 0.000 555.600 1.000 ;
  LAYER ME2 ;
  RECT 554.800 0.000 555.600 1.000 ;
  LAYER ME1 ;
  RECT 554.800 0.000 555.600 1.000 ;
 END
 ANTENNAPARTIALMETALAREA                  4.148 LAYER ME2 ;
 ANTENNADIFFAREA                          5.472 LAYER ME2 ;
 ANTENNADIFFAREA                          5.472 LAYER ME3 ;
 ANTENNADIFFAREA                          5.472 LAYER ME4 ;
END DO26
PIN DI26
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 540.000 0.000 540.800 1.000 ;
  LAYER ME3 ;
  RECT 540.000 0.000 540.800 1.000 ;
  LAYER ME2 ;
  RECT 540.000 0.000 540.800 1.000 ;
  LAYER ME1 ;
  RECT 540.000 0.000 540.800 1.000 ;
 END
 ANTENNAPARTIALMETALAREA                  3.142 LAYER ME2 ;
 ANTENNAGATEAREA                          0.086 LAYER ME2 ;
 ANTENNAGATEAREA                          0.086 LAYER ME3 ;
 ANTENNAGATEAREA                          0.086 LAYER ME4 ;
 ANTENNADIFFAREA                          0.160 LAYER ME2 ;
 ANTENNADIFFAREA                          0.160 LAYER ME3 ;
 ANTENNADIFFAREA                          0.160 LAYER ME4 ;
 ANTENNAMAXAREACAR                       48.708 LAYER ME2 ;
 ANTENNAMAXAREACAR                       57.968 LAYER ME3 ;
 ANTENNAMAXAREACAR                       67.227 LAYER ME4 ;
END DI26
PIN DO25
  DIRECTION OUTPUT ;
 PORT
  LAYER ME4 ;
  RECT 533.600 0.000 534.400 1.000 ;
  LAYER ME3 ;
  RECT 533.600 0.000 534.400 1.000 ;
  LAYER ME2 ;
  RECT 533.600 0.000 534.400 1.000 ;
  LAYER ME1 ;
  RECT 533.600 0.000 534.400 1.000 ;
 END
 ANTENNAPARTIALMETALAREA                  4.156 LAYER ME2 ;
 ANTENNADIFFAREA                          5.472 LAYER ME2 ;
 ANTENNADIFFAREA                          5.472 LAYER ME3 ;
 ANTENNADIFFAREA                          5.472 LAYER ME4 ;
END DO25
PIN DI25
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 519.200 0.000 520.000 1.000 ;
  LAYER ME3 ;
  RECT 519.200 0.000 520.000 1.000 ;
  LAYER ME2 ;
  RECT 519.200 0.000 520.000 1.000 ;
  LAYER ME1 ;
  RECT 519.200 0.000 520.000 1.000 ;
 END
 ANTENNAPARTIALMETALAREA                  3.146 LAYER ME2 ;
 ANTENNAGATEAREA                          0.086 LAYER ME2 ;
 ANTENNAGATEAREA                          0.086 LAYER ME3 ;
 ANTENNAGATEAREA                          0.086 LAYER ME4 ;
 ANTENNADIFFAREA                          0.160 LAYER ME2 ;
 ANTENNADIFFAREA                          0.160 LAYER ME3 ;
 ANTENNADIFFAREA                          0.160 LAYER ME4 ;
 ANTENNAMAXAREACAR                       48.755 LAYER ME2 ;
 ANTENNAMAXAREACAR                       58.014 LAYER ME3 ;
 ANTENNAMAXAREACAR                       67.273 LAYER ME4 ;
END DI25
PIN DO24
  DIRECTION OUTPUT ;
 PORT
  LAYER ME4 ;
  RECT 514.000 0.000 514.800 1.000 ;
  LAYER ME3 ;
  RECT 514.000 0.000 514.800 1.000 ;
  LAYER ME2 ;
  RECT 514.000 0.000 514.800 1.000 ;
  LAYER ME1 ;
  RECT 514.000 0.000 514.800 1.000 ;
 END
 ANTENNAPARTIALMETALAREA                  4.172 LAYER ME2 ;
 ANTENNADIFFAREA                          5.472 LAYER ME2 ;
 ANTENNADIFFAREA                          5.472 LAYER ME3 ;
 ANTENNADIFFAREA                          5.472 LAYER ME4 ;
END DO24
PIN WEB3
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 500.800 0.000 501.600 1.000 ;
  LAYER ME3 ;
  RECT 500.800 0.000 501.600 1.000 ;
  LAYER ME2 ;
  RECT 500.800 0.000 501.600 1.000 ;
  LAYER ME1 ;
  RECT 500.800 0.000 501.600 1.000 ;
 END
 ANTENNAPARTIALMETALAREA                  2.856 LAYER ME2 ;
 ANTENNAGATEAREA                          0.072 LAYER ME2 ;
 ANTENNAGATEAREA                          0.072 LAYER ME3 ;
 ANTENNAGATEAREA                          0.072 LAYER ME4 ;
 ANTENNADIFFAREA                          0.160 LAYER ME2 ;
 ANTENNADIFFAREA                          0.160 LAYER ME3 ;
 ANTENNADIFFAREA                          0.160 LAYER ME4 ;
 ANTENNAMAXAREACAR                       54.678 LAYER ME2 ;
 ANTENNAMAXAREACAR                       65.789 LAYER ME3 ;
 ANTENNAMAXAREACAR                       76.900 LAYER ME4 ;
END WEB3
PIN DI24
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 499.200 0.000 500.000 1.000 ;
  LAYER ME3 ;
  RECT 499.200 0.000 500.000 1.000 ;
  LAYER ME2 ;
  RECT 499.200 0.000 500.000 1.000 ;
  LAYER ME1 ;
  RECT 499.200 0.000 500.000 1.000 ;
 END
 ANTENNAPARTIALMETALAREA                  3.118 LAYER ME2 ;
 ANTENNAGATEAREA                          0.086 LAYER ME2 ;
 ANTENNAGATEAREA                          0.086 LAYER ME3 ;
 ANTENNAGATEAREA                          0.086 LAYER ME4 ;
 ANTENNADIFFAREA                          0.160 LAYER ME2 ;
 ANTENNADIFFAREA                          0.160 LAYER ME3 ;
 ANTENNADIFFAREA                          0.160 LAYER ME4 ;
 ANTENNAMAXAREACAR                       48.431 LAYER ME2 ;
 ANTENNAMAXAREACAR                       57.690 LAYER ME3 ;
 ANTENNAMAXAREACAR                       66.949 LAYER ME4 ;
END DI24
PIN DO23
  DIRECTION OUTPUT ;
 PORT
  LAYER ME4 ;
  RECT 492.800 0.000 493.600 1.000 ;
  LAYER ME3 ;
  RECT 492.800 0.000 493.600 1.000 ;
  LAYER ME2 ;
  RECT 492.800 0.000 493.600 1.000 ;
  LAYER ME1 ;
  RECT 492.800 0.000 493.600 1.000 ;
 END
 ANTENNAPARTIALMETALAREA                  4.148 LAYER ME2 ;
 ANTENNADIFFAREA                          5.472 LAYER ME2 ;
 ANTENNADIFFAREA                          5.472 LAYER ME3 ;
 ANTENNADIFFAREA                          5.472 LAYER ME4 ;
END DO23
PIN DI23
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 478.000 0.000 478.800 1.000 ;
  LAYER ME3 ;
  RECT 478.000 0.000 478.800 1.000 ;
  LAYER ME2 ;
  RECT 478.000 0.000 478.800 1.000 ;
  LAYER ME1 ;
  RECT 478.000 0.000 478.800 1.000 ;
 END
 ANTENNAPARTIALMETALAREA                  3.142 LAYER ME2 ;
 ANTENNAGATEAREA                          0.086 LAYER ME2 ;
 ANTENNAGATEAREA                          0.086 LAYER ME3 ;
 ANTENNAGATEAREA                          0.086 LAYER ME4 ;
 ANTENNADIFFAREA                          0.160 LAYER ME2 ;
 ANTENNADIFFAREA                          0.160 LAYER ME3 ;
 ANTENNADIFFAREA                          0.160 LAYER ME4 ;
 ANTENNAMAXAREACAR                       48.708 LAYER ME2 ;
 ANTENNAMAXAREACAR                       57.968 LAYER ME3 ;
 ANTENNAMAXAREACAR                       67.227 LAYER ME4 ;
END DI23
PIN DO22
  DIRECTION OUTPUT ;
 PORT
  LAYER ME4 ;
  RECT 472.800 0.000 473.600 1.000 ;
  LAYER ME3 ;
  RECT 472.800 0.000 473.600 1.000 ;
  LAYER ME2 ;
  RECT 472.800 0.000 473.600 1.000 ;
  LAYER ME1 ;
  RECT 472.800 0.000 473.600 1.000 ;
 END
 ANTENNAPARTIALMETALAREA                  4.164 LAYER ME2 ;
 ANTENNADIFFAREA                          5.472 LAYER ME2 ;
 ANTENNADIFFAREA                          5.472 LAYER ME3 ;
 ANTENNADIFFAREA                          5.472 LAYER ME4 ;
END DO22
PIN DI22
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 458.400 0.000 459.200 1.000 ;
  LAYER ME3 ;
  RECT 458.400 0.000 459.200 1.000 ;
  LAYER ME2 ;
  RECT 458.400 0.000 459.200 1.000 ;
  LAYER ME1 ;
  RECT 458.400 0.000 459.200 1.000 ;
 END
 ANTENNAPARTIALMETALAREA                  3.138 LAYER ME2 ;
 ANTENNAGATEAREA                          0.086 LAYER ME2 ;
 ANTENNAGATEAREA                          0.086 LAYER ME3 ;
 ANTENNAGATEAREA                          0.086 LAYER ME4 ;
 ANTENNADIFFAREA                          0.160 LAYER ME2 ;
 ANTENNADIFFAREA                          0.160 LAYER ME3 ;
 ANTENNADIFFAREA                          0.160 LAYER ME4 ;
 ANTENNAMAXAREACAR                       48.662 LAYER ME2 ;
 ANTENNAMAXAREACAR                       57.921 LAYER ME3 ;
 ANTENNAMAXAREACAR                       67.181 LAYER ME4 ;
END DI22
PIN DO21
  DIRECTION OUTPUT ;
 PORT
  LAYER ME4 ;
  RECT 452.000 0.000 452.800 1.000 ;
  LAYER ME3 ;
  RECT 452.000 0.000 452.800 1.000 ;
  LAYER ME2 ;
  RECT 452.000 0.000 452.800 1.000 ;
  LAYER ME1 ;
  RECT 452.000 0.000 452.800 1.000 ;
 END
 ANTENNAPARTIALMETALAREA                  4.172 LAYER ME2 ;
 ANTENNADIFFAREA                          5.472 LAYER ME2 ;
 ANTENNADIFFAREA                          5.472 LAYER ME3 ;
 ANTENNADIFFAREA                          5.472 LAYER ME4 ;
END DO21
PIN DI21
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 437.200 0.000 438.000 1.000 ;
  LAYER ME3 ;
  RECT 437.200 0.000 438.000 1.000 ;
  LAYER ME2 ;
  RECT 437.200 0.000 438.000 1.000 ;
  LAYER ME1 ;
  RECT 437.200 0.000 438.000 1.000 ;
 END
 ANTENNAPARTIALMETALAREA                  3.118 LAYER ME2 ;
 ANTENNAGATEAREA                          0.086 LAYER ME2 ;
 ANTENNAGATEAREA                          0.086 LAYER ME3 ;
 ANTENNAGATEAREA                          0.086 LAYER ME4 ;
 ANTENNADIFFAREA                          0.160 LAYER ME2 ;
 ANTENNADIFFAREA                          0.160 LAYER ME3 ;
 ANTENNADIFFAREA                          0.160 LAYER ME4 ;
 ANTENNAMAXAREACAR                       48.431 LAYER ME2 ;
 ANTENNAMAXAREACAR                       57.690 LAYER ME3 ;
 ANTENNAMAXAREACAR                       66.949 LAYER ME4 ;
END DI21
PIN DO20
  DIRECTION OUTPUT ;
 PORT
  LAYER ME4 ;
  RECT 432.000 0.000 432.800 1.000 ;
  LAYER ME3 ;
  RECT 432.000 0.000 432.800 1.000 ;
  LAYER ME2 ;
  RECT 432.000 0.000 432.800 1.000 ;
  LAYER ME1 ;
  RECT 432.000 0.000 432.800 1.000 ;
 END
 ANTENNAPARTIALMETALAREA                  4.140 LAYER ME2 ;
 ANTENNADIFFAREA                          5.472 LAYER ME2 ;
 ANTENNADIFFAREA                          5.472 LAYER ME3 ;
 ANTENNADIFFAREA                          5.472 LAYER ME4 ;
END DO20
PIN DI20
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 417.200 0.000 418.000 1.000 ;
  LAYER ME3 ;
  RECT 417.200 0.000 418.000 1.000 ;
  LAYER ME2 ;
  RECT 417.200 0.000 418.000 1.000 ;
  LAYER ME1 ;
  RECT 417.200 0.000 418.000 1.000 ;
 END
 ANTENNAPARTIALMETALAREA                  3.150 LAYER ME2 ;
 ANTENNAGATEAREA                          0.086 LAYER ME2 ;
 ANTENNAGATEAREA                          0.086 LAYER ME3 ;
 ANTENNAGATEAREA                          0.086 LAYER ME4 ;
 ANTENNADIFFAREA                          0.160 LAYER ME2 ;
 ANTENNADIFFAREA                          0.160 LAYER ME3 ;
 ANTENNADIFFAREA                          0.160 LAYER ME4 ;
 ANTENNAMAXAREACAR                       48.801 LAYER ME2 ;
 ANTENNAMAXAREACAR                       58.060 LAYER ME3 ;
 ANTENNAMAXAREACAR                       67.319 LAYER ME4 ;
END DI20
PIN DO19
  DIRECTION OUTPUT ;
 PORT
  LAYER ME4 ;
  RECT 410.800 0.000 411.600 1.000 ;
  LAYER ME3 ;
  RECT 410.800 0.000 411.600 1.000 ;
  LAYER ME2 ;
  RECT 410.800 0.000 411.600 1.000 ;
  LAYER ME1 ;
  RECT 410.800 0.000 411.600 1.000 ;
 END
 ANTENNAPARTIALMETALAREA                  4.164 LAYER ME2 ;
 ANTENNADIFFAREA                          5.472 LAYER ME2 ;
 ANTENNADIFFAREA                          5.472 LAYER ME3 ;
 ANTENNADIFFAREA                          5.472 LAYER ME4 ;
END DO19
PIN DI19
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 396.400 0.000 397.200 1.000 ;
  LAYER ME3 ;
  RECT 396.400 0.000 397.200 1.000 ;
  LAYER ME2 ;
  RECT 396.400 0.000 397.200 1.000 ;
  LAYER ME1 ;
  RECT 396.400 0.000 397.200 1.000 ;
 END
 ANTENNAPARTIALMETALAREA                  3.138 LAYER ME2 ;
 ANTENNAGATEAREA                          0.086 LAYER ME2 ;
 ANTENNAGATEAREA                          0.086 LAYER ME3 ;
 ANTENNAGATEAREA                          0.086 LAYER ME4 ;
 ANTENNADIFFAREA                          0.160 LAYER ME2 ;
 ANTENNADIFFAREA                          0.160 LAYER ME3 ;
 ANTENNADIFFAREA                          0.160 LAYER ME4 ;
 ANTENNAMAXAREACAR                       48.662 LAYER ME2 ;
 ANTENNAMAXAREACAR                       57.921 LAYER ME3 ;
 ANTENNAMAXAREACAR                       67.181 LAYER ME4 ;
END DI19
PIN DO18
  DIRECTION OUTPUT ;
 PORT
  LAYER ME4 ;
  RECT 391.200 0.000 392.000 1.000 ;
  LAYER ME3 ;
  RECT 391.200 0.000 392.000 1.000 ;
  LAYER ME2 ;
  RECT 391.200 0.000 392.000 1.000 ;
  LAYER ME1 ;
  RECT 391.200 0.000 392.000 1.000 ;
 END
 ANTENNAPARTIALMETALAREA                  4.164 LAYER ME2 ;
 ANTENNADIFFAREA                          5.472 LAYER ME2 ;
 ANTENNADIFFAREA                          5.472 LAYER ME3 ;
 ANTENNADIFFAREA                          5.472 LAYER ME4 ;
END DO18
PIN DI18
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 376.400 0.000 377.200 1.000 ;
  LAYER ME3 ;
  RECT 376.400 0.000 377.200 1.000 ;
  LAYER ME2 ;
  RECT 376.400 0.000 377.200 1.000 ;
  LAYER ME1 ;
  RECT 376.400 0.000 377.200 1.000 ;
 END
 ANTENNAPARTIALMETALAREA                  3.126 LAYER ME2 ;
 ANTENNAGATEAREA                          0.086 LAYER ME2 ;
 ANTENNAGATEAREA                          0.086 LAYER ME3 ;
 ANTENNAGATEAREA                          0.086 LAYER ME4 ;
 ANTENNADIFFAREA                          0.160 LAYER ME2 ;
 ANTENNADIFFAREA                          0.160 LAYER ME3 ;
 ANTENNADIFFAREA                          0.160 LAYER ME4 ;
 ANTENNAMAXAREACAR                       48.523 LAYER ME2 ;
 ANTENNAMAXAREACAR                       57.782 LAYER ME3 ;
 ANTENNAMAXAREACAR                       67.042 LAYER ME4 ;
END DI18
PIN DO17
  DIRECTION OUTPUT ;
 PORT
  LAYER ME4 ;
  RECT 370.000 0.000 370.800 1.000 ;
  LAYER ME3 ;
  RECT 370.000 0.000 370.800 1.000 ;
  LAYER ME2 ;
  RECT 370.000 0.000 370.800 1.000 ;
  LAYER ME1 ;
  RECT 370.000 0.000 370.800 1.000 ;
 END
 ANTENNAPARTIALMETALAREA                  4.140 LAYER ME2 ;
 ANTENNADIFFAREA                          5.472 LAYER ME2 ;
 ANTENNADIFFAREA                          5.472 LAYER ME3 ;
 ANTENNADIFFAREA                          5.472 LAYER ME4 ;
END DO17
PIN DI17
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 355.200 0.000 356.000 1.000 ;
  LAYER ME3 ;
  RECT 355.200 0.000 356.000 1.000 ;
  LAYER ME2 ;
  RECT 355.200 0.000 356.000 1.000 ;
  LAYER ME1 ;
  RECT 355.200 0.000 356.000 1.000 ;
 END
 ANTENNAPARTIALMETALAREA                  3.150 LAYER ME2 ;
 ANTENNAGATEAREA                          0.086 LAYER ME2 ;
 ANTENNAGATEAREA                          0.086 LAYER ME3 ;
 ANTENNAGATEAREA                          0.086 LAYER ME4 ;
 ANTENNADIFFAREA                          0.160 LAYER ME2 ;
 ANTENNADIFFAREA                          0.160 LAYER ME3 ;
 ANTENNADIFFAREA                          0.160 LAYER ME4 ;
 ANTENNAMAXAREACAR                       48.801 LAYER ME2 ;
 ANTENNAMAXAREACAR                       58.060 LAYER ME3 ;
 ANTENNAMAXAREACAR                       67.319 LAYER ME4 ;
END DI17
PIN DO16
  DIRECTION OUTPUT ;
 PORT
  LAYER ME4 ;
  RECT 350.000 0.000 350.800 1.000 ;
  LAYER ME3 ;
  RECT 350.000 0.000 350.800 1.000 ;
  LAYER ME2 ;
  RECT 350.000 0.000 350.800 1.000 ;
  LAYER ME1 ;
  RECT 350.000 0.000 350.800 1.000 ;
 END
 ANTENNAPARTIALMETALAREA                  4.172 LAYER ME2 ;
 ANTENNADIFFAREA                          5.472 LAYER ME2 ;
 ANTENNADIFFAREA                          5.472 LAYER ME3 ;
 ANTENNADIFFAREA                          5.472 LAYER ME4 ;
END DO16
PIN WEB2
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 337.200 0.000 338.000 1.000 ;
  LAYER ME3 ;
  RECT 337.200 0.000 338.000 1.000 ;
  LAYER ME2 ;
  RECT 337.200 0.000 338.000 1.000 ;
  LAYER ME1 ;
  RECT 337.200 0.000 338.000 1.000 ;
 END
 ANTENNAPARTIALMETALAREA                  2.840 LAYER ME2 ;
 ANTENNAGATEAREA                          0.072 LAYER ME2 ;
 ANTENNAGATEAREA                          0.072 LAYER ME3 ;
 ANTENNAGATEAREA                          0.072 LAYER ME4 ;
 ANTENNADIFFAREA                          0.160 LAYER ME2 ;
 ANTENNADIFFAREA                          0.160 LAYER ME3 ;
 ANTENNADIFFAREA                          0.160 LAYER ME4 ;
 ANTENNAMAXAREACAR                       54.456 LAYER ME2 ;
 ANTENNAMAXAREACAR                       65.567 LAYER ME3 ;
 ANTENNAMAXAREACAR                       76.678 LAYER ME4 ;
END WEB2
PIN DI16
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 335.600 0.000 336.400 1.000 ;
  LAYER ME3 ;
  RECT 335.600 0.000 336.400 1.000 ;
  LAYER ME2 ;
  RECT 335.600 0.000 336.400 1.000 ;
  LAYER ME1 ;
  RECT 335.600 0.000 336.400 1.000 ;
 END
 ANTENNAPARTIALMETALAREA                  3.130 LAYER ME2 ;
 ANTENNAGATEAREA                          0.086 LAYER ME2 ;
 ANTENNAGATEAREA                          0.086 LAYER ME3 ;
 ANTENNAGATEAREA                          0.086 LAYER ME4 ;
 ANTENNADIFFAREA                          0.160 LAYER ME2 ;
 ANTENNADIFFAREA                          0.160 LAYER ME3 ;
 ANTENNADIFFAREA                          0.160 LAYER ME4 ;
 ANTENNAMAXAREACAR                       48.569 LAYER ME2 ;
 ANTENNAMAXAREACAR                       57.829 LAYER ME3 ;
 ANTENNAMAXAREACAR                       67.088 LAYER ME4 ;
END DI16
PIN DO15
  DIRECTION OUTPUT ;
 PORT
  LAYER ME4 ;
  RECT 329.200 0.000 330.000 1.000 ;
  LAYER ME3 ;
  RECT 329.200 0.000 330.000 1.000 ;
  LAYER ME2 ;
  RECT 329.200 0.000 330.000 1.000 ;
  LAYER ME1 ;
  RECT 329.200 0.000 330.000 1.000 ;
 END
 ANTENNAPARTIALMETALAREA                  4.164 LAYER ME2 ;
 ANTENNADIFFAREA                          5.472 LAYER ME2 ;
 ANTENNADIFFAREA                          5.472 LAYER ME3 ;
 ANTENNADIFFAREA                          5.472 LAYER ME4 ;
END DO15
PIN DI15
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 314.400 0.000 315.200 1.000 ;
  LAYER ME3 ;
  RECT 314.400 0.000 315.200 1.000 ;
  LAYER ME2 ;
  RECT 314.400 0.000 315.200 1.000 ;
  LAYER ME1 ;
  RECT 314.400 0.000 315.200 1.000 ;
 END
 ANTENNAPARTIALMETALAREA                  3.126 LAYER ME2 ;
 ANTENNAGATEAREA                          0.086 LAYER ME2 ;
 ANTENNAGATEAREA                          0.086 LAYER ME3 ;
 ANTENNAGATEAREA                          0.086 LAYER ME4 ;
 ANTENNADIFFAREA                          0.160 LAYER ME2 ;
 ANTENNADIFFAREA                          0.160 LAYER ME3 ;
 ANTENNADIFFAREA                          0.160 LAYER ME4 ;
 ANTENNAMAXAREACAR                       48.523 LAYER ME2 ;
 ANTENNAMAXAREACAR                       57.782 LAYER ME3 ;
 ANTENNAMAXAREACAR                       67.042 LAYER ME4 ;
END DI15
PIN DO14
  DIRECTION OUTPUT ;
 PORT
  LAYER ME4 ;
  RECT 309.200 0.000 310.000 1.000 ;
  LAYER ME3 ;
  RECT 309.200 0.000 310.000 1.000 ;
  LAYER ME2 ;
  RECT 309.200 0.000 310.000 1.000 ;
  LAYER ME1 ;
  RECT 309.200 0.000 310.000 1.000 ;
 END
 ANTENNAPARTIALMETALAREA                  4.148 LAYER ME2 ;
 ANTENNADIFFAREA                          5.472 LAYER ME2 ;
 ANTENNADIFFAREA                          5.472 LAYER ME3 ;
 ANTENNADIFFAREA                          5.472 LAYER ME4 ;
END DO14
PIN DI14
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 294.800 0.000 295.600 1.000 ;
  LAYER ME3 ;
  RECT 294.800 0.000 295.600 1.000 ;
  LAYER ME2 ;
  RECT 294.800 0.000 295.600 1.000 ;
  LAYER ME1 ;
  RECT 294.800 0.000 295.600 1.000 ;
 END
 ANTENNAPARTIALMETALAREA                  3.154 LAYER ME2 ;
 ANTENNAGATEAREA                          0.086 LAYER ME2 ;
 ANTENNAGATEAREA                          0.086 LAYER ME3 ;
 ANTENNAGATEAREA                          0.086 LAYER ME4 ;
 ANTENNADIFFAREA                          0.160 LAYER ME2 ;
 ANTENNADIFFAREA                          0.160 LAYER ME3 ;
 ANTENNADIFFAREA                          0.160 LAYER ME4 ;
 ANTENNAMAXAREACAR                       48.847 LAYER ME2 ;
 ANTENNAMAXAREACAR                       58.106 LAYER ME3 ;
 ANTENNAMAXAREACAR                       67.366 LAYER ME4 ;
END DI14
PIN DO13
  DIRECTION OUTPUT ;
 PORT
  LAYER ME4 ;
  RECT 288.000 0.000 288.800 1.000 ;
  LAYER ME3 ;
  RECT 288.000 0.000 288.800 1.000 ;
  LAYER ME2 ;
  RECT 288.000 0.000 288.800 1.000 ;
  LAYER ME1 ;
  RECT 288.000 0.000 288.800 1.000 ;
 END
 ANTENNAPARTIALMETALAREA                  4.172 LAYER ME2 ;
 ANTENNADIFFAREA                          5.472 LAYER ME2 ;
 ANTENNADIFFAREA                          5.472 LAYER ME3 ;
 ANTENNADIFFAREA                          5.472 LAYER ME4 ;
END DO13
PIN DI13
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 273.600 0.000 274.400 1.000 ;
  LAYER ME3 ;
  RECT 273.600 0.000 274.400 1.000 ;
  LAYER ME2 ;
  RECT 273.600 0.000 274.400 1.000 ;
  LAYER ME1 ;
  RECT 273.600 0.000 274.400 1.000 ;
 END
 ANTENNAPARTIALMETALAREA                  3.130 LAYER ME2 ;
 ANTENNAGATEAREA                          0.086 LAYER ME2 ;
 ANTENNAGATEAREA                          0.086 LAYER ME3 ;
 ANTENNAGATEAREA                          0.086 LAYER ME4 ;
 ANTENNADIFFAREA                          0.160 LAYER ME2 ;
 ANTENNADIFFAREA                          0.160 LAYER ME3 ;
 ANTENNADIFFAREA                          0.160 LAYER ME4 ;
 ANTENNAMAXAREACAR                       48.569 LAYER ME2 ;
 ANTENNAMAXAREACAR                       57.829 LAYER ME3 ;
 ANTENNAMAXAREACAR                       67.088 LAYER ME4 ;
END DI13
PIN DO12
  DIRECTION OUTPUT ;
 PORT
  LAYER ME4 ;
  RECT 268.400 0.000 269.200 1.000 ;
  LAYER ME3 ;
  RECT 268.400 0.000 269.200 1.000 ;
  LAYER ME2 ;
  RECT 268.400 0.000 269.200 1.000 ;
  LAYER ME1 ;
  RECT 268.400 0.000 269.200 1.000 ;
 END
 ANTENNAPARTIALMETALAREA                  4.156 LAYER ME2 ;
 ANTENNADIFFAREA                          5.472 LAYER ME2 ;
 ANTENNADIFFAREA                          5.472 LAYER ME3 ;
 ANTENNADIFFAREA                          5.472 LAYER ME4 ;
END DO12
PIN DI12
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 253.600 0.000 254.400 1.000 ;
  LAYER ME3 ;
  RECT 253.600 0.000 254.400 1.000 ;
  LAYER ME2 ;
  RECT 253.600 0.000 254.400 1.000 ;
  LAYER ME1 ;
  RECT 253.600 0.000 254.400 1.000 ;
 END
 ANTENNAPARTIALMETALAREA                  3.134 LAYER ME2 ;
 ANTENNAGATEAREA                          0.086 LAYER ME2 ;
 ANTENNAGATEAREA                          0.086 LAYER ME3 ;
 ANTENNAGATEAREA                          0.086 LAYER ME4 ;
 ANTENNADIFFAREA                          0.160 LAYER ME2 ;
 ANTENNADIFFAREA                          0.160 LAYER ME3 ;
 ANTENNADIFFAREA                          0.160 LAYER ME4 ;
 ANTENNAMAXAREACAR                       48.616 LAYER ME2 ;
 ANTENNAMAXAREACAR                       57.875 LAYER ME3 ;
 ANTENNAMAXAREACAR                       67.134 LAYER ME4 ;
END DI12
PIN DO11
  DIRECTION OUTPUT ;
 PORT
  LAYER ME4 ;
  RECT 247.200 0.000 248.000 1.000 ;
  LAYER ME3 ;
  RECT 247.200 0.000 248.000 1.000 ;
  LAYER ME2 ;
  RECT 247.200 0.000 248.000 1.000 ;
  LAYER ME1 ;
  RECT 247.200 0.000 248.000 1.000 ;
 END
 ANTENNAPARTIALMETALAREA                  4.148 LAYER ME2 ;
 ANTENNADIFFAREA                          5.472 LAYER ME2 ;
 ANTENNADIFFAREA                          5.472 LAYER ME3 ;
 ANTENNADIFFAREA                          5.472 LAYER ME4 ;
END DO11
PIN DI11
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 232.800 0.000 233.600 1.000 ;
  LAYER ME3 ;
  RECT 232.800 0.000 233.600 1.000 ;
  LAYER ME2 ;
  RECT 232.800 0.000 233.600 1.000 ;
  LAYER ME1 ;
  RECT 232.800 0.000 233.600 1.000 ;
 END
 ANTENNAPARTIALMETALAREA                  3.154 LAYER ME2 ;
 ANTENNAGATEAREA                          0.086 LAYER ME2 ;
 ANTENNAGATEAREA                          0.086 LAYER ME3 ;
 ANTENNAGATEAREA                          0.086 LAYER ME4 ;
 ANTENNADIFFAREA                          0.160 LAYER ME2 ;
 ANTENNADIFFAREA                          0.160 LAYER ME3 ;
 ANTENNADIFFAREA                          0.160 LAYER ME4 ;
 ANTENNAMAXAREACAR                       48.847 LAYER ME2 ;
 ANTENNAMAXAREACAR                       58.106 LAYER ME3 ;
 ANTENNAMAXAREACAR                       67.366 LAYER ME4 ;
END DI11
PIN DO10
  DIRECTION OUTPUT ;
 PORT
  LAYER ME4 ;
  RECT 227.200 0.000 228.000 1.000 ;
  LAYER ME3 ;
  RECT 227.200 0.000 228.000 1.000 ;
  LAYER ME2 ;
  RECT 227.200 0.000 228.000 1.000 ;
  LAYER ME1 ;
  RECT 227.200 0.000 228.000 1.000 ;
 END
 ANTENNAPARTIALMETALAREA                  4.180 LAYER ME2 ;
 ANTENNADIFFAREA                          5.472 LAYER ME2 ;
 ANTENNADIFFAREA                          5.472 LAYER ME3 ;
 ANTENNADIFFAREA                          5.472 LAYER ME4 ;
END DO10
PIN DI10
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 212.800 0.000 213.600 1.000 ;
  LAYER ME3 ;
  RECT 212.800 0.000 213.600 1.000 ;
  LAYER ME2 ;
  RECT 212.800 0.000 213.600 1.000 ;
  LAYER ME1 ;
  RECT 212.800 0.000 213.600 1.000 ;
 END
 ANTENNAPARTIALMETALAREA                  3.122 LAYER ME2 ;
 ANTENNAGATEAREA                          0.086 LAYER ME2 ;
 ANTENNAGATEAREA                          0.086 LAYER ME3 ;
 ANTENNAGATEAREA                          0.086 LAYER ME4 ;
 ANTENNADIFFAREA                          0.160 LAYER ME2 ;
 ANTENNADIFFAREA                          0.160 LAYER ME3 ;
 ANTENNADIFFAREA                          0.160 LAYER ME4 ;
 ANTENNAMAXAREACAR                       48.477 LAYER ME2 ;
 ANTENNAMAXAREACAR                       57.736 LAYER ME3 ;
 ANTENNAMAXAREACAR                       66.995 LAYER ME4 ;
END DI10
PIN DO9
  DIRECTION OUTPUT ;
 PORT
  LAYER ME4 ;
  RECT 206.400 0.000 207.200 1.000 ;
  LAYER ME3 ;
  RECT 206.400 0.000 207.200 1.000 ;
  LAYER ME2 ;
  RECT 206.400 0.000 207.200 1.000 ;
  LAYER ME1 ;
  RECT 206.400 0.000 207.200 1.000 ;
 END
 ANTENNAPARTIALMETALAREA                  4.156 LAYER ME2 ;
 ANTENNADIFFAREA                          5.472 LAYER ME2 ;
 ANTENNADIFFAREA                          5.472 LAYER ME3 ;
 ANTENNADIFFAREA                          5.472 LAYER ME4 ;
END DO9
PIN DI9
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 191.600 0.000 192.400 1.000 ;
  LAYER ME3 ;
  RECT 191.600 0.000 192.400 1.000 ;
  LAYER ME2 ;
  RECT 191.600 0.000 192.400 1.000 ;
  LAYER ME1 ;
  RECT 191.600 0.000 192.400 1.000 ;
 END
 ANTENNAPARTIALMETALAREA                  3.134 LAYER ME2 ;
 ANTENNAGATEAREA                          0.086 LAYER ME2 ;
 ANTENNAGATEAREA                          0.086 LAYER ME3 ;
 ANTENNAGATEAREA                          0.086 LAYER ME4 ;
 ANTENNADIFFAREA                          0.160 LAYER ME2 ;
 ANTENNADIFFAREA                          0.160 LAYER ME3 ;
 ANTENNADIFFAREA                          0.160 LAYER ME4 ;
 ANTENNAMAXAREACAR                       48.616 LAYER ME2 ;
 ANTENNAMAXAREACAR                       57.875 LAYER ME3 ;
 ANTENNAMAXAREACAR                       67.134 LAYER ME4 ;
END DI9
PIN DO8
  DIRECTION OUTPUT ;
 PORT
  LAYER ME4 ;
  RECT 186.400 0.000 187.200 1.000 ;
  LAYER ME3 ;
  RECT 186.400 0.000 187.200 1.000 ;
  LAYER ME2 ;
  RECT 186.400 0.000 187.200 1.000 ;
  LAYER ME1 ;
  RECT 186.400 0.000 187.200 1.000 ;
 END
 ANTENNAPARTIALMETALAREA                  4.156 LAYER ME2 ;
 ANTENNADIFFAREA                          5.472 LAYER ME2 ;
 ANTENNADIFFAREA                          5.472 LAYER ME3 ;
 ANTENNADIFFAREA                          5.472 LAYER ME4 ;
END DO8
PIN WEB1
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 173.600 0.000 174.400 1.000 ;
  LAYER ME3 ;
  RECT 173.600 0.000 174.400 1.000 ;
  LAYER ME2 ;
  RECT 173.600 0.000 174.400 1.000 ;
  LAYER ME1 ;
  RECT 173.600 0.000 174.400 1.000 ;
 END
 ANTENNAPARTIALMETALAREA                  2.836 LAYER ME2 ;
 ANTENNAGATEAREA                          0.072 LAYER ME2 ;
 ANTENNAGATEAREA                          0.072 LAYER ME3 ;
 ANTENNAGATEAREA                          0.072 LAYER ME4 ;
 ANTENNADIFFAREA                          0.160 LAYER ME2 ;
 ANTENNADIFFAREA                          0.160 LAYER ME3 ;
 ANTENNADIFFAREA                          0.160 LAYER ME4 ;
 ANTENNAMAXAREACAR                       54.400 LAYER ME2 ;
 ANTENNAMAXAREACAR                       65.511 LAYER ME3 ;
 ANTENNAMAXAREACAR                       76.622 LAYER ME4 ;
END WEB1
PIN DI8
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 172.000 0.000 172.800 1.000 ;
  LAYER ME3 ;
  RECT 172.000 0.000 172.800 1.000 ;
  LAYER ME2 ;
  RECT 172.000 0.000 172.800 1.000 ;
  LAYER ME1 ;
  RECT 172.000 0.000 172.800 1.000 ;
 END
 ANTENNAPARTIALMETALAREA                  3.146 LAYER ME2 ;
 ANTENNAGATEAREA                          0.086 LAYER ME2 ;
 ANTENNAGATEAREA                          0.086 LAYER ME3 ;
 ANTENNAGATEAREA                          0.086 LAYER ME4 ;
 ANTENNADIFFAREA                          0.160 LAYER ME2 ;
 ANTENNADIFFAREA                          0.160 LAYER ME3 ;
 ANTENNADIFFAREA                          0.160 LAYER ME4 ;
 ANTENNAMAXAREACAR                       48.755 LAYER ME2 ;
 ANTENNAMAXAREACAR                       58.014 LAYER ME3 ;
 ANTENNAMAXAREACAR                       67.273 LAYER ME4 ;
END DI8
PIN DO7
  DIRECTION OUTPUT ;
 PORT
  LAYER ME4 ;
  RECT 165.200 0.000 166.000 1.000 ;
  LAYER ME3 ;
  RECT 165.200 0.000 166.000 1.000 ;
  LAYER ME2 ;
  RECT 165.200 0.000 166.000 1.000 ;
  LAYER ME1 ;
  RECT 165.200 0.000 166.000 1.000 ;
 END
 ANTENNAPARTIALMETALAREA                  4.180 LAYER ME2 ;
 ANTENNADIFFAREA                          5.472 LAYER ME2 ;
 ANTENNADIFFAREA                          5.472 LAYER ME3 ;
 ANTENNADIFFAREA                          5.472 LAYER ME4 ;
END DO7
PIN DI7
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 150.800 0.000 151.600 1.000 ;
  LAYER ME3 ;
  RECT 150.800 0.000 151.600 1.000 ;
  LAYER ME2 ;
  RECT 150.800 0.000 151.600 1.000 ;
  LAYER ME1 ;
  RECT 150.800 0.000 151.600 1.000 ;
 END
 ANTENNAPARTIALMETALAREA                  3.122 LAYER ME2 ;
 ANTENNAGATEAREA                          0.086 LAYER ME2 ;
 ANTENNAGATEAREA                          0.086 LAYER ME3 ;
 ANTENNAGATEAREA                          0.086 LAYER ME4 ;
 ANTENNADIFFAREA                          0.160 LAYER ME2 ;
 ANTENNADIFFAREA                          0.160 LAYER ME3 ;
 ANTENNADIFFAREA                          0.160 LAYER ME4 ;
 ANTENNAMAXAREACAR                       48.477 LAYER ME2 ;
 ANTENNAMAXAREACAR                       57.736 LAYER ME3 ;
 ANTENNAMAXAREACAR                       66.995 LAYER ME4 ;
END DI7
PIN DO6
  DIRECTION OUTPUT ;
 PORT
  LAYER ME4 ;
  RECT 145.600 0.000 146.400 1.000 ;
  LAYER ME3 ;
  RECT 145.600 0.000 146.400 1.000 ;
  LAYER ME2 ;
  RECT 145.600 0.000 146.400 1.000 ;
  LAYER ME1 ;
  RECT 145.600 0.000 146.400 1.000 ;
 END
 ANTENNAPARTIALMETALAREA                  4.148 LAYER ME2 ;
 ANTENNADIFFAREA                          5.472 LAYER ME2 ;
 ANTENNADIFFAREA                          5.472 LAYER ME3 ;
 ANTENNADIFFAREA                          5.472 LAYER ME4 ;
END DO6
PIN DI6
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 130.800 0.000 131.600 1.000 ;
  LAYER ME3 ;
  RECT 130.800 0.000 131.600 1.000 ;
  LAYER ME2 ;
  RECT 130.800 0.000 131.600 1.000 ;
  LAYER ME1 ;
  RECT 130.800 0.000 131.600 1.000 ;
 END
 ANTENNAPARTIALMETALAREA                  3.142 LAYER ME2 ;
 ANTENNAGATEAREA                          0.086 LAYER ME2 ;
 ANTENNAGATEAREA                          0.086 LAYER ME3 ;
 ANTENNAGATEAREA                          0.086 LAYER ME4 ;
 ANTENNADIFFAREA                          0.160 LAYER ME2 ;
 ANTENNADIFFAREA                          0.160 LAYER ME3 ;
 ANTENNADIFFAREA                          0.160 LAYER ME4 ;
 ANTENNAMAXAREACAR                       48.708 LAYER ME2 ;
 ANTENNAMAXAREACAR                       57.968 LAYER ME3 ;
 ANTENNAMAXAREACAR                       67.227 LAYER ME4 ;
END DI6
PIN DO5
  DIRECTION OUTPUT ;
 PORT
  LAYER ME4 ;
  RECT 124.400 0.000 125.200 1.000 ;
  LAYER ME3 ;
  RECT 124.400 0.000 125.200 1.000 ;
  LAYER ME2 ;
  RECT 124.400 0.000 125.200 1.000 ;
  LAYER ME1 ;
  RECT 124.400 0.000 125.200 1.000 ;
 END
 ANTENNAPARTIALMETALAREA                  4.156 LAYER ME2 ;
 ANTENNADIFFAREA                          5.472 LAYER ME2 ;
 ANTENNADIFFAREA                          5.472 LAYER ME3 ;
 ANTENNADIFFAREA                          5.472 LAYER ME4 ;
END DO5
PIN DI5
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 110.000 0.000 110.800 1.000 ;
  LAYER ME3 ;
  RECT 110.000 0.000 110.800 1.000 ;
  LAYER ME2 ;
  RECT 110.000 0.000 110.800 1.000 ;
  LAYER ME1 ;
  RECT 110.000 0.000 110.800 1.000 ;
 END
 ANTENNAPARTIALMETALAREA                  3.146 LAYER ME2 ;
 ANTENNAGATEAREA                          0.086 LAYER ME2 ;
 ANTENNAGATEAREA                          0.086 LAYER ME3 ;
 ANTENNAGATEAREA                          0.086 LAYER ME4 ;
 ANTENNADIFFAREA                          0.160 LAYER ME2 ;
 ANTENNADIFFAREA                          0.160 LAYER ME3 ;
 ANTENNADIFFAREA                          0.160 LAYER ME4 ;
 ANTENNAMAXAREACAR                       48.755 LAYER ME2 ;
 ANTENNAMAXAREACAR                       58.014 LAYER ME3 ;
 ANTENNAMAXAREACAR                       67.273 LAYER ME4 ;
END DI5
PIN DO4
  DIRECTION OUTPUT ;
 PORT
  LAYER ME4 ;
  RECT 104.800 0.000 105.600 1.000 ;
  LAYER ME3 ;
  RECT 104.800 0.000 105.600 1.000 ;
  LAYER ME2 ;
  RECT 104.800 0.000 105.600 1.000 ;
  LAYER ME1 ;
  RECT 104.800 0.000 105.600 1.000 ;
 END
 ANTENNAPARTIALMETALAREA                  4.172 LAYER ME2 ;
 ANTENNADIFFAREA                          5.472 LAYER ME2 ;
 ANTENNADIFFAREA                          5.472 LAYER ME3 ;
 ANTENNADIFFAREA                          5.472 LAYER ME4 ;
END DO4
PIN DI4
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 90.000 0.000 90.800 1.000 ;
  LAYER ME3 ;
  RECT 90.000 0.000 90.800 1.000 ;
  LAYER ME2 ;
  RECT 90.000 0.000 90.800 1.000 ;
  LAYER ME1 ;
  RECT 90.000 0.000 90.800 1.000 ;
 END
 ANTENNAPARTIALMETALAREA                  3.118 LAYER ME2 ;
 ANTENNAGATEAREA                          0.086 LAYER ME2 ;
 ANTENNAGATEAREA                          0.086 LAYER ME3 ;
 ANTENNAGATEAREA                          0.086 LAYER ME4 ;
 ANTENNADIFFAREA                          0.160 LAYER ME2 ;
 ANTENNADIFFAREA                          0.160 LAYER ME3 ;
 ANTENNADIFFAREA                          0.160 LAYER ME4 ;
 ANTENNAMAXAREACAR                       48.431 LAYER ME2 ;
 ANTENNAMAXAREACAR                       57.690 LAYER ME3 ;
 ANTENNAMAXAREACAR                       66.949 LAYER ME4 ;
END DI4
PIN DO3
  DIRECTION OUTPUT ;
 PORT
  LAYER ME4 ;
  RECT 83.600 0.000 84.400 1.000 ;
  LAYER ME3 ;
  RECT 83.600 0.000 84.400 1.000 ;
  LAYER ME2 ;
  RECT 83.600 0.000 84.400 1.000 ;
  LAYER ME1 ;
  RECT 83.600 0.000 84.400 1.000 ;
 END
 ANTENNAPARTIALMETALAREA                  4.148 LAYER ME2 ;
 ANTENNADIFFAREA                          5.472 LAYER ME2 ;
 ANTENNADIFFAREA                          5.472 LAYER ME3 ;
 ANTENNADIFFAREA                          5.472 LAYER ME4 ;
END DO3
PIN DI3
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 68.800 0.000 69.600 1.000 ;
  LAYER ME3 ;
  RECT 68.800 0.000 69.600 1.000 ;
  LAYER ME2 ;
  RECT 68.800 0.000 69.600 1.000 ;
  LAYER ME1 ;
  RECT 68.800 0.000 69.600 1.000 ;
 END
 ANTENNAPARTIALMETALAREA                  3.142 LAYER ME2 ;
 ANTENNAGATEAREA                          0.086 LAYER ME2 ;
 ANTENNAGATEAREA                          0.086 LAYER ME3 ;
 ANTENNAGATEAREA                          0.086 LAYER ME4 ;
 ANTENNADIFFAREA                          0.160 LAYER ME2 ;
 ANTENNADIFFAREA                          0.160 LAYER ME3 ;
 ANTENNADIFFAREA                          0.160 LAYER ME4 ;
 ANTENNAMAXAREACAR                       48.708 LAYER ME2 ;
 ANTENNAMAXAREACAR                       57.968 LAYER ME3 ;
 ANTENNAMAXAREACAR                       67.227 LAYER ME4 ;
END DI3
PIN DO2
  DIRECTION OUTPUT ;
 PORT
  LAYER ME4 ;
  RECT 63.600 0.000 64.400 1.000 ;
  LAYER ME3 ;
  RECT 63.600 0.000 64.400 1.000 ;
  LAYER ME2 ;
  RECT 63.600 0.000 64.400 1.000 ;
  LAYER ME1 ;
  RECT 63.600 0.000 64.400 1.000 ;
 END
 ANTENNAPARTIALMETALAREA                  4.164 LAYER ME2 ;
 ANTENNADIFFAREA                          5.472 LAYER ME2 ;
 ANTENNADIFFAREA                          5.472 LAYER ME3 ;
 ANTENNADIFFAREA                          5.472 LAYER ME4 ;
END DO2
PIN DI2
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 49.200 0.000 50.000 1.000 ;
  LAYER ME3 ;
  RECT 49.200 0.000 50.000 1.000 ;
  LAYER ME2 ;
  RECT 49.200 0.000 50.000 1.000 ;
  LAYER ME1 ;
  RECT 49.200 0.000 50.000 1.000 ;
 END
 ANTENNAPARTIALMETALAREA                  3.138 LAYER ME2 ;
 ANTENNAGATEAREA                          0.086 LAYER ME2 ;
 ANTENNAGATEAREA                          0.086 LAYER ME3 ;
 ANTENNAGATEAREA                          0.086 LAYER ME4 ;
 ANTENNADIFFAREA                          0.160 LAYER ME2 ;
 ANTENNADIFFAREA                          0.160 LAYER ME3 ;
 ANTENNADIFFAREA                          0.160 LAYER ME4 ;
 ANTENNAMAXAREACAR                       48.662 LAYER ME2 ;
 ANTENNAMAXAREACAR                       57.921 LAYER ME3 ;
 ANTENNAMAXAREACAR                       67.181 LAYER ME4 ;
END DI2
PIN DO1
  DIRECTION OUTPUT ;
 PORT
  LAYER ME4 ;
  RECT 42.800 0.000 43.600 1.000 ;
  LAYER ME3 ;
  RECT 42.800 0.000 43.600 1.000 ;
  LAYER ME2 ;
  RECT 42.800 0.000 43.600 1.000 ;
  LAYER ME1 ;
  RECT 42.800 0.000 43.600 1.000 ;
 END
 ANTENNAPARTIALMETALAREA                  4.172 LAYER ME2 ;
 ANTENNADIFFAREA                          5.472 LAYER ME2 ;
 ANTENNADIFFAREA                          5.472 LAYER ME3 ;
 ANTENNADIFFAREA                          5.472 LAYER ME4 ;
END DO1
PIN DI1
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 28.000 0.000 28.800 1.000 ;
  LAYER ME3 ;
  RECT 28.000 0.000 28.800 1.000 ;
  LAYER ME2 ;
  RECT 28.000 0.000 28.800 1.000 ;
  LAYER ME1 ;
  RECT 28.000 0.000 28.800 1.000 ;
 END
 ANTENNAPARTIALMETALAREA                  3.118 LAYER ME2 ;
 ANTENNAGATEAREA                          0.086 LAYER ME2 ;
 ANTENNAGATEAREA                          0.086 LAYER ME3 ;
 ANTENNAGATEAREA                          0.086 LAYER ME4 ;
 ANTENNADIFFAREA                          0.160 LAYER ME2 ;
 ANTENNADIFFAREA                          0.160 LAYER ME3 ;
 ANTENNADIFFAREA                          0.160 LAYER ME4 ;
 ANTENNAMAXAREACAR                       48.431 LAYER ME2 ;
 ANTENNAMAXAREACAR                       57.690 LAYER ME3 ;
 ANTENNAMAXAREACAR                       66.949 LAYER ME4 ;
END DI1
PIN DO0
  DIRECTION OUTPUT ;
 PORT
  LAYER ME4 ;
  RECT 22.800 0.000 23.600 1.000 ;
  LAYER ME3 ;
  RECT 22.800 0.000 23.600 1.000 ;
  LAYER ME2 ;
  RECT 22.800 0.000 23.600 1.000 ;
  LAYER ME1 ;
  RECT 22.800 0.000 23.600 1.000 ;
 END
 ANTENNAPARTIALMETALAREA                  4.140 LAYER ME2 ;
 ANTENNADIFFAREA                          5.472 LAYER ME2 ;
 ANTENNADIFFAREA                          5.472 LAYER ME3 ;
 ANTENNADIFFAREA                          5.472 LAYER ME4 ;
END DO0
PIN WEB0
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 10.000 0.000 10.800 1.000 ;
  LAYER ME3 ;
  RECT 10.000 0.000 10.800 1.000 ;
  LAYER ME2 ;
  RECT 10.000 0.000 10.800 1.000 ;
  LAYER ME1 ;
  RECT 10.000 0.000 10.800 1.000 ;
 END
 ANTENNAPARTIALMETALAREA                  2.852 LAYER ME2 ;
 ANTENNAGATEAREA                          0.072 LAYER ME2 ;
 ANTENNAGATEAREA                          0.072 LAYER ME3 ;
 ANTENNAGATEAREA                          0.072 LAYER ME4 ;
 ANTENNADIFFAREA                          0.160 LAYER ME2 ;
 ANTENNADIFFAREA                          0.160 LAYER ME3 ;
 ANTENNADIFFAREA                          0.160 LAYER ME4 ;
 ANTENNAMAXAREACAR                       54.622 LAYER ME2 ;
 ANTENNAMAXAREACAR                       65.733 LAYER ME3 ;
 ANTENNAMAXAREACAR                       76.844 LAYER ME4 ;
END WEB0
PIN DI0
  DIRECTION INPUT ;
 PORT
  LAYER ME4 ;
  RECT 8.000 0.000 8.800 1.000 ;
  LAYER ME3 ;
  RECT 8.000 0.000 8.800 1.000 ;
  LAYER ME2 ;
  RECT 8.000 0.000 8.800 1.000 ;
  LAYER ME1 ;
  RECT 8.000 0.000 8.800 1.000 ;
 END
 ANTENNAPARTIALMETALAREA                  3.150 LAYER ME2 ;
 ANTENNAGATEAREA                          0.086 LAYER ME2 ;
 ANTENNAGATEAREA                          0.086 LAYER ME3 ;
 ANTENNAGATEAREA                          0.086 LAYER ME4 ;
 ANTENNADIFFAREA                          0.160 LAYER ME2 ;
 ANTENNADIFFAREA                          0.160 LAYER ME3 ;
 ANTENNADIFFAREA                          0.160 LAYER ME4 ;
 ANTENNAMAXAREACAR                       48.801 LAYER ME2 ;
 ANTENNAMAXAREACAR                       58.060 LAYER ME3 ;
 ANTENNAMAXAREACAR                       67.319 LAYER ME4 ;
END DI0
PIN VCC
  DIRECTION INOUT ;
  USE POWER ;
  SHAPE RING ;
 PORT
  LAYER ME4 ;
  RECT 2.000 547.210 1377.500 549.210 ;
  RECT 2.000 3.600 1377.500 5.600 ;
  RECT 1375.500 3.600 1377.500 549.210 ;
  RECT 2.000 3.600 4.000 549.210 ;
 END
END VCC
PIN GND
  DIRECTION INOUT ;
  USE GROUND ;
  SHAPE RING ;
 PORT
  LAYER ME3 ;
  RECT 0.000 549.210 1379.500 551.210 ;
  RECT 0.000 1.600 1379.500 3.600 ;
  RECT 1377.500 1.600 1379.500 551.210 ;
  RECT 0.000 1.600 2.000 551.210 ;
 END
END GND
OBS
  LAYER ME4 ;
  RECT 5.420 7.020 1374.080 545.790 ;
  RECT 1375.500 5.600 1377.500 547.210 ;
  RECT 2.000 5.600 4.000 547.210 ;
  RECT 4.000 547.210 1375.500 549.210 ;
  RECT 4.000 3.600 1375.500 5.600 ;
  RECT 2.000 547.210 4.000 549.210 ;
  RECT 1375.500 3.600 1377.500 5.600 ;
  RECT 1375.500 547.210 1377.500 549.210 ;
  RECT 2.000 3.600 4.000 5.600 ;
  RECT 1367.600 0.000 1368.400 1.000 ;
  RECT 1352.800 0.000 1353.600 1.000 ;
  RECT 1347.600 0.000 1348.400 1.000 ;
  RECT 1333.200 0.000 1334.000 1.000 ;
  RECT 1326.800 0.000 1327.600 1.000 ;
  RECT 1312.000 0.000 1312.800 1.000 ;
  RECT 1306.800 0.000 1307.600 1.000 ;
  RECT 1292.000 0.000 1292.800 1.000 ;
  RECT 1285.600 0.000 1286.400 1.000 ;
  RECT 1271.200 0.000 1272.000 1.000 ;
  RECT 1266.000 0.000 1266.800 1.000 ;
  RECT 1251.200 0.000 1252.000 1.000 ;
  RECT 1244.800 0.000 1245.600 1.000 ;
  RECT 1230.000 0.000 1230.800 1.000 ;
  RECT 1224.800 0.000 1225.600 1.000 ;
  RECT 1212.000 0.000 1212.800 1.000 ;
  RECT 1210.400 0.000 1211.200 1.000 ;
  RECT 1204.000 0.000 1204.800 1.000 ;
  RECT 1189.200 0.000 1190.000 1.000 ;
  RECT 1184.000 0.000 1184.800 1.000 ;
  RECT 1169.200 0.000 1170.000 1.000 ;
  RECT 1162.800 0.000 1163.600 1.000 ;
  RECT 1148.400 0.000 1149.200 1.000 ;
  RECT 1143.200 0.000 1144.000 1.000 ;
  RECT 1128.400 0.000 1129.200 1.000 ;
  RECT 1122.000 0.000 1122.800 1.000 ;
  RECT 1107.200 0.000 1108.000 1.000 ;
  RECT 1102.000 0.000 1102.800 1.000 ;
  RECT 1087.600 0.000 1088.400 1.000 ;
  RECT 1081.200 0.000 1082.000 1.000 ;
  RECT 1066.400 0.000 1067.200 1.000 ;
  RECT 1061.200 0.000 1062.000 1.000 ;
  RECT 1048.400 0.000 1049.200 1.000 ;
  RECT 1046.800 0.000 1047.600 1.000 ;
  RECT 1040.000 0.000 1040.800 1.000 ;
  RECT 1025.600 0.000 1026.400 1.000 ;
  RECT 1020.400 0.000 1021.200 1.000 ;
  RECT 1005.600 0.000 1006.400 1.000 ;
  RECT 999.200 0.000 1000.000 1.000 ;
  RECT 984.800 0.000 985.600 1.000 ;
  RECT 979.600 0.000 980.400 1.000 ;
  RECT 964.800 0.000 965.600 1.000 ;
  RECT 958.400 0.000 959.200 1.000 ;
  RECT 943.600 0.000 944.400 1.000 ;
  RECT 938.400 0.000 939.200 1.000 ;
  RECT 924.000 0.000 924.800 1.000 ;
  RECT 917.600 0.000 918.400 1.000 ;
  RECT 902.800 0.000 903.600 1.000 ;
  RECT 897.600 0.000 898.400 1.000 ;
  RECT 884.800 0.000 885.600 1.000 ;
  RECT 882.800 0.000 883.600 1.000 ;
  RECT 876.400 0.000 877.200 1.000 ;
  RECT 862.000 0.000 862.800 1.000 ;
  RECT 856.800 0.000 857.600 1.000 ;
  RECT 842.000 0.000 842.800 1.000 ;
  RECT 835.600 0.000 836.400 1.000 ;
  RECT 820.800 0.000 821.600 1.000 ;
  RECT 815.600 0.000 816.400 1.000 ;
  RECT 801.200 0.000 802.000 1.000 ;
  RECT 794.800 0.000 795.600 1.000 ;
  RECT 780.000 0.000 780.800 1.000 ;
  RECT 774.800 0.000 775.600 1.000 ;
  RECT 760.000 0.000 760.800 1.000 ;
  RECT 753.600 0.000 754.400 1.000 ;
  RECT 739.200 0.000 740.000 1.000 ;
  RECT 734.000 0.000 734.800 1.000 ;
  RECT 720.800 0.000 721.600 1.000 ;
  RECT 719.200 0.000 720.000 1.000 ;
  RECT 698.400 0.000 699.200 1.000 ;
  RECT 697.200 0.000 698.000 1.000 ;
  RECT 696.000 0.000 696.800 1.000 ;
  RECT 694.800 0.000 695.600 1.000 ;
  RECT 693.600 0.000 694.400 1.000 ;
  RECT 692.400 0.000 693.200 1.000 ;
  RECT 686.400 0.000 687.200 1.000 ;
  RECT 679.200 0.000 680.000 1.000 ;
  RECT 676.800 0.000 677.600 1.000 ;
  RECT 674.000 0.000 674.800 1.000 ;
  RECT 671.200 0.000 672.000 1.000 ;
  RECT 670.000 0.000 670.800 1.000 ;
  RECT 667.200 0.000 668.000 1.000 ;
  RECT 666.000 0.000 666.800 1.000 ;
  RECT 663.200 0.000 664.000 1.000 ;
  RECT 656.400 0.000 657.200 1.000 ;
  RECT 642.000 0.000 642.800 1.000 ;
  RECT 636.400 0.000 637.200 1.000 ;
  RECT 622.000 0.000 622.800 1.000 ;
  RECT 615.600 0.000 616.400 1.000 ;
  RECT 600.800 0.000 601.600 1.000 ;
  RECT 595.600 0.000 596.400 1.000 ;
  RECT 581.200 0.000 582.000 1.000 ;
  RECT 574.400 0.000 575.200 1.000 ;
  RECT 560.000 0.000 560.800 1.000 ;
  RECT 554.800 0.000 555.600 1.000 ;
  RECT 540.000 0.000 540.800 1.000 ;
  RECT 533.600 0.000 534.400 1.000 ;
  RECT 519.200 0.000 520.000 1.000 ;
  RECT 514.000 0.000 514.800 1.000 ;
  RECT 500.800 0.000 501.600 1.000 ;
  RECT 499.200 0.000 500.000 1.000 ;
  RECT 492.800 0.000 493.600 1.000 ;
  RECT 478.000 0.000 478.800 1.000 ;
  RECT 472.800 0.000 473.600 1.000 ;
  RECT 458.400 0.000 459.200 1.000 ;
  RECT 452.000 0.000 452.800 1.000 ;
  RECT 437.200 0.000 438.000 1.000 ;
  RECT 432.000 0.000 432.800 1.000 ;
  RECT 417.200 0.000 418.000 1.000 ;
  RECT 410.800 0.000 411.600 1.000 ;
  RECT 396.400 0.000 397.200 1.000 ;
  RECT 391.200 0.000 392.000 1.000 ;
  RECT 376.400 0.000 377.200 1.000 ;
  RECT 370.000 0.000 370.800 1.000 ;
  RECT 355.200 0.000 356.000 1.000 ;
  RECT 350.000 0.000 350.800 1.000 ;
  RECT 337.200 0.000 338.000 1.000 ;
  RECT 335.600 0.000 336.400 1.000 ;
  RECT 329.200 0.000 330.000 1.000 ;
  RECT 314.400 0.000 315.200 1.000 ;
  RECT 309.200 0.000 310.000 1.000 ;
  RECT 294.800 0.000 295.600 1.000 ;
  RECT 288.000 0.000 288.800 1.000 ;
  RECT 273.600 0.000 274.400 1.000 ;
  RECT 268.400 0.000 269.200 1.000 ;
  RECT 253.600 0.000 254.400 1.000 ;
  RECT 247.200 0.000 248.000 1.000 ;
  RECT 232.800 0.000 233.600 1.000 ;
  RECT 227.200 0.000 228.000 1.000 ;
  RECT 212.800 0.000 213.600 1.000 ;
  RECT 206.400 0.000 207.200 1.000 ;
  RECT 191.600 0.000 192.400 1.000 ;
  RECT 186.400 0.000 187.200 1.000 ;
  RECT 173.600 0.000 174.400 1.000 ;
  RECT 172.000 0.000 172.800 1.000 ;
  RECT 165.200 0.000 166.000 1.000 ;
  RECT 150.800 0.000 151.600 1.000 ;
  RECT 145.600 0.000 146.400 1.000 ;
  RECT 130.800 0.000 131.600 1.000 ;
  RECT 124.400 0.000 125.200 1.000 ;
  RECT 110.000 0.000 110.800 1.000 ;
  RECT 104.800 0.000 105.600 1.000 ;
  RECT 90.000 0.000 90.800 1.000 ;
  RECT 83.600 0.000 84.400 1.000 ;
  RECT 68.800 0.000 69.600 1.000 ;
  RECT 63.600 0.000 64.400 1.000 ;
  RECT 49.200 0.000 50.000 1.000 ;
  RECT 42.800 0.000 43.600 1.000 ;
  RECT 28.000 0.000 28.800 1.000 ;
  RECT 22.800 0.000 23.600 1.000 ;
  RECT 10.000 0.000 10.800 1.000 ;
  RECT 8.000 0.000 8.800 1.000 ;
  RECT 1374.360 9.570 1375.500 11.170 ;
  RECT 1374.360 14.200 1375.500 15.200 ;
  RECT 1374.360 18.730 1375.500 19.730 ;
  RECT 1374.360 21.230 1375.500 22.070 ;
  RECT 1374.360 24.170 1375.500 25.170 ;
  RECT 1374.360 36.320 1375.500 37.320 ;
  RECT 1374.360 39.480 1375.500 40.080 ;
  RECT 1374.360 45.560 1375.500 46.160 ;
  RECT 1374.360 57.100 1375.500 61.420 ;
  RECT 1372.940 5.880 1374.080 7.020 ;
  RECT 729.500 5.600 737.500 7.020 ;
  RECT 719.460 5.880 727.460 7.020 ;
  RECT 739.300 5.880 747.300 7.020 ;
  RECT 749.340 5.600 757.340 7.020 ;
  RECT 760.380 5.880 768.380 7.020 ;
  RECT 770.420 5.600 778.420 7.020 ;
  RECT 780.220 5.880 788.220 7.020 ;
  RECT 790.260 5.600 798.260 7.020 ;
  RECT 801.300 5.880 809.300 7.020 ;
  RECT 811.340 5.600 819.340 7.020 ;
  RECT 821.140 5.880 829.140 7.020 ;
  RECT 831.180 5.600 839.180 7.020 ;
  RECT 842.220 5.880 850.220 7.020 ;
  RECT 852.260 5.600 860.260 7.020 ;
  RECT 862.060 5.880 870.060 7.020 ;
  RECT 872.100 5.600 880.100 7.020 ;
  RECT 893.180 5.600 901.180 7.020 ;
  RECT 883.140 5.880 891.140 7.020 ;
  RECT 902.980 5.880 910.980 7.020 ;
  RECT 913.020 5.600 921.020 7.020 ;
  RECT 924.060 5.880 932.060 7.020 ;
  RECT 934.100 5.600 942.100 7.020 ;
  RECT 943.900 5.880 951.900 7.020 ;
  RECT 953.940 5.600 961.940 7.020 ;
  RECT 964.980 5.880 972.980 7.020 ;
  RECT 975.020 5.600 983.020 7.020 ;
  RECT 984.820 5.880 992.820 7.020 ;
  RECT 994.860 5.600 1002.860 7.020 ;
  RECT 1005.900 5.880 1013.900 7.020 ;
  RECT 1015.940 5.600 1023.940 7.020 ;
  RECT 1025.740 5.880 1033.740 7.020 ;
  RECT 1035.780 5.600 1043.780 7.020 ;
  RECT 1056.860 5.600 1064.860 7.020 ;
  RECT 1046.820 5.880 1054.820 7.020 ;
  RECT 1066.660 5.880 1074.660 7.020 ;
  RECT 1076.700 5.600 1084.700 7.020 ;
  RECT 1087.740 5.880 1095.740 7.020 ;
  RECT 1097.780 5.600 1105.780 7.020 ;
  RECT 1107.580 5.880 1115.580 7.020 ;
  RECT 1117.620 5.600 1125.620 7.020 ;
  RECT 1128.660 5.880 1136.660 7.020 ;
  RECT 1138.700 5.600 1146.700 7.020 ;
  RECT 1148.500 5.880 1156.500 7.020 ;
  RECT 1158.540 5.600 1166.540 7.020 ;
  RECT 1169.580 5.880 1177.580 7.020 ;
  RECT 1179.620 5.600 1187.620 7.020 ;
  RECT 1189.420 5.880 1197.420 7.020 ;
  RECT 1199.460 5.600 1207.460 7.020 ;
  RECT 1220.540 5.600 1228.540 7.020 ;
  RECT 1210.500 5.880 1218.500 7.020 ;
  RECT 1230.340 5.880 1238.340 7.020 ;
  RECT 1240.380 5.600 1248.380 7.020 ;
  RECT 1251.420 5.880 1259.420 7.020 ;
  RECT 1261.460 5.600 1269.460 7.020 ;
  RECT 1271.260 5.880 1279.260 7.020 ;
  RECT 1281.300 5.600 1289.300 7.020 ;
  RECT 1292.340 5.880 1300.340 7.020 ;
  RECT 1302.380 5.600 1310.380 7.020 ;
  RECT 1312.180 5.880 1320.180 7.020 ;
  RECT 1322.220 5.600 1330.220 7.020 ;
  RECT 1333.260 5.880 1341.260 7.020 ;
  RECT 1343.300 5.600 1351.300 7.020 ;
  RECT 1353.100 5.880 1361.100 7.020 ;
  RECT 1363.140 5.600 1371.140 7.020 ;
  RECT 681.160 5.600 684.220 7.020 ;
  RECT 684.720 5.880 688.170 7.020 ;
  RECT 688.670 5.600 692.420 7.020 ;
  RECT 693.570 5.880 699.490 7.020 ;
  RECT 700.640 5.600 704.390 7.020 ;
  RECT 704.890 5.600 708.640 7.020 ;
  RECT 709.140 5.600 712.890 7.020 ;
  RECT 678.440 5.600 680.200 7.020 ;
  RECT 676.440 5.880 678.200 7.020 ;
  RECT 673.100 5.600 674.860 7.020 ;
  RECT 671.100 5.880 672.860 7.020 ;
  RECT 669.100 5.600 670.860 7.020 ;
  RECT 667.100 5.880 668.860 7.020 ;
  RECT 665.100 5.600 666.860 7.020 ;
  RECT 663.100 5.880 664.860 7.020 ;
  RECT 4.000 57.100 5.140 61.420 ;
  RECT 4.000 45.560 5.140 46.160 ;
  RECT 4.000 39.480 5.140 40.080 ;
  RECT 4.000 36.320 5.140 37.320 ;
  RECT 4.000 24.170 5.140 25.170 ;
  RECT 4.000 21.230 5.140 22.070 ;
  RECT 4.000 18.730 5.140 19.730 ;
  RECT 4.000 14.200 5.140 15.200 ;
  RECT 4.000 9.570 5.140 11.170 ;
  RECT 5.420 5.880 6.560 7.020 ;
  RECT 18.400 5.600 26.400 7.020 ;
  RECT 8.360 5.880 16.360 7.020 ;
  RECT 28.200 5.880 36.200 7.020 ;
  RECT 38.240 5.600 46.240 7.020 ;
  RECT 49.280 5.880 57.280 7.020 ;
  RECT 59.320 5.600 67.320 7.020 ;
  RECT 69.120 5.880 77.120 7.020 ;
  RECT 79.160 5.600 87.160 7.020 ;
  RECT 90.200 5.880 98.200 7.020 ;
  RECT 100.240 5.600 108.240 7.020 ;
  RECT 110.040 5.880 118.040 7.020 ;
  RECT 120.080 5.600 128.080 7.020 ;
  RECT 131.120 5.880 139.120 7.020 ;
  RECT 141.160 5.600 149.160 7.020 ;
  RECT 150.960 5.880 158.960 7.020 ;
  RECT 161.000 5.600 169.000 7.020 ;
  RECT 182.080 5.600 190.080 7.020 ;
  RECT 172.040 5.880 180.040 7.020 ;
  RECT 191.880 5.880 199.880 7.020 ;
  RECT 201.920 5.600 209.920 7.020 ;
  RECT 212.960 5.880 220.960 7.020 ;
  RECT 223.000 5.600 231.000 7.020 ;
  RECT 232.800 5.880 240.800 7.020 ;
  RECT 242.840 5.600 250.840 7.020 ;
  RECT 253.880 5.880 261.880 7.020 ;
  RECT 263.920 5.600 271.920 7.020 ;
  RECT 273.720 5.880 281.720 7.020 ;
  RECT 283.760 5.600 291.760 7.020 ;
  RECT 294.800 5.880 302.800 7.020 ;
  RECT 304.840 5.600 312.840 7.020 ;
  RECT 314.640 5.880 322.640 7.020 ;
  RECT 324.680 5.600 332.680 7.020 ;
  RECT 345.760 5.600 353.760 7.020 ;
  RECT 335.720 5.880 343.720 7.020 ;
  RECT 355.560 5.880 363.560 7.020 ;
  RECT 365.600 5.600 373.600 7.020 ;
  RECT 376.640 5.880 384.640 7.020 ;
  RECT 386.680 5.600 394.680 7.020 ;
  RECT 396.480 5.880 404.480 7.020 ;
  RECT 406.520 5.600 414.520 7.020 ;
  RECT 417.560 5.880 425.560 7.020 ;
  RECT 427.600 5.600 435.600 7.020 ;
  RECT 437.400 5.880 445.400 7.020 ;
  RECT 447.440 5.600 455.440 7.020 ;
  RECT 458.480 5.880 466.480 7.020 ;
  RECT 468.520 5.600 476.520 7.020 ;
  RECT 478.320 5.880 486.320 7.020 ;
  RECT 488.360 5.600 496.360 7.020 ;
  RECT 509.440 5.600 517.440 7.020 ;
  RECT 499.400 5.880 507.400 7.020 ;
  RECT 519.240 5.880 527.240 7.020 ;
  RECT 529.280 5.600 537.280 7.020 ;
  RECT 540.320 5.880 548.320 7.020 ;
  RECT 550.360 5.600 558.360 7.020 ;
  RECT 560.160 5.880 568.160 7.020 ;
  RECT 570.200 5.600 578.200 7.020 ;
  RECT 581.240 5.880 589.240 7.020 ;
  RECT 591.280 5.600 599.280 7.020 ;
  RECT 601.080 5.880 609.080 7.020 ;
  RECT 611.120 5.600 619.120 7.020 ;
  RECT 622.160 5.880 630.160 7.020 ;
  RECT 632.200 5.600 640.200 7.020 ;
  RECT 642.000 5.880 650.000 7.020 ;
  RECT 652.040 5.600 660.040 7.020 ;
  RECT 1374.360 545.220 1375.500 545.600 ;
  RECT 1374.360 537.300 1375.500 537.580 ;
  RECT 1374.360 533.620 1375.500 533.900 ;
  RECT 1374.360 529.940 1375.500 530.220 ;
  RECT 1374.360 526.260 1375.500 526.540 ;
  RECT 1374.360 522.580 1375.500 522.860 ;
  RECT 1374.360 518.900 1375.500 519.180 ;
  RECT 1374.360 515.220 1375.500 515.500 ;
  RECT 1374.360 511.540 1375.500 511.820 ;
  RECT 1374.360 507.860 1375.500 508.140 ;
  RECT 1374.360 504.180 1375.500 504.460 ;
  RECT 1374.360 500.500 1375.500 500.780 ;
  RECT 1374.360 496.820 1375.500 497.100 ;
  RECT 1374.360 493.140 1375.500 493.420 ;
  RECT 1374.360 489.460 1375.500 489.740 ;
  RECT 1374.360 485.780 1375.500 486.060 ;
  RECT 1374.360 482.100 1375.500 482.380 ;
  RECT 1374.360 478.420 1375.500 478.700 ;
  RECT 1374.360 474.740 1375.500 475.020 ;
  RECT 1374.360 471.060 1375.500 471.340 ;
  RECT 1374.360 467.380 1375.500 467.660 ;
  RECT 1374.360 463.700 1375.500 463.980 ;
  RECT 1374.360 460.020 1375.500 460.300 ;
  RECT 1374.360 456.340 1375.500 456.620 ;
  RECT 1374.360 452.660 1375.500 452.940 ;
  RECT 1374.360 448.980 1375.500 449.260 ;
  RECT 1374.360 445.300 1375.500 445.580 ;
  RECT 1374.360 441.620 1375.500 441.900 ;
  RECT 1374.360 437.940 1375.500 438.220 ;
  RECT 1374.360 434.260 1375.500 434.540 ;
  RECT 1374.360 430.580 1375.500 430.860 ;
  RECT 1374.360 426.900 1375.500 427.180 ;
  RECT 1374.360 423.220 1375.500 423.500 ;
  RECT 1374.360 419.540 1375.500 419.820 ;
  RECT 1374.360 415.860 1375.500 416.140 ;
  RECT 1374.360 412.180 1375.500 412.460 ;
  RECT 1374.360 408.500 1375.500 408.780 ;
  RECT 1374.360 404.820 1375.500 405.100 ;
  RECT 1374.360 401.140 1375.500 401.420 ;
  RECT 1374.360 397.460 1375.500 397.740 ;
  RECT 1374.360 393.780 1375.500 394.060 ;
  RECT 1374.360 390.100 1375.500 390.380 ;
  RECT 1374.360 386.420 1375.500 386.700 ;
  RECT 1374.360 382.740 1375.500 383.020 ;
  RECT 1374.360 379.060 1375.500 379.340 ;
  RECT 1374.360 375.380 1375.500 375.660 ;
  RECT 1374.360 371.700 1375.500 371.980 ;
  RECT 1374.360 368.020 1375.500 368.300 ;
  RECT 1374.360 364.340 1375.500 364.620 ;
  RECT 1374.360 360.660 1375.500 360.940 ;
  RECT 1374.360 356.980 1375.500 357.260 ;
  RECT 1374.360 353.300 1375.500 353.580 ;
  RECT 1374.360 349.620 1375.500 349.900 ;
  RECT 1374.360 345.940 1375.500 346.220 ;
  RECT 1374.360 342.260 1375.500 342.540 ;
  RECT 1374.360 338.580 1375.500 338.860 ;
  RECT 1374.360 334.900 1375.500 335.180 ;
  RECT 1374.360 331.220 1375.500 331.500 ;
  RECT 1374.360 327.540 1375.500 327.820 ;
  RECT 1374.360 323.860 1375.500 324.140 ;
  RECT 1374.360 320.180 1375.500 320.460 ;
  RECT 1374.360 316.500 1375.500 316.780 ;
  RECT 1374.360 312.820 1375.500 313.100 ;
  RECT 1374.360 309.140 1375.500 309.420 ;
  RECT 1374.360 305.460 1375.500 305.740 ;
  RECT 1374.360 301.780 1375.500 302.060 ;
  RECT 1374.360 298.100 1375.500 298.380 ;
  RECT 1374.360 294.420 1375.500 294.700 ;
  RECT 1374.360 290.740 1375.500 291.020 ;
  RECT 1374.360 287.060 1375.500 287.340 ;
  RECT 1374.360 283.380 1375.500 283.660 ;
  RECT 1374.360 279.700 1375.500 279.980 ;
  RECT 1374.360 276.020 1375.500 276.300 ;
  RECT 1374.360 272.340 1375.500 272.620 ;
  RECT 1374.360 268.660 1375.500 268.940 ;
  RECT 1374.360 264.980 1375.500 265.260 ;
  RECT 1374.360 261.300 1375.500 261.580 ;
  RECT 1374.360 257.620 1375.500 257.900 ;
  RECT 1374.360 253.940 1375.500 254.220 ;
  RECT 1374.360 250.260 1375.500 250.540 ;
  RECT 1374.360 246.580 1375.500 246.860 ;
  RECT 1374.360 242.900 1375.500 243.180 ;
  RECT 1374.360 239.220 1375.500 239.500 ;
  RECT 1374.360 235.540 1375.500 235.820 ;
  RECT 1374.360 231.860 1375.500 232.140 ;
  RECT 1374.360 228.180 1375.500 228.460 ;
  RECT 1374.360 224.500 1375.500 224.780 ;
  RECT 1374.360 220.820 1375.500 221.100 ;
  RECT 1374.360 217.140 1375.500 217.420 ;
  RECT 1374.360 213.460 1375.500 213.740 ;
  RECT 1374.360 209.780 1375.500 210.060 ;
  RECT 1374.360 206.100 1375.500 206.380 ;
  RECT 1374.360 202.420 1375.500 202.700 ;
  RECT 1374.360 198.740 1375.500 199.020 ;
  RECT 1374.360 195.060 1375.500 195.340 ;
  RECT 1374.360 191.380 1375.500 191.660 ;
  RECT 1374.360 187.700 1375.500 187.980 ;
  RECT 1374.360 184.020 1375.500 184.300 ;
  RECT 1374.360 180.340 1375.500 180.620 ;
  RECT 1374.360 176.660 1375.500 176.940 ;
  RECT 1374.360 172.980 1375.500 173.260 ;
  RECT 1374.360 169.300 1375.500 169.580 ;
  RECT 1374.360 165.620 1375.500 165.900 ;
  RECT 1374.360 161.940 1375.500 162.220 ;
  RECT 1374.360 158.260 1375.500 158.540 ;
  RECT 1374.360 154.580 1375.500 154.860 ;
  RECT 1374.360 150.900 1375.500 151.180 ;
  RECT 1374.360 147.220 1375.500 147.500 ;
  RECT 1374.360 143.540 1375.500 143.820 ;
  RECT 1374.360 139.860 1375.500 140.140 ;
  RECT 1374.360 136.180 1375.500 136.460 ;
  RECT 1374.360 132.500 1375.500 132.780 ;
  RECT 1374.360 128.820 1375.500 129.100 ;
  RECT 1374.360 125.140 1375.500 125.420 ;
  RECT 1374.360 121.460 1375.500 121.740 ;
  RECT 1374.360 117.780 1375.500 118.060 ;
  RECT 1374.360 114.100 1375.500 114.380 ;
  RECT 1374.360 110.420 1375.500 110.700 ;
  RECT 1374.360 106.740 1375.500 107.020 ;
  RECT 1374.360 103.060 1375.500 103.340 ;
  RECT 1374.360 99.380 1375.500 99.660 ;
  RECT 1374.360 95.700 1375.500 95.980 ;
  RECT 1374.360 92.020 1375.500 92.300 ;
  RECT 1374.360 88.340 1375.500 88.620 ;
  RECT 1374.360 84.660 1375.500 84.940 ;
  RECT 1374.360 80.980 1375.500 81.260 ;
  RECT 1374.360 77.300 1375.500 77.580 ;
  RECT 1374.360 73.620 1375.500 73.900 ;
  RECT 1374.360 69.940 1375.500 70.220 ;
  RECT 1374.360 65.600 1375.500 65.980 ;
  RECT 718.100 546.070 718.350 547.210 ;
  RECT 759.020 546.070 759.270 547.210 ;
  RECT 799.940 546.070 800.190 547.210 ;
  RECT 840.860 546.070 841.110 547.210 ;
  RECT 881.780 546.070 882.030 547.210 ;
  RECT 922.700 546.070 922.950 547.210 ;
  RECT 963.620 546.070 963.870 547.210 ;
  RECT 1004.540 546.070 1004.790 547.210 ;
  RECT 1045.460 546.070 1045.710 547.210 ;
  RECT 1086.380 546.070 1086.630 547.210 ;
  RECT 1127.300 546.070 1127.550 547.210 ;
  RECT 1168.220 546.070 1168.470 547.210 ;
  RECT 1209.140 546.070 1209.390 547.210 ;
  RECT 1250.060 546.070 1250.310 547.210 ;
  RECT 1290.980 546.070 1291.230 547.210 ;
  RECT 1331.900 546.070 1332.150 547.210 ;
  RECT 701.090 546.070 703.600 547.210 ;
  RECT 688.670 546.070 691.060 547.210 ;
  RECT 681.160 546.070 684.220 547.210 ;
  RECT 705.340 546.070 708.190 547.210 ;
  RECT 709.640 546.070 712.890 547.210 ;
  RECT 678.440 546.070 680.200 547.210 ;
  RECT 673.100 546.070 674.860 547.210 ;
  RECT 669.100 546.070 670.860 547.210 ;
  RECT 665.100 546.070 666.860 547.210 ;
  RECT 4.000 65.600 5.140 65.980 ;
  RECT 4.000 69.940 5.140 70.220 ;
  RECT 4.000 73.620 5.140 73.900 ;
  RECT 4.000 77.300 5.140 77.580 ;
  RECT 4.000 80.980 5.140 81.260 ;
  RECT 4.000 84.660 5.140 84.940 ;
  RECT 4.000 88.340 5.140 88.620 ;
  RECT 4.000 92.020 5.140 92.300 ;
  RECT 4.000 95.700 5.140 95.980 ;
  RECT 4.000 99.380 5.140 99.660 ;
  RECT 4.000 103.060 5.140 103.340 ;
  RECT 4.000 106.740 5.140 107.020 ;
  RECT 4.000 110.420 5.140 110.700 ;
  RECT 4.000 114.100 5.140 114.380 ;
  RECT 4.000 117.780 5.140 118.060 ;
  RECT 4.000 121.460 5.140 121.740 ;
  RECT 4.000 125.140 5.140 125.420 ;
  RECT 4.000 128.820 5.140 129.100 ;
  RECT 4.000 132.500 5.140 132.780 ;
  RECT 4.000 136.180 5.140 136.460 ;
  RECT 4.000 139.860 5.140 140.140 ;
  RECT 4.000 143.540 5.140 143.820 ;
  RECT 4.000 147.220 5.140 147.500 ;
  RECT 4.000 150.900 5.140 151.180 ;
  RECT 4.000 154.580 5.140 154.860 ;
  RECT 4.000 158.260 5.140 158.540 ;
  RECT 4.000 161.940 5.140 162.220 ;
  RECT 4.000 165.620 5.140 165.900 ;
  RECT 4.000 169.300 5.140 169.580 ;
  RECT 4.000 172.980 5.140 173.260 ;
  RECT 4.000 176.660 5.140 176.940 ;
  RECT 4.000 180.340 5.140 180.620 ;
  RECT 4.000 184.020 5.140 184.300 ;
  RECT 4.000 187.700 5.140 187.980 ;
  RECT 4.000 191.380 5.140 191.660 ;
  RECT 4.000 195.060 5.140 195.340 ;
  RECT 4.000 198.740 5.140 199.020 ;
  RECT 4.000 202.420 5.140 202.700 ;
  RECT 4.000 206.100 5.140 206.380 ;
  RECT 4.000 209.780 5.140 210.060 ;
  RECT 4.000 213.460 5.140 213.740 ;
  RECT 4.000 217.140 5.140 217.420 ;
  RECT 4.000 220.820 5.140 221.100 ;
  RECT 4.000 224.500 5.140 224.780 ;
  RECT 4.000 228.180 5.140 228.460 ;
  RECT 4.000 231.860 5.140 232.140 ;
  RECT 4.000 235.540 5.140 235.820 ;
  RECT 4.000 239.220 5.140 239.500 ;
  RECT 4.000 242.900 5.140 243.180 ;
  RECT 4.000 246.580 5.140 246.860 ;
  RECT 4.000 250.260 5.140 250.540 ;
  RECT 4.000 253.940 5.140 254.220 ;
  RECT 4.000 257.620 5.140 257.900 ;
  RECT 4.000 261.300 5.140 261.580 ;
  RECT 4.000 264.980 5.140 265.260 ;
  RECT 4.000 268.660 5.140 268.940 ;
  RECT 4.000 272.340 5.140 272.620 ;
  RECT 4.000 276.020 5.140 276.300 ;
  RECT 4.000 279.700 5.140 279.980 ;
  RECT 4.000 283.380 5.140 283.660 ;
  RECT 4.000 287.060 5.140 287.340 ;
  RECT 4.000 290.740 5.140 291.020 ;
  RECT 4.000 294.420 5.140 294.700 ;
  RECT 4.000 298.100 5.140 298.380 ;
  RECT 4.000 301.780 5.140 302.060 ;
  RECT 4.000 305.460 5.140 305.740 ;
  RECT 4.000 309.140 5.140 309.420 ;
  RECT 4.000 312.820 5.140 313.100 ;
  RECT 4.000 316.500 5.140 316.780 ;
  RECT 4.000 320.180 5.140 320.460 ;
  RECT 4.000 323.860 5.140 324.140 ;
  RECT 4.000 327.540 5.140 327.820 ;
  RECT 4.000 331.220 5.140 331.500 ;
  RECT 4.000 334.900 5.140 335.180 ;
  RECT 4.000 338.580 5.140 338.860 ;
  RECT 4.000 342.260 5.140 342.540 ;
  RECT 4.000 345.940 5.140 346.220 ;
  RECT 4.000 349.620 5.140 349.900 ;
  RECT 4.000 353.300 5.140 353.580 ;
  RECT 4.000 356.980 5.140 357.260 ;
  RECT 4.000 360.660 5.140 360.940 ;
  RECT 4.000 364.340 5.140 364.620 ;
  RECT 4.000 368.020 5.140 368.300 ;
  RECT 4.000 371.700 5.140 371.980 ;
  RECT 4.000 375.380 5.140 375.660 ;
  RECT 4.000 379.060 5.140 379.340 ;
  RECT 4.000 382.740 5.140 383.020 ;
  RECT 4.000 386.420 5.140 386.700 ;
  RECT 4.000 390.100 5.140 390.380 ;
  RECT 4.000 393.780 5.140 394.060 ;
  RECT 4.000 397.460 5.140 397.740 ;
  RECT 4.000 401.140 5.140 401.420 ;
  RECT 4.000 404.820 5.140 405.100 ;
  RECT 4.000 408.500 5.140 408.780 ;
  RECT 4.000 412.180 5.140 412.460 ;
  RECT 4.000 415.860 5.140 416.140 ;
  RECT 4.000 419.540 5.140 419.820 ;
  RECT 4.000 423.220 5.140 423.500 ;
  RECT 4.000 426.900 5.140 427.180 ;
  RECT 4.000 430.580 5.140 430.860 ;
  RECT 4.000 434.260 5.140 434.540 ;
  RECT 4.000 437.940 5.140 438.220 ;
  RECT 4.000 441.620 5.140 441.900 ;
  RECT 4.000 445.300 5.140 445.580 ;
  RECT 4.000 448.980 5.140 449.260 ;
  RECT 4.000 452.660 5.140 452.940 ;
  RECT 4.000 456.340 5.140 456.620 ;
  RECT 4.000 460.020 5.140 460.300 ;
  RECT 4.000 463.700 5.140 463.980 ;
  RECT 4.000 467.380 5.140 467.660 ;
  RECT 4.000 471.060 5.140 471.340 ;
  RECT 4.000 474.740 5.140 475.020 ;
  RECT 4.000 478.420 5.140 478.700 ;
  RECT 4.000 482.100 5.140 482.380 ;
  RECT 4.000 485.780 5.140 486.060 ;
  RECT 4.000 489.460 5.140 489.740 ;
  RECT 4.000 493.140 5.140 493.420 ;
  RECT 4.000 496.820 5.140 497.100 ;
  RECT 4.000 500.500 5.140 500.780 ;
  RECT 4.000 504.180 5.140 504.460 ;
  RECT 4.000 507.860 5.140 508.140 ;
  RECT 4.000 511.540 5.140 511.820 ;
  RECT 4.000 515.220 5.140 515.500 ;
  RECT 4.000 518.900 5.140 519.180 ;
  RECT 4.000 522.580 5.140 522.860 ;
  RECT 4.000 526.260 5.140 526.540 ;
  RECT 4.000 529.940 5.140 530.220 ;
  RECT 4.000 533.620 5.140 533.900 ;
  RECT 4.000 537.300 5.140 537.580 ;
  RECT 4.000 545.220 5.140 545.600 ;
  RECT 47.350 546.070 47.600 547.210 ;
  RECT 88.270 546.070 88.520 547.210 ;
  RECT 129.190 546.070 129.440 547.210 ;
  RECT 170.110 546.070 170.360 547.210 ;
  RECT 211.030 546.070 211.280 547.210 ;
  RECT 251.950 546.070 252.200 547.210 ;
  RECT 292.870 546.070 293.120 547.210 ;
  RECT 333.790 546.070 334.040 547.210 ;
  RECT 374.710 546.070 374.960 547.210 ;
  RECT 415.630 546.070 415.880 547.210 ;
  RECT 456.550 546.070 456.800 547.210 ;
  RECT 497.470 546.070 497.720 547.210 ;
  RECT 538.390 546.070 538.640 547.210 ;
  RECT 579.310 546.070 579.560 547.210 ;
  RECT 620.230 546.070 620.480 547.210 ;
  RECT 2.000 547.210 1377.500 549.210 ;
  RECT 2.000 3.600 1377.500 5.600 ;
  RECT 1375.500 3.600 1377.500 549.210 ;
  RECT 2.000 3.600 4.000 549.210 ;
  LAYER ME3 ;
  RECT 5.420 7.020 1374.080 545.790 ;
  RECT 1377.500 3.600 1379.500 549.210 ;
  RECT 0.000 3.600 2.000 549.210 ;
  RECT 2.000 549.210 1377.500 551.210 ;
  RECT 2.000 1.600 1377.500 3.600 ;
  RECT 1375.500 540.280 1377.220 547.210 ;
  RECT 1375.500 64.930 1377.220 67.240 ;
  RECT 1375.500 44.080 1377.220 61.260 ;
  RECT 1375.500 39.620 1377.220 41.480 ;
  RECT 1375.500 29.870 1377.220 33.520 ;
  RECT 1375.500 24.270 1377.220 26.870 ;
  RECT 1375.500 18.130 1377.220 21.270 ;
  RECT 1375.500 5.600 1377.220 11.230 ;
  RECT 2.280 540.280 4.000 547.210 ;
  RECT 2.280 64.930 4.000 67.240 ;
  RECT 2.280 44.080 4.000 61.260 ;
  RECT 2.280 39.620 4.000 41.480 ;
  RECT 2.280 29.870 4.000 33.520 ;
  RECT 2.280 24.270 4.000 26.870 ;
  RECT 2.280 18.130 4.000 21.270 ;
  RECT 2.280 5.600 4.000 11.230 ;
  RECT 1332.580 547.210 1375.500 548.930 ;
  RECT 1291.660 547.210 1330.330 548.930 ;
  RECT 1250.740 547.210 1289.410 548.930 ;
  RECT 1209.820 547.210 1248.490 548.930 ;
  RECT 1168.900 547.210 1207.570 548.930 ;
  RECT 1127.980 547.210 1166.650 548.930 ;
  RECT 1087.060 547.210 1125.730 548.930 ;
  RECT 1046.140 547.210 1084.810 548.930 ;
  RECT 1005.220 547.210 1043.890 548.930 ;
  RECT 964.300 547.210 1002.970 548.930 ;
  RECT 923.380 547.210 962.050 548.930 ;
  RECT 882.460 547.210 921.130 548.930 ;
  RECT 841.540 547.210 880.210 548.930 ;
  RECT 800.620 547.210 839.290 548.930 ;
  RECT 759.700 547.210 798.370 548.930 ;
  RECT 718.780 547.210 757.450 548.930 ;
  RECT 700.040 547.210 713.040 548.930 ;
  RECT 688.910 547.210 693.720 548.930 ;
  RECT 679.200 547.210 683.720 548.930 ;
  RECT 673.860 547.210 675.440 548.930 ;
  RECT 622.050 547.210 661.080 548.930 ;
  RECT 581.130 547.210 619.800 548.930 ;
  RECT 540.210 547.210 578.880 548.930 ;
  RECT 499.290 547.210 537.960 548.930 ;
  RECT 458.370 547.210 497.040 548.930 ;
  RECT 417.450 547.210 456.120 548.930 ;
  RECT 376.530 547.210 415.200 548.930 ;
  RECT 335.610 547.210 374.280 548.930 ;
  RECT 294.690 547.210 333.360 548.930 ;
  RECT 253.770 547.210 292.440 548.930 ;
  RECT 212.850 547.210 251.520 548.930 ;
  RECT 171.930 547.210 210.600 548.930 ;
  RECT 131.010 547.210 169.680 548.930 ;
  RECT 90.090 547.210 128.760 548.930 ;
  RECT 49.170 547.210 87.840 548.930 ;
  RECT 4.000 547.210 46.920 548.930 ;
  RECT 1362.100 3.880 1371.940 5.600 ;
  RECT 1342.260 3.880 1352.100 5.600 ;
  RECT 1321.180 3.880 1332.260 5.600 ;
  RECT 1301.340 3.880 1311.180 5.600 ;
  RECT 1280.260 3.880 1291.340 5.600 ;
  RECT 1260.420 3.880 1270.260 5.600 ;
  RECT 1239.340 3.880 1250.420 5.600 ;
  RECT 1219.500 3.880 1229.340 5.600 ;
  RECT 1198.420 3.880 1209.500 5.600 ;
  RECT 1178.580 3.880 1188.420 5.600 ;
  RECT 1157.500 3.880 1168.580 5.600 ;
  RECT 1137.660 3.880 1147.500 5.600 ;
  RECT 1116.580 3.880 1127.660 5.600 ;
  RECT 1096.740 3.880 1106.580 5.600 ;
  RECT 1075.660 3.880 1086.740 5.600 ;
  RECT 1055.820 3.880 1065.660 5.600 ;
  RECT 1034.740 3.880 1045.820 5.600 ;
  RECT 1014.900 3.880 1024.740 5.600 ;
  RECT 993.820 3.880 1004.900 5.600 ;
  RECT 973.980 3.880 983.820 5.600 ;
  RECT 952.900 3.880 963.980 5.600 ;
  RECT 933.060 3.880 942.900 5.600 ;
  RECT 911.980 3.880 923.060 5.600 ;
  RECT 892.140 3.880 901.980 5.600 ;
  RECT 871.060 3.880 882.140 5.600 ;
  RECT 851.220 3.880 861.060 5.600 ;
  RECT 830.140 3.880 841.220 5.600 ;
  RECT 810.300 3.880 820.140 5.600 ;
  RECT 789.220 3.880 800.300 5.600 ;
  RECT 769.380 3.880 779.220 5.600 ;
  RECT 748.300 3.880 759.380 5.600 ;
  RECT 728.460 3.880 738.300 5.600 ;
  RECT 700.490 3.880 718.460 5.600 ;
  RECT 689.170 3.880 692.570 5.600 ;
  RECT 679.200 3.880 683.720 5.600 ;
  RECT 673.860 3.880 675.440 5.600 ;
  RECT 651.000 3.880 662.100 5.600 ;
  RECT 631.160 3.880 641.000 5.600 ;
  RECT 610.080 3.880 621.160 5.600 ;
  RECT 590.240 3.880 600.080 5.600 ;
  RECT 569.160 3.880 580.240 5.600 ;
  RECT 549.320 3.880 559.160 5.600 ;
  RECT 528.240 3.880 539.320 5.600 ;
  RECT 508.400 3.880 518.240 5.600 ;
  RECT 487.320 3.880 498.400 5.600 ;
  RECT 467.480 3.880 477.320 5.600 ;
  RECT 446.400 3.880 457.480 5.600 ;
  RECT 426.560 3.880 436.400 5.600 ;
  RECT 405.480 3.880 416.560 5.600 ;
  RECT 385.640 3.880 395.480 5.600 ;
  RECT 364.560 3.880 375.640 5.600 ;
  RECT 344.720 3.880 354.560 5.600 ;
  RECT 323.640 3.880 334.720 5.600 ;
  RECT 303.800 3.880 313.640 5.600 ;
  RECT 282.720 3.880 293.800 5.600 ;
  RECT 262.880 3.880 272.720 5.600 ;
  RECT 241.800 3.880 252.880 5.600 ;
  RECT 221.960 3.880 231.800 5.600 ;
  RECT 200.880 3.880 211.960 5.600 ;
  RECT 181.040 3.880 190.880 5.600 ;
  RECT 159.960 3.880 171.040 5.600 ;
  RECT 140.120 3.880 149.960 5.600 ;
  RECT 119.040 3.880 130.120 5.600 ;
  RECT 99.200 3.880 109.040 5.600 ;
  RECT 78.120 3.880 89.200 5.600 ;
  RECT 58.280 3.880 68.120 5.600 ;
  RECT 37.200 3.880 48.280 5.600 ;
  RECT 17.360 3.880 27.200 5.600 ;
  RECT 2.280 547.210 4.000 548.930 ;
  RECT 0.000 549.210 2.000 551.210 ;
  RECT 1375.500 3.880 1377.220 5.600 ;
  RECT 1377.500 1.600 1379.500 3.600 ;
  RECT 1375.500 547.210 1377.220 548.930 ;
  RECT 1377.500 549.210 1379.500 551.210 ;
  RECT 2.280 3.880 4.000 5.600 ;
  RECT 0.000 1.600 2.000 3.600 ;
  RECT 1367.600 0.000 1368.400 1.000 ;
  RECT 1352.800 0.000 1353.600 1.000 ;
  RECT 1347.600 0.000 1348.400 1.000 ;
  RECT 1333.200 0.000 1334.000 1.000 ;
  RECT 1326.800 0.000 1327.600 1.000 ;
  RECT 1312.000 0.000 1312.800 1.000 ;
  RECT 1306.800 0.000 1307.600 1.000 ;
  RECT 1292.000 0.000 1292.800 1.000 ;
  RECT 1285.600 0.000 1286.400 1.000 ;
  RECT 1271.200 0.000 1272.000 1.000 ;
  RECT 1266.000 0.000 1266.800 1.000 ;
  RECT 1251.200 0.000 1252.000 1.000 ;
  RECT 1244.800 0.000 1245.600 1.000 ;
  RECT 1230.000 0.000 1230.800 1.000 ;
  RECT 1224.800 0.000 1225.600 1.000 ;
  RECT 1212.000 0.000 1212.800 1.000 ;
  RECT 1210.400 0.000 1211.200 1.000 ;
  RECT 1204.000 0.000 1204.800 1.000 ;
  RECT 1189.200 0.000 1190.000 1.000 ;
  RECT 1184.000 0.000 1184.800 1.000 ;
  RECT 1169.200 0.000 1170.000 1.000 ;
  RECT 1162.800 0.000 1163.600 1.000 ;
  RECT 1148.400 0.000 1149.200 1.000 ;
  RECT 1143.200 0.000 1144.000 1.000 ;
  RECT 1128.400 0.000 1129.200 1.000 ;
  RECT 1122.000 0.000 1122.800 1.000 ;
  RECT 1107.200 0.000 1108.000 1.000 ;
  RECT 1102.000 0.000 1102.800 1.000 ;
  RECT 1087.600 0.000 1088.400 1.000 ;
  RECT 1081.200 0.000 1082.000 1.000 ;
  RECT 1066.400 0.000 1067.200 1.000 ;
  RECT 1061.200 0.000 1062.000 1.000 ;
  RECT 1048.400 0.000 1049.200 1.000 ;
  RECT 1046.800 0.000 1047.600 1.000 ;
  RECT 1040.000 0.000 1040.800 1.000 ;
  RECT 1025.600 0.000 1026.400 1.000 ;
  RECT 1020.400 0.000 1021.200 1.000 ;
  RECT 1005.600 0.000 1006.400 1.000 ;
  RECT 999.200 0.000 1000.000 1.000 ;
  RECT 984.800 0.000 985.600 1.000 ;
  RECT 979.600 0.000 980.400 1.000 ;
  RECT 964.800 0.000 965.600 1.000 ;
  RECT 958.400 0.000 959.200 1.000 ;
  RECT 943.600 0.000 944.400 1.000 ;
  RECT 938.400 0.000 939.200 1.000 ;
  RECT 924.000 0.000 924.800 1.000 ;
  RECT 917.600 0.000 918.400 1.000 ;
  RECT 902.800 0.000 903.600 1.000 ;
  RECT 897.600 0.000 898.400 1.000 ;
  RECT 884.800 0.000 885.600 1.000 ;
  RECT 882.800 0.000 883.600 1.000 ;
  RECT 876.400 0.000 877.200 1.000 ;
  RECT 862.000 0.000 862.800 1.000 ;
  RECT 856.800 0.000 857.600 1.000 ;
  RECT 842.000 0.000 842.800 1.000 ;
  RECT 835.600 0.000 836.400 1.000 ;
  RECT 820.800 0.000 821.600 1.000 ;
  RECT 815.600 0.000 816.400 1.000 ;
  RECT 801.200 0.000 802.000 1.000 ;
  RECT 794.800 0.000 795.600 1.000 ;
  RECT 780.000 0.000 780.800 1.000 ;
  RECT 774.800 0.000 775.600 1.000 ;
  RECT 760.000 0.000 760.800 1.000 ;
  RECT 753.600 0.000 754.400 1.000 ;
  RECT 739.200 0.000 740.000 1.000 ;
  RECT 734.000 0.000 734.800 1.000 ;
  RECT 720.800 0.000 721.600 1.000 ;
  RECT 719.200 0.000 720.000 1.000 ;
  RECT 698.400 0.000 699.200 1.000 ;
  RECT 697.200 0.000 698.000 1.000 ;
  RECT 696.000 0.000 696.800 1.000 ;
  RECT 694.800 0.000 695.600 1.000 ;
  RECT 693.600 0.000 694.400 1.000 ;
  RECT 692.400 0.000 693.200 1.000 ;
  RECT 686.400 0.000 687.200 1.000 ;
  RECT 679.200 0.000 680.000 1.000 ;
  RECT 676.800 0.000 677.600 1.000 ;
  RECT 674.000 0.000 674.800 1.000 ;
  RECT 671.200 0.000 672.000 1.000 ;
  RECT 670.000 0.000 670.800 1.000 ;
  RECT 667.200 0.000 668.000 1.000 ;
  RECT 666.000 0.000 666.800 1.000 ;
  RECT 663.200 0.000 664.000 1.000 ;
  RECT 656.400 0.000 657.200 1.000 ;
  RECT 642.000 0.000 642.800 1.000 ;
  RECT 636.400 0.000 637.200 1.000 ;
  RECT 622.000 0.000 622.800 1.000 ;
  RECT 615.600 0.000 616.400 1.000 ;
  RECT 600.800 0.000 601.600 1.000 ;
  RECT 595.600 0.000 596.400 1.000 ;
  RECT 581.200 0.000 582.000 1.000 ;
  RECT 574.400 0.000 575.200 1.000 ;
  RECT 560.000 0.000 560.800 1.000 ;
  RECT 554.800 0.000 555.600 1.000 ;
  RECT 540.000 0.000 540.800 1.000 ;
  RECT 533.600 0.000 534.400 1.000 ;
  RECT 519.200 0.000 520.000 1.000 ;
  RECT 514.000 0.000 514.800 1.000 ;
  RECT 500.800 0.000 501.600 1.000 ;
  RECT 499.200 0.000 500.000 1.000 ;
  RECT 492.800 0.000 493.600 1.000 ;
  RECT 478.000 0.000 478.800 1.000 ;
  RECT 472.800 0.000 473.600 1.000 ;
  RECT 458.400 0.000 459.200 1.000 ;
  RECT 452.000 0.000 452.800 1.000 ;
  RECT 437.200 0.000 438.000 1.000 ;
  RECT 432.000 0.000 432.800 1.000 ;
  RECT 417.200 0.000 418.000 1.000 ;
  RECT 410.800 0.000 411.600 1.000 ;
  RECT 396.400 0.000 397.200 1.000 ;
  RECT 391.200 0.000 392.000 1.000 ;
  RECT 376.400 0.000 377.200 1.000 ;
  RECT 370.000 0.000 370.800 1.000 ;
  RECT 355.200 0.000 356.000 1.000 ;
  RECT 350.000 0.000 350.800 1.000 ;
  RECT 337.200 0.000 338.000 1.000 ;
  RECT 335.600 0.000 336.400 1.000 ;
  RECT 329.200 0.000 330.000 1.000 ;
  RECT 314.400 0.000 315.200 1.000 ;
  RECT 309.200 0.000 310.000 1.000 ;
  RECT 294.800 0.000 295.600 1.000 ;
  RECT 288.000 0.000 288.800 1.000 ;
  RECT 273.600 0.000 274.400 1.000 ;
  RECT 268.400 0.000 269.200 1.000 ;
  RECT 253.600 0.000 254.400 1.000 ;
  RECT 247.200 0.000 248.000 1.000 ;
  RECT 232.800 0.000 233.600 1.000 ;
  RECT 227.200 0.000 228.000 1.000 ;
  RECT 212.800 0.000 213.600 1.000 ;
  RECT 206.400 0.000 207.200 1.000 ;
  RECT 191.600 0.000 192.400 1.000 ;
  RECT 186.400 0.000 187.200 1.000 ;
  RECT 173.600 0.000 174.400 1.000 ;
  RECT 172.000 0.000 172.800 1.000 ;
  RECT 165.200 0.000 166.000 1.000 ;
  RECT 150.800 0.000 151.600 1.000 ;
  RECT 145.600 0.000 146.400 1.000 ;
  RECT 130.800 0.000 131.600 1.000 ;
  RECT 124.400 0.000 125.200 1.000 ;
  RECT 110.000 0.000 110.800 1.000 ;
  RECT 104.800 0.000 105.600 1.000 ;
  RECT 90.000 0.000 90.800 1.000 ;
  RECT 83.600 0.000 84.400 1.000 ;
  RECT 68.800 0.000 69.600 1.000 ;
  RECT 63.600 0.000 64.400 1.000 ;
  RECT 49.200 0.000 50.000 1.000 ;
  RECT 42.800 0.000 43.600 1.000 ;
  RECT 28.000 0.000 28.800 1.000 ;
  RECT 22.800 0.000 23.600 1.000 ;
  RECT 10.000 0.000 10.800 1.000 ;
  RECT 8.000 0.000 8.800 1.000 ;
  RECT 1374.080 62.260 1377.500 63.930 ;
  RECT 1374.080 22.270 1377.500 23.270 ;
  RECT 1374.080 16.130 1377.500 17.130 ;
  RECT 1374.080 12.230 1377.500 13.230 ;
  RECT 1374.080 27.870 1377.500 28.870 ;
  RECT 1374.080 42.480 1377.500 43.080 ;
  RECT 1374.080 37.620 1377.500 38.620 ;
  RECT 1374.080 34.520 1377.500 36.020 ;
  RECT 1374.360 9.570 1375.220 11.170 ;
  RECT 1374.360 14.200 1375.220 15.200 ;
  RECT 1374.360 18.730 1375.220 19.730 ;
  RECT 1374.360 21.230 1375.220 22.070 ;
  RECT 1374.360 24.170 1375.220 25.170 ;
  RECT 1374.360 36.320 1375.220 37.320 ;
  RECT 1374.360 39.480 1375.220 40.080 ;
  RECT 1374.360 45.560 1375.220 46.160 ;
  RECT 1374.360 57.100 1375.220 61.420 ;
  RECT 1372.940 3.600 1374.080 6.740 ;
  RECT 719.460 3.600 727.460 6.740 ;
  RECT 739.300 3.600 747.300 6.740 ;
  RECT 760.380 3.600 768.380 6.740 ;
  RECT 780.220 3.600 788.220 6.740 ;
  RECT 801.300 3.600 809.300 6.740 ;
  RECT 821.140 3.600 829.140 6.740 ;
  RECT 842.220 3.600 850.220 6.740 ;
  RECT 862.060 3.600 870.060 6.740 ;
  RECT 883.140 3.600 891.140 6.740 ;
  RECT 902.980 3.600 910.980 6.740 ;
  RECT 924.060 3.600 932.060 6.740 ;
  RECT 943.900 3.600 951.900 6.740 ;
  RECT 964.980 3.600 972.980 6.740 ;
  RECT 984.820 3.600 992.820 6.740 ;
  RECT 1005.900 3.600 1013.900 6.740 ;
  RECT 1025.740 3.600 1033.740 6.740 ;
  RECT 1046.820 3.600 1054.820 6.740 ;
  RECT 1066.660 3.600 1074.660 6.740 ;
  RECT 1087.740 3.600 1095.740 6.740 ;
  RECT 1107.580 3.600 1115.580 6.740 ;
  RECT 1128.660 3.600 1136.660 6.740 ;
  RECT 1148.500 3.600 1156.500 6.740 ;
  RECT 1169.580 3.600 1177.580 6.740 ;
  RECT 1189.420 3.600 1197.420 6.740 ;
  RECT 1210.500 3.600 1218.500 6.740 ;
  RECT 1230.340 3.600 1238.340 6.740 ;
  RECT 1251.420 3.600 1259.420 6.740 ;
  RECT 1271.260 3.600 1279.260 6.740 ;
  RECT 1292.340 3.600 1300.340 6.740 ;
  RECT 1312.180 3.600 1320.180 6.740 ;
  RECT 1333.260 3.600 1341.260 6.740 ;
  RECT 1353.100 3.600 1361.100 6.740 ;
  RECT 684.720 3.600 688.170 6.740 ;
  RECT 693.570 3.600 699.490 6.740 ;
  RECT 676.440 3.600 678.200 6.740 ;
  RECT 671.100 3.600 672.860 6.740 ;
  RECT 667.100 3.600 668.860 6.740 ;
  RECT 663.100 3.600 664.860 6.740 ;
  RECT 4.280 57.100 5.140 61.420 ;
  RECT 4.280 45.560 5.140 46.160 ;
  RECT 4.280 39.480 5.140 40.080 ;
  RECT 4.280 36.320 5.140 37.320 ;
  RECT 4.280 24.170 5.140 25.170 ;
  RECT 4.280 21.230 5.140 22.070 ;
  RECT 4.280 18.730 5.140 19.730 ;
  RECT 4.280 14.200 5.140 15.200 ;
  RECT 4.280 9.570 5.140 11.170 ;
  RECT 2.000 34.520 5.420 36.020 ;
  RECT 2.000 37.620 5.420 38.620 ;
  RECT 2.000 42.480 5.420 43.080 ;
  RECT 2.000 27.870 5.420 28.870 ;
  RECT 2.000 12.230 5.420 13.230 ;
  RECT 2.000 16.130 5.420 17.130 ;
  RECT 2.000 22.270 5.420 23.270 ;
  RECT 2.000 62.260 5.420 63.930 ;
  RECT 5.420 3.600 6.560 6.740 ;
  RECT 8.360 3.600 16.360 6.740 ;
  RECT 28.200 3.600 36.200 6.740 ;
  RECT 49.280 3.600 57.280 6.740 ;
  RECT 69.120 3.600 77.120 6.740 ;
  RECT 90.200 3.600 98.200 6.740 ;
  RECT 110.040 3.600 118.040 6.740 ;
  RECT 131.120 3.600 139.120 6.740 ;
  RECT 150.960 3.600 158.960 6.740 ;
  RECT 172.040 3.600 180.040 6.740 ;
  RECT 191.880 3.600 199.880 6.740 ;
  RECT 212.960 3.600 220.960 6.740 ;
  RECT 232.800 3.600 240.800 6.740 ;
  RECT 253.880 3.600 261.880 6.740 ;
  RECT 273.720 3.600 281.720 6.740 ;
  RECT 294.800 3.600 302.800 6.740 ;
  RECT 314.640 3.600 322.640 6.740 ;
  RECT 335.720 3.600 343.720 6.740 ;
  RECT 355.560 3.600 363.560 6.740 ;
  RECT 376.640 3.600 384.640 6.740 ;
  RECT 396.480 3.600 404.480 6.740 ;
  RECT 417.560 3.600 425.560 6.740 ;
  RECT 437.400 3.600 445.400 6.740 ;
  RECT 458.480 3.600 466.480 6.740 ;
  RECT 478.320 3.600 486.320 6.740 ;
  RECT 499.400 3.600 507.400 6.740 ;
  RECT 519.240 3.600 527.240 6.740 ;
  RECT 540.320 3.600 548.320 6.740 ;
  RECT 560.160 3.600 568.160 6.740 ;
  RECT 581.240 3.600 589.240 6.740 ;
  RECT 601.080 3.600 609.080 6.740 ;
  RECT 622.160 3.600 630.160 6.740 ;
  RECT 642.000 3.600 650.000 6.740 ;
  RECT 1374.360 545.220 1375.220 545.600 ;
  RECT 1374.360 537.300 1375.220 537.580 ;
  RECT 1374.080 538.080 1377.500 539.280 ;
  RECT 1374.080 535.600 1377.500 536.800 ;
  RECT 1374.360 533.620 1375.220 533.900 ;
  RECT 1374.080 534.400 1377.500 535.600 ;
  RECT 1374.080 531.920 1377.500 533.120 ;
  RECT 1374.360 529.940 1375.220 530.220 ;
  RECT 1374.080 530.720 1377.500 531.920 ;
  RECT 1374.080 528.240 1377.500 529.440 ;
  RECT 1374.360 526.260 1375.220 526.540 ;
  RECT 1374.080 527.040 1377.500 528.240 ;
  RECT 1374.080 524.560 1377.500 525.760 ;
  RECT 1374.360 522.580 1375.220 522.860 ;
  RECT 1374.080 523.360 1377.500 524.560 ;
  RECT 1374.080 520.880 1377.500 522.080 ;
  RECT 1374.360 518.900 1375.220 519.180 ;
  RECT 1374.080 519.680 1377.500 520.880 ;
  RECT 1374.080 517.200 1377.500 518.400 ;
  RECT 1374.360 515.220 1375.220 515.500 ;
  RECT 1374.080 516.000 1377.500 517.200 ;
  RECT 1374.080 513.520 1377.500 514.720 ;
  RECT 1374.360 511.540 1375.220 511.820 ;
  RECT 1374.080 512.320 1377.500 513.520 ;
  RECT 1374.080 509.840 1377.500 511.040 ;
  RECT 1374.360 507.860 1375.220 508.140 ;
  RECT 1374.080 508.640 1377.500 509.840 ;
  RECT 1374.080 506.160 1377.500 507.360 ;
  RECT 1374.360 504.180 1375.220 504.460 ;
  RECT 1374.080 504.960 1377.500 506.160 ;
  RECT 1374.080 502.480 1377.500 503.680 ;
  RECT 1374.360 500.500 1375.220 500.780 ;
  RECT 1374.080 501.280 1377.500 502.480 ;
  RECT 1374.080 498.800 1377.500 500.000 ;
  RECT 1374.360 496.820 1375.220 497.100 ;
  RECT 1374.080 497.600 1377.500 498.800 ;
  RECT 1374.080 495.120 1377.500 496.320 ;
  RECT 1374.360 493.140 1375.220 493.420 ;
  RECT 1374.080 493.920 1377.500 495.120 ;
  RECT 1374.080 491.440 1377.500 492.640 ;
  RECT 1374.360 489.460 1375.220 489.740 ;
  RECT 1374.080 490.240 1377.500 491.440 ;
  RECT 1374.080 487.760 1377.500 488.960 ;
  RECT 1374.360 485.780 1375.220 486.060 ;
  RECT 1374.080 486.560 1377.500 487.760 ;
  RECT 1374.080 484.080 1377.500 485.280 ;
  RECT 1374.360 482.100 1375.220 482.380 ;
  RECT 1374.080 482.880 1377.500 484.080 ;
  RECT 1374.080 480.400 1377.500 481.600 ;
  RECT 1374.360 478.420 1375.220 478.700 ;
  RECT 1374.080 479.200 1377.500 480.400 ;
  RECT 1374.080 476.720 1377.500 477.920 ;
  RECT 1374.360 474.740 1375.220 475.020 ;
  RECT 1374.080 475.520 1377.500 476.720 ;
  RECT 1374.080 473.040 1377.500 474.240 ;
  RECT 1374.360 471.060 1375.220 471.340 ;
  RECT 1374.080 471.840 1377.500 473.040 ;
  RECT 1374.080 469.360 1377.500 470.560 ;
  RECT 1374.360 467.380 1375.220 467.660 ;
  RECT 1374.080 468.160 1377.500 469.360 ;
  RECT 1374.080 465.680 1377.500 466.880 ;
  RECT 1374.360 463.700 1375.220 463.980 ;
  RECT 1374.080 464.480 1377.500 465.680 ;
  RECT 1374.080 462.000 1377.500 463.200 ;
  RECT 1374.360 460.020 1375.220 460.300 ;
  RECT 1374.080 460.800 1377.500 462.000 ;
  RECT 1374.080 458.320 1377.500 459.520 ;
  RECT 1374.360 456.340 1375.220 456.620 ;
  RECT 1374.080 457.120 1377.500 458.320 ;
  RECT 1374.080 454.640 1377.500 455.840 ;
  RECT 1374.360 452.660 1375.220 452.940 ;
  RECT 1374.080 453.440 1377.500 454.640 ;
  RECT 1374.080 450.960 1377.500 452.160 ;
  RECT 1374.360 448.980 1375.220 449.260 ;
  RECT 1374.080 449.760 1377.500 450.960 ;
  RECT 1374.080 447.280 1377.500 448.480 ;
  RECT 1374.360 445.300 1375.220 445.580 ;
  RECT 1374.080 446.080 1377.500 447.280 ;
  RECT 1374.080 443.600 1377.500 444.800 ;
  RECT 1374.360 441.620 1375.220 441.900 ;
  RECT 1374.080 442.400 1377.500 443.600 ;
  RECT 1374.080 439.920 1377.500 441.120 ;
  RECT 1374.360 437.940 1375.220 438.220 ;
  RECT 1374.080 438.720 1377.500 439.920 ;
  RECT 1374.080 436.240 1377.500 437.440 ;
  RECT 1374.360 434.260 1375.220 434.540 ;
  RECT 1374.080 435.040 1377.500 436.240 ;
  RECT 1374.080 432.560 1377.500 433.760 ;
  RECT 1374.360 430.580 1375.220 430.860 ;
  RECT 1374.080 431.360 1377.500 432.560 ;
  RECT 1374.080 428.880 1377.500 430.080 ;
  RECT 1374.360 426.900 1375.220 427.180 ;
  RECT 1374.080 427.680 1377.500 428.880 ;
  RECT 1374.080 425.200 1377.500 426.400 ;
  RECT 1374.360 423.220 1375.220 423.500 ;
  RECT 1374.080 424.000 1377.500 425.200 ;
  RECT 1374.080 421.520 1377.500 422.720 ;
  RECT 1374.360 419.540 1375.220 419.820 ;
  RECT 1374.080 420.320 1377.500 421.520 ;
  RECT 1374.080 417.840 1377.500 419.040 ;
  RECT 1374.360 415.860 1375.220 416.140 ;
  RECT 1374.080 416.640 1377.500 417.840 ;
  RECT 1374.080 414.160 1377.500 415.360 ;
  RECT 1374.360 412.180 1375.220 412.460 ;
  RECT 1374.080 412.960 1377.500 414.160 ;
  RECT 1374.080 410.480 1377.500 411.680 ;
  RECT 1374.360 408.500 1375.220 408.780 ;
  RECT 1374.080 409.280 1377.500 410.480 ;
  RECT 1374.080 406.800 1377.500 408.000 ;
  RECT 1374.360 404.820 1375.220 405.100 ;
  RECT 1374.080 405.600 1377.500 406.800 ;
  RECT 1374.080 403.120 1377.500 404.320 ;
  RECT 1374.360 401.140 1375.220 401.420 ;
  RECT 1374.080 401.920 1377.500 403.120 ;
  RECT 1374.080 399.440 1377.500 400.640 ;
  RECT 1374.360 397.460 1375.220 397.740 ;
  RECT 1374.080 398.240 1377.500 399.440 ;
  RECT 1374.080 395.760 1377.500 396.960 ;
  RECT 1374.360 393.780 1375.220 394.060 ;
  RECT 1374.080 394.560 1377.500 395.760 ;
  RECT 1374.080 392.080 1377.500 393.280 ;
  RECT 1374.360 390.100 1375.220 390.380 ;
  RECT 1374.080 390.880 1377.500 392.080 ;
  RECT 1374.080 388.400 1377.500 389.600 ;
  RECT 1374.360 386.420 1375.220 386.700 ;
  RECT 1374.080 387.200 1377.500 388.400 ;
  RECT 1374.080 384.720 1377.500 385.920 ;
  RECT 1374.360 382.740 1375.220 383.020 ;
  RECT 1374.080 383.520 1377.500 384.720 ;
  RECT 1374.080 381.040 1377.500 382.240 ;
  RECT 1374.360 379.060 1375.220 379.340 ;
  RECT 1374.080 379.840 1377.500 381.040 ;
  RECT 1374.080 377.360 1377.500 378.560 ;
  RECT 1374.360 375.380 1375.220 375.660 ;
  RECT 1374.080 376.160 1377.500 377.360 ;
  RECT 1374.080 373.680 1377.500 374.880 ;
  RECT 1374.360 371.700 1375.220 371.980 ;
  RECT 1374.080 372.480 1377.500 373.680 ;
  RECT 1374.080 370.000 1377.500 371.200 ;
  RECT 1374.360 368.020 1375.220 368.300 ;
  RECT 1374.080 368.800 1377.500 370.000 ;
  RECT 1374.080 366.320 1377.500 367.520 ;
  RECT 1374.360 364.340 1375.220 364.620 ;
  RECT 1374.080 365.120 1377.500 366.320 ;
  RECT 1374.080 362.640 1377.500 363.840 ;
  RECT 1374.360 360.660 1375.220 360.940 ;
  RECT 1374.080 361.440 1377.500 362.640 ;
  RECT 1374.080 358.960 1377.500 360.160 ;
  RECT 1374.360 356.980 1375.220 357.260 ;
  RECT 1374.080 357.760 1377.500 358.960 ;
  RECT 1374.080 355.280 1377.500 356.480 ;
  RECT 1374.360 353.300 1375.220 353.580 ;
  RECT 1374.080 354.080 1377.500 355.280 ;
  RECT 1374.080 351.600 1377.500 352.800 ;
  RECT 1374.360 349.620 1375.220 349.900 ;
  RECT 1374.080 350.400 1377.500 351.600 ;
  RECT 1374.080 347.920 1377.500 349.120 ;
  RECT 1374.360 345.940 1375.220 346.220 ;
  RECT 1374.080 346.720 1377.500 347.920 ;
  RECT 1374.080 344.240 1377.500 345.440 ;
  RECT 1374.360 342.260 1375.220 342.540 ;
  RECT 1374.080 343.040 1377.500 344.240 ;
  RECT 1374.080 340.560 1377.500 341.760 ;
  RECT 1374.360 338.580 1375.220 338.860 ;
  RECT 1374.080 339.360 1377.500 340.560 ;
  RECT 1374.080 336.880 1377.500 338.080 ;
  RECT 1374.360 334.900 1375.220 335.180 ;
  RECT 1374.080 335.680 1377.500 336.880 ;
  RECT 1374.080 333.200 1377.500 334.400 ;
  RECT 1374.360 331.220 1375.220 331.500 ;
  RECT 1374.080 332.000 1377.500 333.200 ;
  RECT 1374.080 329.520 1377.500 330.720 ;
  RECT 1374.360 327.540 1375.220 327.820 ;
  RECT 1374.080 328.320 1377.500 329.520 ;
  RECT 1374.080 325.840 1377.500 327.040 ;
  RECT 1374.360 323.860 1375.220 324.140 ;
  RECT 1374.080 324.640 1377.500 325.840 ;
  RECT 1374.080 322.160 1377.500 323.360 ;
  RECT 1374.360 320.180 1375.220 320.460 ;
  RECT 1374.080 320.960 1377.500 322.160 ;
  RECT 1374.080 318.480 1377.500 319.680 ;
  RECT 1374.360 316.500 1375.220 316.780 ;
  RECT 1374.080 317.280 1377.500 318.480 ;
  RECT 1374.080 314.800 1377.500 316.000 ;
  RECT 1374.360 312.820 1375.220 313.100 ;
  RECT 1374.080 313.600 1377.500 314.800 ;
  RECT 1374.080 311.120 1377.500 312.320 ;
  RECT 1374.360 309.140 1375.220 309.420 ;
  RECT 1374.080 309.920 1377.500 311.120 ;
  RECT 1374.080 307.440 1377.500 308.640 ;
  RECT 1374.360 305.460 1375.220 305.740 ;
  RECT 1374.080 306.240 1377.500 307.440 ;
  RECT 1374.080 303.760 1377.500 304.960 ;
  RECT 1374.360 301.780 1375.220 302.060 ;
  RECT 1374.080 302.560 1377.500 303.760 ;
  RECT 1374.080 300.080 1377.500 301.280 ;
  RECT 1374.360 298.100 1375.220 298.380 ;
  RECT 1374.080 298.880 1377.500 300.080 ;
  RECT 1374.080 296.400 1377.500 297.600 ;
  RECT 1374.360 294.420 1375.220 294.700 ;
  RECT 1374.080 295.200 1377.500 296.400 ;
  RECT 1374.080 292.720 1377.500 293.920 ;
  RECT 1374.360 290.740 1375.220 291.020 ;
  RECT 1374.080 291.520 1377.500 292.720 ;
  RECT 1374.080 289.040 1377.500 290.240 ;
  RECT 1374.360 287.060 1375.220 287.340 ;
  RECT 1374.080 287.840 1377.500 289.040 ;
  RECT 1374.080 285.360 1377.500 286.560 ;
  RECT 1374.360 283.380 1375.220 283.660 ;
  RECT 1374.080 284.160 1377.500 285.360 ;
  RECT 1374.080 281.680 1377.500 282.880 ;
  RECT 1374.360 279.700 1375.220 279.980 ;
  RECT 1374.080 280.480 1377.500 281.680 ;
  RECT 1374.080 278.000 1377.500 279.200 ;
  RECT 1374.360 276.020 1375.220 276.300 ;
  RECT 1374.080 276.800 1377.500 278.000 ;
  RECT 1374.080 274.320 1377.500 275.520 ;
  RECT 1374.360 272.340 1375.220 272.620 ;
  RECT 1374.080 273.120 1377.500 274.320 ;
  RECT 1374.080 270.640 1377.500 271.840 ;
  RECT 1374.360 268.660 1375.220 268.940 ;
  RECT 1374.080 269.440 1377.500 270.640 ;
  RECT 1374.080 266.960 1377.500 268.160 ;
  RECT 1374.360 264.980 1375.220 265.260 ;
  RECT 1374.080 265.760 1377.500 266.960 ;
  RECT 1374.080 263.280 1377.500 264.480 ;
  RECT 1374.360 261.300 1375.220 261.580 ;
  RECT 1374.080 262.080 1377.500 263.280 ;
  RECT 1374.080 259.600 1377.500 260.800 ;
  RECT 1374.360 257.620 1375.220 257.900 ;
  RECT 1374.080 258.400 1377.500 259.600 ;
  RECT 1374.080 255.920 1377.500 257.120 ;
  RECT 1374.360 253.940 1375.220 254.220 ;
  RECT 1374.080 254.720 1377.500 255.920 ;
  RECT 1374.080 252.240 1377.500 253.440 ;
  RECT 1374.360 250.260 1375.220 250.540 ;
  RECT 1374.080 251.040 1377.500 252.240 ;
  RECT 1374.080 248.560 1377.500 249.760 ;
  RECT 1374.360 246.580 1375.220 246.860 ;
  RECT 1374.080 247.360 1377.500 248.560 ;
  RECT 1374.080 244.880 1377.500 246.080 ;
  RECT 1374.360 242.900 1375.220 243.180 ;
  RECT 1374.080 243.680 1377.500 244.880 ;
  RECT 1374.080 241.200 1377.500 242.400 ;
  RECT 1374.360 239.220 1375.220 239.500 ;
  RECT 1374.080 240.000 1377.500 241.200 ;
  RECT 1374.080 237.520 1377.500 238.720 ;
  RECT 1374.360 235.540 1375.220 235.820 ;
  RECT 1374.080 236.320 1377.500 237.520 ;
  RECT 1374.080 233.840 1377.500 235.040 ;
  RECT 1374.360 231.860 1375.220 232.140 ;
  RECT 1374.080 232.640 1377.500 233.840 ;
  RECT 1374.080 230.160 1377.500 231.360 ;
  RECT 1374.360 228.180 1375.220 228.460 ;
  RECT 1374.080 228.960 1377.500 230.160 ;
  RECT 1374.080 226.480 1377.500 227.680 ;
  RECT 1374.360 224.500 1375.220 224.780 ;
  RECT 1374.080 225.280 1377.500 226.480 ;
  RECT 1374.080 222.800 1377.500 224.000 ;
  RECT 1374.360 220.820 1375.220 221.100 ;
  RECT 1374.080 221.600 1377.500 222.800 ;
  RECT 1374.080 219.120 1377.500 220.320 ;
  RECT 1374.360 217.140 1375.220 217.420 ;
  RECT 1374.080 217.920 1377.500 219.120 ;
  RECT 1374.080 215.440 1377.500 216.640 ;
  RECT 1374.360 213.460 1375.220 213.740 ;
  RECT 1374.080 214.240 1377.500 215.440 ;
  RECT 1374.080 211.760 1377.500 212.960 ;
  RECT 1374.360 209.780 1375.220 210.060 ;
  RECT 1374.080 210.560 1377.500 211.760 ;
  RECT 1374.080 208.080 1377.500 209.280 ;
  RECT 1374.360 206.100 1375.220 206.380 ;
  RECT 1374.080 206.880 1377.500 208.080 ;
  RECT 1374.080 204.400 1377.500 205.600 ;
  RECT 1374.360 202.420 1375.220 202.700 ;
  RECT 1374.080 203.200 1377.500 204.400 ;
  RECT 1374.080 200.720 1377.500 201.920 ;
  RECT 1374.360 198.740 1375.220 199.020 ;
  RECT 1374.080 199.520 1377.500 200.720 ;
  RECT 1374.080 197.040 1377.500 198.240 ;
  RECT 1374.360 195.060 1375.220 195.340 ;
  RECT 1374.080 195.840 1377.500 197.040 ;
  RECT 1374.080 193.360 1377.500 194.560 ;
  RECT 1374.360 191.380 1375.220 191.660 ;
  RECT 1374.080 192.160 1377.500 193.360 ;
  RECT 1374.080 189.680 1377.500 190.880 ;
  RECT 1374.360 187.700 1375.220 187.980 ;
  RECT 1374.080 188.480 1377.500 189.680 ;
  RECT 1374.080 186.000 1377.500 187.200 ;
  RECT 1374.360 184.020 1375.220 184.300 ;
  RECT 1374.080 184.800 1377.500 186.000 ;
  RECT 1374.080 182.320 1377.500 183.520 ;
  RECT 1374.360 180.340 1375.220 180.620 ;
  RECT 1374.080 181.120 1377.500 182.320 ;
  RECT 1374.080 178.640 1377.500 179.840 ;
  RECT 1374.360 176.660 1375.220 176.940 ;
  RECT 1374.080 177.440 1377.500 178.640 ;
  RECT 1374.080 174.960 1377.500 176.160 ;
  RECT 1374.360 172.980 1375.220 173.260 ;
  RECT 1374.080 173.760 1377.500 174.960 ;
  RECT 1374.080 171.280 1377.500 172.480 ;
  RECT 1374.360 169.300 1375.220 169.580 ;
  RECT 1374.080 170.080 1377.500 171.280 ;
  RECT 1374.080 167.600 1377.500 168.800 ;
  RECT 1374.360 165.620 1375.220 165.900 ;
  RECT 1374.080 166.400 1377.500 167.600 ;
  RECT 1374.080 163.920 1377.500 165.120 ;
  RECT 1374.360 161.940 1375.220 162.220 ;
  RECT 1374.080 162.720 1377.500 163.920 ;
  RECT 1374.080 160.240 1377.500 161.440 ;
  RECT 1374.360 158.260 1375.220 158.540 ;
  RECT 1374.080 159.040 1377.500 160.240 ;
  RECT 1374.080 156.560 1377.500 157.760 ;
  RECT 1374.360 154.580 1375.220 154.860 ;
  RECT 1374.080 155.360 1377.500 156.560 ;
  RECT 1374.080 152.880 1377.500 154.080 ;
  RECT 1374.360 150.900 1375.220 151.180 ;
  RECT 1374.080 151.680 1377.500 152.880 ;
  RECT 1374.080 149.200 1377.500 150.400 ;
  RECT 1374.360 147.220 1375.220 147.500 ;
  RECT 1374.080 148.000 1377.500 149.200 ;
  RECT 1374.080 145.520 1377.500 146.720 ;
  RECT 1374.360 143.540 1375.220 143.820 ;
  RECT 1374.080 144.320 1377.500 145.520 ;
  RECT 1374.080 141.840 1377.500 143.040 ;
  RECT 1374.360 139.860 1375.220 140.140 ;
  RECT 1374.080 140.640 1377.500 141.840 ;
  RECT 1374.080 138.160 1377.500 139.360 ;
  RECT 1374.360 136.180 1375.220 136.460 ;
  RECT 1374.080 136.960 1377.500 138.160 ;
  RECT 1374.080 134.480 1377.500 135.680 ;
  RECT 1374.360 132.500 1375.220 132.780 ;
  RECT 1374.080 133.280 1377.500 134.480 ;
  RECT 1374.080 130.800 1377.500 132.000 ;
  RECT 1374.360 128.820 1375.220 129.100 ;
  RECT 1374.080 129.600 1377.500 130.800 ;
  RECT 1374.080 127.120 1377.500 128.320 ;
  RECT 1374.360 125.140 1375.220 125.420 ;
  RECT 1374.080 125.920 1377.500 127.120 ;
  RECT 1374.080 123.440 1377.500 124.640 ;
  RECT 1374.360 121.460 1375.220 121.740 ;
  RECT 1374.080 122.240 1377.500 123.440 ;
  RECT 1374.080 119.760 1377.500 120.960 ;
  RECT 1374.360 117.780 1375.220 118.060 ;
  RECT 1374.080 118.560 1377.500 119.760 ;
  RECT 1374.080 116.080 1377.500 117.280 ;
  RECT 1374.360 114.100 1375.220 114.380 ;
  RECT 1374.080 114.880 1377.500 116.080 ;
  RECT 1374.080 112.400 1377.500 113.600 ;
  RECT 1374.360 110.420 1375.220 110.700 ;
  RECT 1374.080 111.200 1377.500 112.400 ;
  RECT 1374.080 108.720 1377.500 109.920 ;
  RECT 1374.360 106.740 1375.220 107.020 ;
  RECT 1374.080 107.520 1377.500 108.720 ;
  RECT 1374.080 105.040 1377.500 106.240 ;
  RECT 1374.360 103.060 1375.220 103.340 ;
  RECT 1374.080 103.840 1377.500 105.040 ;
  RECT 1374.080 101.360 1377.500 102.560 ;
  RECT 1374.360 99.380 1375.220 99.660 ;
  RECT 1374.080 100.160 1377.500 101.360 ;
  RECT 1374.080 97.680 1377.500 98.880 ;
  RECT 1374.360 95.700 1375.220 95.980 ;
  RECT 1374.080 96.480 1377.500 97.680 ;
  RECT 1374.080 94.000 1377.500 95.200 ;
  RECT 1374.360 92.020 1375.220 92.300 ;
  RECT 1374.080 92.800 1377.500 94.000 ;
  RECT 1374.080 90.320 1377.500 91.520 ;
  RECT 1374.360 88.340 1375.220 88.620 ;
  RECT 1374.080 89.120 1377.500 90.320 ;
  RECT 1374.080 86.640 1377.500 87.840 ;
  RECT 1374.360 84.660 1375.220 84.940 ;
  RECT 1374.080 85.440 1377.500 86.640 ;
  RECT 1374.080 82.960 1377.500 84.160 ;
  RECT 1374.360 80.980 1375.220 81.260 ;
  RECT 1374.080 81.760 1377.500 82.960 ;
  RECT 1374.080 79.280 1377.500 80.480 ;
  RECT 1374.360 77.300 1375.220 77.580 ;
  RECT 1374.080 78.080 1377.500 79.280 ;
  RECT 1374.080 75.600 1377.500 76.800 ;
  RECT 1374.360 73.620 1375.220 73.900 ;
  RECT 1374.080 74.400 1377.500 75.600 ;
  RECT 1374.080 71.920 1377.500 73.120 ;
  RECT 1374.360 69.940 1375.220 70.220 ;
  RECT 1374.080 70.720 1377.500 71.920 ;
  RECT 1374.080 68.240 1377.500 69.440 ;
  RECT 1374.360 65.600 1375.220 65.980 ;
  RECT 717.530 545.790 717.780 549.210 ;
  RECT 718.100 546.070 718.350 546.930 ;
  RECT 758.450 545.790 758.700 549.210 ;
  RECT 759.020 546.070 759.270 546.930 ;
  RECT 799.370 545.790 799.620 549.210 ;
  RECT 799.940 546.070 800.190 546.930 ;
  RECT 840.290 545.790 840.540 549.210 ;
  RECT 840.860 546.070 841.110 546.930 ;
  RECT 881.210 545.790 881.460 549.210 ;
  RECT 881.780 546.070 882.030 546.930 ;
  RECT 922.130 545.790 922.380 549.210 ;
  RECT 922.700 546.070 922.950 546.930 ;
  RECT 963.050 545.790 963.300 549.210 ;
  RECT 963.620 546.070 963.870 546.930 ;
  RECT 1003.970 545.790 1004.220 549.210 ;
  RECT 1004.540 546.070 1004.790 546.930 ;
  RECT 1044.890 545.790 1045.140 549.210 ;
  RECT 1045.460 546.070 1045.710 546.930 ;
  RECT 1085.810 545.790 1086.060 549.210 ;
  RECT 1086.380 546.070 1086.630 546.930 ;
  RECT 1126.730 545.790 1126.980 549.210 ;
  RECT 1127.300 546.070 1127.550 546.930 ;
  RECT 1167.650 545.790 1167.900 549.210 ;
  RECT 1168.220 546.070 1168.470 546.930 ;
  RECT 1208.570 545.790 1208.820 549.210 ;
  RECT 1209.140 546.070 1209.390 546.930 ;
  RECT 1249.490 545.790 1249.740 549.210 ;
  RECT 1250.060 546.070 1250.310 546.930 ;
  RECT 1290.410 545.790 1290.660 549.210 ;
  RECT 1290.980 546.070 1291.230 546.930 ;
  RECT 1331.330 545.790 1331.580 549.210 ;
  RECT 1331.900 546.070 1332.150 546.930 ;
  RECT 714.040 545.790 714.940 549.210 ;
  RECT 684.720 545.790 687.910 549.210 ;
  RECT 694.720 545.790 699.040 549.210 ;
  RECT 701.090 546.070 703.600 546.930 ;
  RECT 688.670 546.070 691.060 546.930 ;
  RECT 681.160 546.070 684.220 546.930 ;
  RECT 705.340 546.070 708.190 546.930 ;
  RECT 709.640 546.070 712.890 546.930 ;
  RECT 676.440 545.790 678.200 549.210 ;
  RECT 678.440 546.070 680.200 546.930 ;
  RECT 671.100 545.790 672.860 549.210 ;
  RECT 667.100 545.790 668.860 549.210 ;
  RECT 663.180 545.790 664.860 549.210 ;
  RECT 673.100 546.070 674.860 546.930 ;
  RECT 669.100 546.070 670.860 546.930 ;
  RECT 665.100 546.070 666.860 546.930 ;
  RECT 662.080 545.790 662.980 549.210 ;
  RECT 4.280 65.600 5.140 65.980 ;
  RECT 2.000 68.240 5.420 69.440 ;
  RECT 2.000 70.720 5.420 71.920 ;
  RECT 4.280 69.940 5.140 70.220 ;
  RECT 2.000 71.920 5.420 73.120 ;
  RECT 2.000 74.400 5.420 75.600 ;
  RECT 4.280 73.620 5.140 73.900 ;
  RECT 2.000 75.600 5.420 76.800 ;
  RECT 2.000 78.080 5.420 79.280 ;
  RECT 4.280 77.300 5.140 77.580 ;
  RECT 2.000 79.280 5.420 80.480 ;
  RECT 2.000 81.760 5.420 82.960 ;
  RECT 4.280 80.980 5.140 81.260 ;
  RECT 2.000 82.960 5.420 84.160 ;
  RECT 2.000 85.440 5.420 86.640 ;
  RECT 4.280 84.660 5.140 84.940 ;
  RECT 2.000 86.640 5.420 87.840 ;
  RECT 2.000 89.120 5.420 90.320 ;
  RECT 4.280 88.340 5.140 88.620 ;
  RECT 2.000 90.320 5.420 91.520 ;
  RECT 2.000 92.800 5.420 94.000 ;
  RECT 4.280 92.020 5.140 92.300 ;
  RECT 2.000 94.000 5.420 95.200 ;
  RECT 2.000 96.480 5.420 97.680 ;
  RECT 4.280 95.700 5.140 95.980 ;
  RECT 2.000 97.680 5.420 98.880 ;
  RECT 2.000 100.160 5.420 101.360 ;
  RECT 4.280 99.380 5.140 99.660 ;
  RECT 2.000 101.360 5.420 102.560 ;
  RECT 2.000 103.840 5.420 105.040 ;
  RECT 4.280 103.060 5.140 103.340 ;
  RECT 2.000 105.040 5.420 106.240 ;
  RECT 2.000 107.520 5.420 108.720 ;
  RECT 4.280 106.740 5.140 107.020 ;
  RECT 2.000 108.720 5.420 109.920 ;
  RECT 2.000 111.200 5.420 112.400 ;
  RECT 4.280 110.420 5.140 110.700 ;
  RECT 2.000 112.400 5.420 113.600 ;
  RECT 2.000 114.880 5.420 116.080 ;
  RECT 4.280 114.100 5.140 114.380 ;
  RECT 2.000 116.080 5.420 117.280 ;
  RECT 2.000 118.560 5.420 119.760 ;
  RECT 4.280 117.780 5.140 118.060 ;
  RECT 2.000 119.760 5.420 120.960 ;
  RECT 2.000 122.240 5.420 123.440 ;
  RECT 4.280 121.460 5.140 121.740 ;
  RECT 2.000 123.440 5.420 124.640 ;
  RECT 2.000 125.920 5.420 127.120 ;
  RECT 4.280 125.140 5.140 125.420 ;
  RECT 2.000 127.120 5.420 128.320 ;
  RECT 2.000 129.600 5.420 130.800 ;
  RECT 4.280 128.820 5.140 129.100 ;
  RECT 2.000 130.800 5.420 132.000 ;
  RECT 2.000 133.280 5.420 134.480 ;
  RECT 4.280 132.500 5.140 132.780 ;
  RECT 2.000 134.480 5.420 135.680 ;
  RECT 2.000 136.960 5.420 138.160 ;
  RECT 4.280 136.180 5.140 136.460 ;
  RECT 2.000 138.160 5.420 139.360 ;
  RECT 2.000 140.640 5.420 141.840 ;
  RECT 4.280 139.860 5.140 140.140 ;
  RECT 2.000 141.840 5.420 143.040 ;
  RECT 2.000 144.320 5.420 145.520 ;
  RECT 4.280 143.540 5.140 143.820 ;
  RECT 2.000 145.520 5.420 146.720 ;
  RECT 2.000 148.000 5.420 149.200 ;
  RECT 4.280 147.220 5.140 147.500 ;
  RECT 2.000 149.200 5.420 150.400 ;
  RECT 2.000 151.680 5.420 152.880 ;
  RECT 4.280 150.900 5.140 151.180 ;
  RECT 2.000 152.880 5.420 154.080 ;
  RECT 2.000 155.360 5.420 156.560 ;
  RECT 4.280 154.580 5.140 154.860 ;
  RECT 2.000 156.560 5.420 157.760 ;
  RECT 2.000 159.040 5.420 160.240 ;
  RECT 4.280 158.260 5.140 158.540 ;
  RECT 2.000 160.240 5.420 161.440 ;
  RECT 2.000 162.720 5.420 163.920 ;
  RECT 4.280 161.940 5.140 162.220 ;
  RECT 2.000 163.920 5.420 165.120 ;
  RECT 2.000 166.400 5.420 167.600 ;
  RECT 4.280 165.620 5.140 165.900 ;
  RECT 2.000 167.600 5.420 168.800 ;
  RECT 2.000 170.080 5.420 171.280 ;
  RECT 4.280 169.300 5.140 169.580 ;
  RECT 2.000 171.280 5.420 172.480 ;
  RECT 2.000 173.760 5.420 174.960 ;
  RECT 4.280 172.980 5.140 173.260 ;
  RECT 2.000 174.960 5.420 176.160 ;
  RECT 2.000 177.440 5.420 178.640 ;
  RECT 4.280 176.660 5.140 176.940 ;
  RECT 2.000 178.640 5.420 179.840 ;
  RECT 2.000 181.120 5.420 182.320 ;
  RECT 4.280 180.340 5.140 180.620 ;
  RECT 2.000 182.320 5.420 183.520 ;
  RECT 2.000 184.800 5.420 186.000 ;
  RECT 4.280 184.020 5.140 184.300 ;
  RECT 2.000 186.000 5.420 187.200 ;
  RECT 2.000 188.480 5.420 189.680 ;
  RECT 4.280 187.700 5.140 187.980 ;
  RECT 2.000 189.680 5.420 190.880 ;
  RECT 2.000 192.160 5.420 193.360 ;
  RECT 4.280 191.380 5.140 191.660 ;
  RECT 2.000 193.360 5.420 194.560 ;
  RECT 2.000 195.840 5.420 197.040 ;
  RECT 4.280 195.060 5.140 195.340 ;
  RECT 2.000 197.040 5.420 198.240 ;
  RECT 2.000 199.520 5.420 200.720 ;
  RECT 4.280 198.740 5.140 199.020 ;
  RECT 2.000 200.720 5.420 201.920 ;
  RECT 2.000 203.200 5.420 204.400 ;
  RECT 4.280 202.420 5.140 202.700 ;
  RECT 2.000 204.400 5.420 205.600 ;
  RECT 2.000 206.880 5.420 208.080 ;
  RECT 4.280 206.100 5.140 206.380 ;
  RECT 2.000 208.080 5.420 209.280 ;
  RECT 2.000 210.560 5.420 211.760 ;
  RECT 4.280 209.780 5.140 210.060 ;
  RECT 2.000 211.760 5.420 212.960 ;
  RECT 2.000 214.240 5.420 215.440 ;
  RECT 4.280 213.460 5.140 213.740 ;
  RECT 2.000 215.440 5.420 216.640 ;
  RECT 2.000 217.920 5.420 219.120 ;
  RECT 4.280 217.140 5.140 217.420 ;
  RECT 2.000 219.120 5.420 220.320 ;
  RECT 2.000 221.600 5.420 222.800 ;
  RECT 4.280 220.820 5.140 221.100 ;
  RECT 2.000 222.800 5.420 224.000 ;
  RECT 2.000 225.280 5.420 226.480 ;
  RECT 4.280 224.500 5.140 224.780 ;
  RECT 2.000 226.480 5.420 227.680 ;
  RECT 2.000 228.960 5.420 230.160 ;
  RECT 4.280 228.180 5.140 228.460 ;
  RECT 2.000 230.160 5.420 231.360 ;
  RECT 2.000 232.640 5.420 233.840 ;
  RECT 4.280 231.860 5.140 232.140 ;
  RECT 2.000 233.840 5.420 235.040 ;
  RECT 2.000 236.320 5.420 237.520 ;
  RECT 4.280 235.540 5.140 235.820 ;
  RECT 2.000 237.520 5.420 238.720 ;
  RECT 2.000 240.000 5.420 241.200 ;
  RECT 4.280 239.220 5.140 239.500 ;
  RECT 2.000 241.200 5.420 242.400 ;
  RECT 2.000 243.680 5.420 244.880 ;
  RECT 4.280 242.900 5.140 243.180 ;
  RECT 2.000 244.880 5.420 246.080 ;
  RECT 2.000 247.360 5.420 248.560 ;
  RECT 4.280 246.580 5.140 246.860 ;
  RECT 2.000 248.560 5.420 249.760 ;
  RECT 2.000 251.040 5.420 252.240 ;
  RECT 4.280 250.260 5.140 250.540 ;
  RECT 2.000 252.240 5.420 253.440 ;
  RECT 2.000 254.720 5.420 255.920 ;
  RECT 4.280 253.940 5.140 254.220 ;
  RECT 2.000 255.920 5.420 257.120 ;
  RECT 2.000 258.400 5.420 259.600 ;
  RECT 4.280 257.620 5.140 257.900 ;
  RECT 2.000 259.600 5.420 260.800 ;
  RECT 2.000 262.080 5.420 263.280 ;
  RECT 4.280 261.300 5.140 261.580 ;
  RECT 2.000 263.280 5.420 264.480 ;
  RECT 2.000 265.760 5.420 266.960 ;
  RECT 4.280 264.980 5.140 265.260 ;
  RECT 2.000 266.960 5.420 268.160 ;
  RECT 2.000 269.440 5.420 270.640 ;
  RECT 4.280 268.660 5.140 268.940 ;
  RECT 2.000 270.640 5.420 271.840 ;
  RECT 2.000 273.120 5.420 274.320 ;
  RECT 4.280 272.340 5.140 272.620 ;
  RECT 2.000 274.320 5.420 275.520 ;
  RECT 2.000 276.800 5.420 278.000 ;
  RECT 4.280 276.020 5.140 276.300 ;
  RECT 2.000 278.000 5.420 279.200 ;
  RECT 2.000 280.480 5.420 281.680 ;
  RECT 4.280 279.700 5.140 279.980 ;
  RECT 2.000 281.680 5.420 282.880 ;
  RECT 2.000 284.160 5.420 285.360 ;
  RECT 4.280 283.380 5.140 283.660 ;
  RECT 2.000 285.360 5.420 286.560 ;
  RECT 2.000 287.840 5.420 289.040 ;
  RECT 4.280 287.060 5.140 287.340 ;
  RECT 2.000 289.040 5.420 290.240 ;
  RECT 2.000 291.520 5.420 292.720 ;
  RECT 4.280 290.740 5.140 291.020 ;
  RECT 2.000 292.720 5.420 293.920 ;
  RECT 2.000 295.200 5.420 296.400 ;
  RECT 4.280 294.420 5.140 294.700 ;
  RECT 2.000 296.400 5.420 297.600 ;
  RECT 2.000 298.880 5.420 300.080 ;
  RECT 4.280 298.100 5.140 298.380 ;
  RECT 2.000 300.080 5.420 301.280 ;
  RECT 2.000 302.560 5.420 303.760 ;
  RECT 4.280 301.780 5.140 302.060 ;
  RECT 2.000 303.760 5.420 304.960 ;
  RECT 2.000 306.240 5.420 307.440 ;
  RECT 4.280 305.460 5.140 305.740 ;
  RECT 2.000 307.440 5.420 308.640 ;
  RECT 2.000 309.920 5.420 311.120 ;
  RECT 4.280 309.140 5.140 309.420 ;
  RECT 2.000 311.120 5.420 312.320 ;
  RECT 2.000 313.600 5.420 314.800 ;
  RECT 4.280 312.820 5.140 313.100 ;
  RECT 2.000 314.800 5.420 316.000 ;
  RECT 2.000 317.280 5.420 318.480 ;
  RECT 4.280 316.500 5.140 316.780 ;
  RECT 2.000 318.480 5.420 319.680 ;
  RECT 2.000 320.960 5.420 322.160 ;
  RECT 4.280 320.180 5.140 320.460 ;
  RECT 2.000 322.160 5.420 323.360 ;
  RECT 2.000 324.640 5.420 325.840 ;
  RECT 4.280 323.860 5.140 324.140 ;
  RECT 2.000 325.840 5.420 327.040 ;
  RECT 2.000 328.320 5.420 329.520 ;
  RECT 4.280 327.540 5.140 327.820 ;
  RECT 2.000 329.520 5.420 330.720 ;
  RECT 2.000 332.000 5.420 333.200 ;
  RECT 4.280 331.220 5.140 331.500 ;
  RECT 2.000 333.200 5.420 334.400 ;
  RECT 2.000 335.680 5.420 336.880 ;
  RECT 4.280 334.900 5.140 335.180 ;
  RECT 2.000 336.880 5.420 338.080 ;
  RECT 2.000 339.360 5.420 340.560 ;
  RECT 4.280 338.580 5.140 338.860 ;
  RECT 2.000 340.560 5.420 341.760 ;
  RECT 2.000 343.040 5.420 344.240 ;
  RECT 4.280 342.260 5.140 342.540 ;
  RECT 2.000 344.240 5.420 345.440 ;
  RECT 2.000 346.720 5.420 347.920 ;
  RECT 4.280 345.940 5.140 346.220 ;
  RECT 2.000 347.920 5.420 349.120 ;
  RECT 2.000 350.400 5.420 351.600 ;
  RECT 4.280 349.620 5.140 349.900 ;
  RECT 2.000 351.600 5.420 352.800 ;
  RECT 2.000 354.080 5.420 355.280 ;
  RECT 4.280 353.300 5.140 353.580 ;
  RECT 2.000 355.280 5.420 356.480 ;
  RECT 2.000 357.760 5.420 358.960 ;
  RECT 4.280 356.980 5.140 357.260 ;
  RECT 2.000 358.960 5.420 360.160 ;
  RECT 2.000 361.440 5.420 362.640 ;
  RECT 4.280 360.660 5.140 360.940 ;
  RECT 2.000 362.640 5.420 363.840 ;
  RECT 2.000 365.120 5.420 366.320 ;
  RECT 4.280 364.340 5.140 364.620 ;
  RECT 2.000 366.320 5.420 367.520 ;
  RECT 2.000 368.800 5.420 370.000 ;
  RECT 4.280 368.020 5.140 368.300 ;
  RECT 2.000 370.000 5.420 371.200 ;
  RECT 2.000 372.480 5.420 373.680 ;
  RECT 4.280 371.700 5.140 371.980 ;
  RECT 2.000 373.680 5.420 374.880 ;
  RECT 2.000 376.160 5.420 377.360 ;
  RECT 4.280 375.380 5.140 375.660 ;
  RECT 2.000 377.360 5.420 378.560 ;
  RECT 2.000 379.840 5.420 381.040 ;
  RECT 4.280 379.060 5.140 379.340 ;
  RECT 2.000 381.040 5.420 382.240 ;
  RECT 2.000 383.520 5.420 384.720 ;
  RECT 4.280 382.740 5.140 383.020 ;
  RECT 2.000 384.720 5.420 385.920 ;
  RECT 2.000 387.200 5.420 388.400 ;
  RECT 4.280 386.420 5.140 386.700 ;
  RECT 2.000 388.400 5.420 389.600 ;
  RECT 2.000 390.880 5.420 392.080 ;
  RECT 4.280 390.100 5.140 390.380 ;
  RECT 2.000 392.080 5.420 393.280 ;
  RECT 2.000 394.560 5.420 395.760 ;
  RECT 4.280 393.780 5.140 394.060 ;
  RECT 2.000 395.760 5.420 396.960 ;
  RECT 2.000 398.240 5.420 399.440 ;
  RECT 4.280 397.460 5.140 397.740 ;
  RECT 2.000 399.440 5.420 400.640 ;
  RECT 2.000 401.920 5.420 403.120 ;
  RECT 4.280 401.140 5.140 401.420 ;
  RECT 2.000 403.120 5.420 404.320 ;
  RECT 2.000 405.600 5.420 406.800 ;
  RECT 4.280 404.820 5.140 405.100 ;
  RECT 2.000 406.800 5.420 408.000 ;
  RECT 2.000 409.280 5.420 410.480 ;
  RECT 4.280 408.500 5.140 408.780 ;
  RECT 2.000 410.480 5.420 411.680 ;
  RECT 2.000 412.960 5.420 414.160 ;
  RECT 4.280 412.180 5.140 412.460 ;
  RECT 2.000 414.160 5.420 415.360 ;
  RECT 2.000 416.640 5.420 417.840 ;
  RECT 4.280 415.860 5.140 416.140 ;
  RECT 2.000 417.840 5.420 419.040 ;
  RECT 2.000 420.320 5.420 421.520 ;
  RECT 4.280 419.540 5.140 419.820 ;
  RECT 2.000 421.520 5.420 422.720 ;
  RECT 2.000 424.000 5.420 425.200 ;
  RECT 4.280 423.220 5.140 423.500 ;
  RECT 2.000 425.200 5.420 426.400 ;
  RECT 2.000 427.680 5.420 428.880 ;
  RECT 4.280 426.900 5.140 427.180 ;
  RECT 2.000 428.880 5.420 430.080 ;
  RECT 2.000 431.360 5.420 432.560 ;
  RECT 4.280 430.580 5.140 430.860 ;
  RECT 2.000 432.560 5.420 433.760 ;
  RECT 2.000 435.040 5.420 436.240 ;
  RECT 4.280 434.260 5.140 434.540 ;
  RECT 2.000 436.240 5.420 437.440 ;
  RECT 2.000 438.720 5.420 439.920 ;
  RECT 4.280 437.940 5.140 438.220 ;
  RECT 2.000 439.920 5.420 441.120 ;
  RECT 2.000 442.400 5.420 443.600 ;
  RECT 4.280 441.620 5.140 441.900 ;
  RECT 2.000 443.600 5.420 444.800 ;
  RECT 2.000 446.080 5.420 447.280 ;
  RECT 4.280 445.300 5.140 445.580 ;
  RECT 2.000 447.280 5.420 448.480 ;
  RECT 2.000 449.760 5.420 450.960 ;
  RECT 4.280 448.980 5.140 449.260 ;
  RECT 2.000 450.960 5.420 452.160 ;
  RECT 2.000 453.440 5.420 454.640 ;
  RECT 4.280 452.660 5.140 452.940 ;
  RECT 2.000 454.640 5.420 455.840 ;
  RECT 2.000 457.120 5.420 458.320 ;
  RECT 4.280 456.340 5.140 456.620 ;
  RECT 2.000 458.320 5.420 459.520 ;
  RECT 2.000 460.800 5.420 462.000 ;
  RECT 4.280 460.020 5.140 460.300 ;
  RECT 2.000 462.000 5.420 463.200 ;
  RECT 2.000 464.480 5.420 465.680 ;
  RECT 4.280 463.700 5.140 463.980 ;
  RECT 2.000 465.680 5.420 466.880 ;
  RECT 2.000 468.160 5.420 469.360 ;
  RECT 4.280 467.380 5.140 467.660 ;
  RECT 2.000 469.360 5.420 470.560 ;
  RECT 2.000 471.840 5.420 473.040 ;
  RECT 4.280 471.060 5.140 471.340 ;
  RECT 2.000 473.040 5.420 474.240 ;
  RECT 2.000 475.520 5.420 476.720 ;
  RECT 4.280 474.740 5.140 475.020 ;
  RECT 2.000 476.720 5.420 477.920 ;
  RECT 2.000 479.200 5.420 480.400 ;
  RECT 4.280 478.420 5.140 478.700 ;
  RECT 2.000 480.400 5.420 481.600 ;
  RECT 2.000 482.880 5.420 484.080 ;
  RECT 4.280 482.100 5.140 482.380 ;
  RECT 2.000 484.080 5.420 485.280 ;
  RECT 2.000 486.560 5.420 487.760 ;
  RECT 4.280 485.780 5.140 486.060 ;
  RECT 2.000 487.760 5.420 488.960 ;
  RECT 2.000 490.240 5.420 491.440 ;
  RECT 4.280 489.460 5.140 489.740 ;
  RECT 2.000 491.440 5.420 492.640 ;
  RECT 2.000 493.920 5.420 495.120 ;
  RECT 4.280 493.140 5.140 493.420 ;
  RECT 2.000 495.120 5.420 496.320 ;
  RECT 2.000 497.600 5.420 498.800 ;
  RECT 4.280 496.820 5.140 497.100 ;
  RECT 2.000 498.800 5.420 500.000 ;
  RECT 2.000 501.280 5.420 502.480 ;
  RECT 4.280 500.500 5.140 500.780 ;
  RECT 2.000 502.480 5.420 503.680 ;
  RECT 2.000 504.960 5.420 506.160 ;
  RECT 4.280 504.180 5.140 504.460 ;
  RECT 2.000 506.160 5.420 507.360 ;
  RECT 2.000 508.640 5.420 509.840 ;
  RECT 4.280 507.860 5.140 508.140 ;
  RECT 2.000 509.840 5.420 511.040 ;
  RECT 2.000 512.320 5.420 513.520 ;
  RECT 4.280 511.540 5.140 511.820 ;
  RECT 2.000 513.520 5.420 514.720 ;
  RECT 2.000 516.000 5.420 517.200 ;
  RECT 4.280 515.220 5.140 515.500 ;
  RECT 2.000 517.200 5.420 518.400 ;
  RECT 2.000 519.680 5.420 520.880 ;
  RECT 4.280 518.900 5.140 519.180 ;
  RECT 2.000 520.880 5.420 522.080 ;
  RECT 2.000 523.360 5.420 524.560 ;
  RECT 4.280 522.580 5.140 522.860 ;
  RECT 2.000 524.560 5.420 525.760 ;
  RECT 2.000 527.040 5.420 528.240 ;
  RECT 4.280 526.260 5.140 526.540 ;
  RECT 2.000 528.240 5.420 529.440 ;
  RECT 2.000 530.720 5.420 531.920 ;
  RECT 4.280 529.940 5.140 530.220 ;
  RECT 2.000 531.920 5.420 533.120 ;
  RECT 2.000 534.400 5.420 535.600 ;
  RECT 4.280 533.620 5.140 533.900 ;
  RECT 2.000 535.600 5.420 536.800 ;
  RECT 2.000 538.080 5.420 539.280 ;
  RECT 4.280 537.300 5.140 537.580 ;
  RECT 4.280 545.220 5.140 545.600 ;
  RECT 47.920 545.790 48.170 549.210 ;
  RECT 47.350 546.070 47.600 546.930 ;
  RECT 88.840 545.790 89.090 549.210 ;
  RECT 88.270 546.070 88.520 546.930 ;
  RECT 129.760 545.790 130.010 549.210 ;
  RECT 129.190 546.070 129.440 546.930 ;
  RECT 170.680 545.790 170.930 549.210 ;
  RECT 170.110 546.070 170.360 546.930 ;
  RECT 211.600 545.790 211.850 549.210 ;
  RECT 211.030 546.070 211.280 546.930 ;
  RECT 252.520 545.790 252.770 549.210 ;
  RECT 251.950 546.070 252.200 546.930 ;
  RECT 293.440 545.790 293.690 549.210 ;
  RECT 292.870 546.070 293.120 546.930 ;
  RECT 334.360 545.790 334.610 549.210 ;
  RECT 333.790 546.070 334.040 546.930 ;
  RECT 375.280 545.790 375.530 549.210 ;
  RECT 374.710 546.070 374.960 546.930 ;
  RECT 416.200 545.790 416.450 549.210 ;
  RECT 415.630 546.070 415.880 546.930 ;
  RECT 457.120 545.790 457.370 549.210 ;
  RECT 456.550 546.070 456.800 546.930 ;
  RECT 498.040 545.790 498.290 549.210 ;
  RECT 497.470 546.070 497.720 546.930 ;
  RECT 538.960 545.790 539.210 549.210 ;
  RECT 538.390 546.070 538.640 546.930 ;
  RECT 579.880 545.790 580.130 549.210 ;
  RECT 579.310 546.070 579.560 546.930 ;
  RECT 620.800 545.790 621.050 549.210 ;
  RECT 620.230 546.070 620.480 546.930 ;
  RECT 0.000 549.210 1379.500 551.210 ;
  RECT 0.000 1.600 1379.500 3.600 ;
  RECT 1377.500 1.600 1379.500 551.210 ;
  RECT 0.000 1.600 2.000 551.210 ;
  LAYER ME2 ;
  RECT 5.420 7.020 1374.080 545.790 ;
  RECT 1377.640 3.460 1379.500 549.350 ;
  RECT 0.000 3.460 1.860 549.350 ;
  RECT 1.860 549.350 1377.640 551.210 ;
  RECT 1369.400 1.600 1377.640 3.460 ;
  RECT 1354.600 1.600 1366.840 3.460 ;
  RECT 1349.400 1.600 1352.210 3.460 ;
  RECT 1335.000 1.600 1347.000 3.460 ;
  RECT 1328.600 1.600 1332.370 3.460 ;
  RECT 1313.800 1.600 1325.920 3.460 ;
  RECT 1308.600 1.600 1311.290 3.460 ;
  RECT 1293.800 1.600 1306.080 3.460 ;
  RECT 1287.400 1.600 1291.450 3.460 ;
  RECT 1273.000 1.600 1285.000 3.460 ;
  RECT 1267.800 1.600 1270.370 3.460 ;
  RECT 1253.000 1.600 1265.160 3.460 ;
  RECT 1246.600 1.600 1250.530 3.460 ;
  RECT 1231.800 1.600 1244.080 3.460 ;
  RECT 1226.600 1.600 1229.450 3.460 ;
  RECT 1213.800 1.600 1224.240 3.460 ;
  RECT 1205.800 1.600 1209.610 3.460 ;
  RECT 1191.000 1.600 1203.160 3.460 ;
  RECT 1185.800 1.600 1188.530 3.460 ;
  RECT 1171.000 1.600 1183.320 3.460 ;
  RECT 1164.600 1.600 1168.690 3.460 ;
  RECT 1150.200 1.600 1162.240 3.460 ;
  RECT 1145.000 1.600 1147.610 3.460 ;
  RECT 1130.200 1.600 1142.400 3.460 ;
  RECT 1123.800 1.600 1127.770 3.460 ;
  RECT 1109.000 1.600 1121.320 3.460 ;
  RECT 1103.800 1.600 1106.690 3.460 ;
  RECT 1089.400 1.600 1101.480 3.460 ;
  RECT 1083.000 1.600 1086.850 3.460 ;
  RECT 1068.200 1.600 1080.400 3.460 ;
  RECT 1063.000 1.600 1065.770 3.460 ;
  RECT 1050.200 1.600 1060.560 3.460 ;
  RECT 1041.800 1.600 1045.930 3.460 ;
  RECT 1027.400 1.600 1039.480 3.460 ;
  RECT 1022.200 1.600 1024.850 3.460 ;
  RECT 1007.400 1.600 1019.640 3.460 ;
  RECT 1001.000 1.600 1005.010 3.460 ;
  RECT 986.600 1.600 998.560 3.460 ;
  RECT 981.400 1.600 983.930 3.460 ;
  RECT 966.600 1.600 978.720 3.460 ;
  RECT 960.200 1.600 964.090 3.460 ;
  RECT 945.400 1.600 957.640 3.460 ;
  RECT 940.200 1.600 943.010 3.460 ;
  RECT 925.800 1.600 937.800 3.460 ;
  RECT 919.400 1.600 923.170 3.460 ;
  RECT 904.600 1.600 916.720 3.460 ;
  RECT 899.400 1.600 902.090 3.460 ;
  RECT 886.600 1.600 896.880 3.460 ;
  RECT 878.200 1.600 882.250 3.460 ;
  RECT 863.800 1.600 875.800 3.460 ;
  RECT 858.600 1.600 861.170 3.460 ;
  RECT 843.800 1.600 855.960 3.460 ;
  RECT 837.400 1.600 841.330 3.460 ;
  RECT 822.600 1.600 834.880 3.460 ;
  RECT 817.400 1.600 820.250 3.460 ;
  RECT 803.000 1.600 815.040 3.460 ;
  RECT 796.600 1.600 800.410 3.460 ;
  RECT 781.800 1.600 793.960 3.460 ;
  RECT 776.600 1.600 779.330 3.460 ;
  RECT 761.800 1.600 774.120 3.460 ;
  RECT 755.400 1.600 759.490 3.460 ;
  RECT 741.000 1.600 753.040 3.460 ;
  RECT 735.800 1.600 738.410 3.460 ;
  RECT 722.600 1.600 733.200 3.460 ;
  RECT 700.200 1.600 718.570 3.460 ;
  RECT 688.200 1.600 691.730 3.460 ;
  RECT 681.000 1.600 685.760 3.460 ;
  RECT 658.200 1.600 662.640 3.460 ;
  RECT 643.800 1.600 655.740 3.460 ;
  RECT 638.200 1.600 641.110 3.460 ;
  RECT 623.800 1.600 635.900 3.460 ;
  RECT 617.400 1.600 621.270 3.460 ;
  RECT 602.600 1.600 614.820 3.460 ;
  RECT 597.400 1.600 600.190 3.460 ;
  RECT 583.000 1.600 594.980 3.460 ;
  RECT 576.200 1.600 580.350 3.460 ;
  RECT 561.800 1.600 573.900 3.460 ;
  RECT 556.600 1.600 559.270 3.460 ;
  RECT 541.800 1.600 554.060 3.460 ;
  RECT 535.400 1.600 539.430 3.460 ;
  RECT 521.000 1.600 532.980 3.460 ;
  RECT 515.800 1.600 518.350 3.460 ;
  RECT 502.600 1.600 513.140 3.460 ;
  RECT 494.600 1.600 498.510 3.460 ;
  RECT 479.800 1.600 492.060 3.460 ;
  RECT 474.600 1.600 477.430 3.460 ;
  RECT 460.200 1.600 472.220 3.460 ;
  RECT 453.800 1.600 457.590 3.460 ;
  RECT 439.000 1.600 451.140 3.460 ;
  RECT 433.800 1.600 436.510 3.460 ;
  RECT 419.000 1.600 431.300 3.460 ;
  RECT 412.600 1.600 416.670 3.460 ;
  RECT 398.200 1.600 410.220 3.460 ;
  RECT 393.000 1.600 395.590 3.460 ;
  RECT 378.200 1.600 390.380 3.460 ;
  RECT 371.800 1.600 375.750 3.460 ;
  RECT 357.000 1.600 369.300 3.460 ;
  RECT 351.800 1.600 354.670 3.460 ;
  RECT 339.000 1.600 349.460 3.460 ;
  RECT 331.000 1.600 334.830 3.460 ;
  RECT 316.200 1.600 328.380 3.460 ;
  RECT 311.000 1.600 313.750 3.460 ;
  RECT 296.600 1.600 308.540 3.460 ;
  RECT 289.800 1.600 293.910 3.460 ;
  RECT 275.400 1.600 287.460 3.460 ;
  RECT 270.200 1.600 272.830 3.460 ;
  RECT 255.400 1.600 267.620 3.460 ;
  RECT 249.000 1.600 252.990 3.460 ;
  RECT 234.600 1.600 246.540 3.460 ;
  RECT 229.000 1.600 231.910 3.460 ;
  RECT 214.600 1.600 226.700 3.460 ;
  RECT 208.200 1.600 212.070 3.460 ;
  RECT 193.400 1.600 205.620 3.460 ;
  RECT 188.200 1.600 190.990 3.460 ;
  RECT 175.400 1.600 185.780 3.460 ;
  RECT 167.000 1.600 171.150 3.460 ;
  RECT 152.600 1.600 164.700 3.460 ;
  RECT 147.400 1.600 150.070 3.460 ;
  RECT 132.600 1.600 144.860 3.460 ;
  RECT 126.200 1.600 130.230 3.460 ;
  RECT 111.800 1.600 123.780 3.460 ;
  RECT 106.600 1.600 109.150 3.460 ;
  RECT 91.800 1.600 103.940 3.460 ;
  RECT 85.400 1.600 89.310 3.460 ;
  RECT 70.600 1.600 82.860 3.460 ;
  RECT 65.400 1.600 68.230 3.460 ;
  RECT 51.000 1.600 63.020 3.460 ;
  RECT 44.600 1.600 48.390 3.460 ;
  RECT 29.800 1.600 41.940 3.460 ;
  RECT 24.600 1.600 27.310 3.460 ;
  RECT 11.800 1.600 22.100 3.460 ;
  RECT 1.860 1.600 7.470 3.460 ;
  RECT 1375.500 5.600 1377.360 547.210 ;
  RECT 2.140 5.600 4.000 547.210 ;
  RECT 4.000 547.210 1375.500 549.070 ;
  RECT 1369.400 3.740 1375.500 5.600 ;
  RECT 1354.600 3.740 1366.840 5.600 ;
  RECT 1349.400 3.740 1352.210 5.600 ;
  RECT 1335.000 3.740 1347.000 5.600 ;
  RECT 1328.600 3.740 1332.370 5.600 ;
  RECT 1313.800 3.740 1325.920 5.600 ;
  RECT 1308.600 3.740 1311.290 5.600 ;
  RECT 1293.800 3.740 1306.080 5.600 ;
  RECT 1287.400 3.740 1291.450 5.600 ;
  RECT 1273.000 3.740 1285.000 5.600 ;
  RECT 1267.800 3.740 1270.370 5.600 ;
  RECT 1253.000 3.740 1265.160 5.600 ;
  RECT 1246.600 3.740 1250.530 5.600 ;
  RECT 1231.800 3.740 1244.080 5.600 ;
  RECT 1226.600 3.740 1229.450 5.600 ;
  RECT 1213.800 3.740 1224.240 5.600 ;
  RECT 1205.800 3.740 1209.610 5.600 ;
  RECT 1191.000 3.740 1203.160 5.600 ;
  RECT 1185.800 3.740 1188.530 5.600 ;
  RECT 1171.000 3.740 1183.320 5.600 ;
  RECT 1164.600 3.740 1168.690 5.600 ;
  RECT 1150.200 3.740 1162.240 5.600 ;
  RECT 1145.000 3.740 1147.610 5.600 ;
  RECT 1130.200 3.740 1142.400 5.600 ;
  RECT 1123.800 3.740 1127.770 5.600 ;
  RECT 1109.000 3.740 1121.320 5.600 ;
  RECT 1103.800 3.740 1106.690 5.600 ;
  RECT 1089.400 3.740 1101.480 5.600 ;
  RECT 1083.000 3.740 1086.850 5.600 ;
  RECT 1068.200 3.740 1080.400 5.600 ;
  RECT 1063.000 3.740 1065.770 5.600 ;
  RECT 1050.200 3.740 1060.560 5.600 ;
  RECT 1041.800 3.740 1045.930 5.600 ;
  RECT 1027.400 3.740 1039.480 5.600 ;
  RECT 1022.200 3.740 1024.850 5.600 ;
  RECT 1007.400 3.740 1019.640 5.600 ;
  RECT 1001.000 3.740 1005.010 5.600 ;
  RECT 986.600 3.740 998.560 5.600 ;
  RECT 981.400 3.740 983.930 5.600 ;
  RECT 966.600 3.740 978.720 5.600 ;
  RECT 960.200 3.740 964.090 5.600 ;
  RECT 945.400 3.740 957.640 5.600 ;
  RECT 940.200 3.740 943.010 5.600 ;
  RECT 925.800 3.740 937.800 5.600 ;
  RECT 919.400 3.740 923.170 5.600 ;
  RECT 904.600 3.740 916.720 5.600 ;
  RECT 899.400 3.740 902.090 5.600 ;
  RECT 886.600 3.740 896.880 5.600 ;
  RECT 878.200 3.740 882.250 5.600 ;
  RECT 863.800 3.740 875.800 5.600 ;
  RECT 858.600 3.740 861.170 5.600 ;
  RECT 843.800 3.740 855.960 5.600 ;
  RECT 837.400 3.740 841.330 5.600 ;
  RECT 822.600 3.740 834.880 5.600 ;
  RECT 817.400 3.740 820.250 5.600 ;
  RECT 803.000 3.740 815.040 5.600 ;
  RECT 796.600 3.740 800.410 5.600 ;
  RECT 781.800 3.740 793.960 5.600 ;
  RECT 776.600 3.740 779.330 5.600 ;
  RECT 761.800 3.740 774.120 5.600 ;
  RECT 755.400 3.740 759.490 5.600 ;
  RECT 741.000 3.740 753.040 5.600 ;
  RECT 735.800 3.740 738.410 5.600 ;
  RECT 722.600 3.740 733.200 5.600 ;
  RECT 700.200 3.740 718.570 5.600 ;
  RECT 688.200 3.740 691.730 5.600 ;
  RECT 681.000 3.740 685.760 5.600 ;
  RECT 658.200 3.740 662.640 5.600 ;
  RECT 643.800 3.740 655.740 5.600 ;
  RECT 638.200 3.740 641.110 5.600 ;
  RECT 623.800 3.740 635.900 5.600 ;
  RECT 617.400 3.740 621.270 5.600 ;
  RECT 602.600 3.740 614.820 5.600 ;
  RECT 597.400 3.740 600.190 5.600 ;
  RECT 583.000 3.740 594.980 5.600 ;
  RECT 576.200 3.740 580.350 5.600 ;
  RECT 561.800 3.740 573.900 5.600 ;
  RECT 556.600 3.740 559.270 5.600 ;
  RECT 541.800 3.740 554.060 5.600 ;
  RECT 535.400 3.740 539.430 5.600 ;
  RECT 521.000 3.740 532.980 5.600 ;
  RECT 515.800 3.740 518.350 5.600 ;
  RECT 502.600 3.740 513.140 5.600 ;
  RECT 494.600 3.740 498.510 5.600 ;
  RECT 479.800 3.740 492.060 5.600 ;
  RECT 474.600 3.740 477.430 5.600 ;
  RECT 460.200 3.740 472.220 5.600 ;
  RECT 453.800 3.740 457.590 5.600 ;
  RECT 439.000 3.740 451.140 5.600 ;
  RECT 433.800 3.740 436.510 5.600 ;
  RECT 419.000 3.740 431.300 5.600 ;
  RECT 412.600 3.740 416.670 5.600 ;
  RECT 398.200 3.740 410.220 5.600 ;
  RECT 393.000 3.740 395.590 5.600 ;
  RECT 378.200 3.740 390.380 5.600 ;
  RECT 371.800 3.740 375.750 5.600 ;
  RECT 357.000 3.740 369.300 5.600 ;
  RECT 351.800 3.740 354.670 5.600 ;
  RECT 339.000 3.740 349.460 5.600 ;
  RECT 331.000 3.740 334.830 5.600 ;
  RECT 316.200 3.740 328.380 5.600 ;
  RECT 311.000 3.740 313.750 5.600 ;
  RECT 296.600 3.740 308.540 5.600 ;
  RECT 289.800 3.740 293.910 5.600 ;
  RECT 275.400 3.740 287.460 5.600 ;
  RECT 270.200 3.740 272.830 5.600 ;
  RECT 255.400 3.740 267.620 5.600 ;
  RECT 249.000 3.740 252.990 5.600 ;
  RECT 234.600 3.740 246.540 5.600 ;
  RECT 229.000 3.740 231.910 5.600 ;
  RECT 214.600 3.740 226.700 5.600 ;
  RECT 208.200 3.740 212.070 5.600 ;
  RECT 193.400 3.740 205.620 5.600 ;
  RECT 188.200 3.740 190.990 5.600 ;
  RECT 175.400 3.740 185.780 5.600 ;
  RECT 167.000 3.740 171.150 5.600 ;
  RECT 152.600 3.740 164.700 5.600 ;
  RECT 147.400 3.740 150.070 5.600 ;
  RECT 132.600 3.740 144.860 5.600 ;
  RECT 126.200 3.740 130.230 5.600 ;
  RECT 111.800 3.740 123.780 5.600 ;
  RECT 106.600 3.740 109.150 5.600 ;
  RECT 91.800 3.740 103.940 5.600 ;
  RECT 85.400 3.740 89.310 5.600 ;
  RECT 70.600 3.740 82.860 5.600 ;
  RECT 65.400 3.740 68.230 5.600 ;
  RECT 51.000 3.740 63.020 5.600 ;
  RECT 44.600 3.740 48.390 5.600 ;
  RECT 29.800 3.740 41.940 5.600 ;
  RECT 24.600 3.740 27.310 5.600 ;
  RECT 11.800 3.740 22.100 5.600 ;
  RECT 4.000 3.740 7.470 5.600 ;
  RECT 2.140 547.210 4.000 549.070 ;
  RECT 0.000 549.350 1.860 551.210 ;
  RECT 1375.500 3.740 1377.360 5.600 ;
  RECT 1377.640 1.600 1379.500 3.460 ;
  RECT 1375.500 547.210 1377.360 549.070 ;
  RECT 1377.640 549.350 1379.500 551.210 ;
  RECT 2.140 3.740 4.000 5.600 ;
  RECT 0.000 1.600 1.860 3.460 ;
  RECT 1367.600 0.000 1368.400 1.000 ;
  RECT 1367.900 1.000 1368.100 5.200 ;
  RECT 1367.840 5.200 1368.100 5.400 ;
  RECT 1367.840 5.400 1368.040 7.020 ;
  RECT 1352.800 0.000 1353.600 1.000 ;
  RECT 1353.100 1.000 1353.300 5.200 ;
  RECT 1353.100 5.200 1353.410 5.400 ;
  RECT 1353.210 5.400 1353.410 7.020 ;
  RECT 1347.600 0.000 1348.400 1.000 ;
  RECT 1347.900 1.000 1348.100 5.200 ;
  RECT 1347.900 5.200 1348.200 5.400 ;
  RECT 1348.000 5.400 1348.200 7.020 ;
  RECT 1333.200 0.000 1334.000 1.000 ;
  RECT 1333.500 1.000 1333.700 5.200 ;
  RECT 1333.370 5.200 1333.700 5.400 ;
  RECT 1333.370 5.400 1333.570 7.020 ;
  RECT 1326.800 0.000 1327.600 1.000 ;
  RECT 1327.100 1.000 1327.300 5.200 ;
  RECT 1326.920 5.200 1327.300 5.400 ;
  RECT 1326.920 5.400 1327.120 7.020 ;
  RECT 1312.000 0.000 1312.800 1.000 ;
  RECT 1312.300 1.000 1312.500 5.200 ;
  RECT 1312.290 5.200 1312.500 5.400 ;
  RECT 1312.290 5.400 1312.490 7.020 ;
  RECT 1306.800 0.000 1307.600 1.000 ;
  RECT 1307.100 1.000 1307.300 5.200 ;
  RECT 1307.080 5.200 1307.300 5.400 ;
  RECT 1307.080 5.400 1307.280 7.020 ;
  RECT 1292.000 0.000 1292.800 1.000 ;
  RECT 1292.300 1.000 1292.500 5.200 ;
  RECT 1292.300 5.200 1292.650 5.400 ;
  RECT 1292.450 5.400 1292.650 7.020 ;
  RECT 1285.600 0.000 1286.400 1.000 ;
  RECT 1285.900 1.000 1286.100 5.200 ;
  RECT 1285.900 5.200 1286.200 5.400 ;
  RECT 1286.000 5.400 1286.200 7.020 ;
  RECT 1271.200 0.000 1272.000 1.000 ;
  RECT 1271.500 1.000 1271.700 5.200 ;
  RECT 1271.370 5.200 1271.700 5.400 ;
  RECT 1271.370 5.400 1271.570 7.020 ;
  RECT 1266.000 0.000 1266.800 1.000 ;
  RECT 1266.300 1.000 1266.500 5.200 ;
  RECT 1266.160 5.200 1266.500 5.400 ;
  RECT 1266.160 5.400 1266.360 7.020 ;
  RECT 1251.200 0.000 1252.000 1.000 ;
  RECT 1251.500 1.000 1251.700 5.200 ;
  RECT 1251.500 5.200 1251.730 5.400 ;
  RECT 1251.530 5.400 1251.730 7.020 ;
  RECT 1244.800 0.000 1245.600 1.000 ;
  RECT 1245.100 1.000 1245.300 5.200 ;
  RECT 1245.080 5.200 1245.300 5.400 ;
  RECT 1245.080 5.400 1245.280 7.020 ;
  RECT 1230.000 0.000 1230.800 1.000 ;
  RECT 1230.300 1.000 1230.500 5.200 ;
  RECT 1230.300 5.200 1230.650 5.400 ;
  RECT 1230.450 5.400 1230.650 7.020 ;
  RECT 1224.800 0.000 1225.600 1.000 ;
  RECT 1225.100 1.000 1225.300 5.200 ;
  RECT 1225.100 5.200 1225.440 5.400 ;
  RECT 1225.240 5.400 1225.440 7.020 ;
  RECT 1212.000 0.000 1212.800 1.000 ;
  RECT 1212.300 1.000 1212.500 5.200 ;
  RECT 1212.300 5.200 1212.530 5.400 ;
  RECT 1212.330 5.400 1212.530 7.020 ;
  RECT 1210.400 0.000 1211.200 1.000 ;
  RECT 1210.700 1.000 1210.900 5.200 ;
  RECT 1210.610 5.200 1210.900 5.400 ;
  RECT 1210.610 5.400 1210.810 7.020 ;
  RECT 1204.000 0.000 1204.800 1.000 ;
  RECT 1204.300 1.000 1204.500 5.200 ;
  RECT 1204.160 5.200 1204.500 5.400 ;
  RECT 1204.160 5.400 1204.360 7.020 ;
  RECT 1189.200 0.000 1190.000 1.000 ;
  RECT 1189.500 1.000 1189.700 5.200 ;
  RECT 1189.500 5.200 1189.730 5.400 ;
  RECT 1189.530 5.400 1189.730 7.020 ;
  RECT 1184.000 0.000 1184.800 1.000 ;
  RECT 1184.300 1.000 1184.500 5.200 ;
  RECT 1184.300 5.200 1184.520 5.400 ;
  RECT 1184.320 5.400 1184.520 7.020 ;
  RECT 1169.200 0.000 1170.000 1.000 ;
  RECT 1169.500 1.000 1169.700 5.200 ;
  RECT 1169.500 5.200 1169.890 5.400 ;
  RECT 1169.690 5.400 1169.890 7.020 ;
  RECT 1162.800 0.000 1163.600 1.000 ;
  RECT 1163.100 1.000 1163.300 5.200 ;
  RECT 1163.100 5.200 1163.440 5.400 ;
  RECT 1163.240 5.400 1163.440 7.020 ;
  RECT 1148.400 0.000 1149.200 1.000 ;
  RECT 1148.700 1.000 1148.900 5.200 ;
  RECT 1148.610 5.200 1148.900 5.400 ;
  RECT 1148.610 5.400 1148.810 7.020 ;
  RECT 1143.200 0.000 1144.000 1.000 ;
  RECT 1143.500 1.000 1143.700 5.200 ;
  RECT 1143.400 5.200 1143.700 5.400 ;
  RECT 1143.400 5.400 1143.600 7.020 ;
  RECT 1128.400 0.000 1129.200 1.000 ;
  RECT 1128.700 1.000 1128.900 5.200 ;
  RECT 1128.700 5.200 1128.970 5.400 ;
  RECT 1128.770 5.400 1128.970 7.020 ;
  RECT 1122.000 0.000 1122.800 1.000 ;
  RECT 1122.300 1.000 1122.500 5.200 ;
  RECT 1122.300 5.200 1122.520 5.400 ;
  RECT 1122.320 5.400 1122.520 7.020 ;
  RECT 1107.200 0.000 1108.000 1.000 ;
  RECT 1107.500 1.000 1107.700 5.200 ;
  RECT 1107.500 5.200 1107.890 5.400 ;
  RECT 1107.690 5.400 1107.890 7.020 ;
  RECT 1102.000 0.000 1102.800 1.000 ;
  RECT 1102.300 1.000 1102.500 5.200 ;
  RECT 1102.300 5.200 1102.680 5.400 ;
  RECT 1102.480 5.400 1102.680 7.020 ;
  RECT 1087.600 0.000 1088.400 1.000 ;
  RECT 1087.900 1.000 1088.100 5.200 ;
  RECT 1087.850 5.200 1088.100 5.400 ;
  RECT 1087.850 5.400 1088.050 7.020 ;
  RECT 1081.200 0.000 1082.000 1.000 ;
  RECT 1081.500 1.000 1081.700 5.200 ;
  RECT 1081.400 5.200 1081.700 5.400 ;
  RECT 1081.400 5.400 1081.600 7.020 ;
  RECT 1066.400 0.000 1067.200 1.000 ;
  RECT 1066.700 1.000 1066.900 5.200 ;
  RECT 1066.700 5.200 1066.970 5.400 ;
  RECT 1066.770 5.400 1066.970 7.020 ;
  RECT 1061.200 0.000 1062.000 1.000 ;
  RECT 1061.500 1.000 1061.700 5.200 ;
  RECT 1061.500 5.200 1061.760 5.400 ;
  RECT 1061.560 5.400 1061.760 7.020 ;
  RECT 1048.400 0.000 1049.200 1.000 ;
  RECT 1048.700 1.000 1048.900 5.200 ;
  RECT 1048.650 5.200 1048.900 5.400 ;
  RECT 1048.650 5.400 1048.850 7.020 ;
  RECT 1046.800 0.000 1047.600 1.000 ;
  RECT 1047.100 1.000 1047.300 5.200 ;
  RECT 1046.930 5.200 1047.300 5.400 ;
  RECT 1046.930 5.400 1047.130 7.020 ;
  RECT 1040.000 0.000 1040.800 1.000 ;
  RECT 1040.300 1.000 1040.500 5.200 ;
  RECT 1040.300 5.200 1040.680 5.400 ;
  RECT 1040.480 5.400 1040.680 7.020 ;
  RECT 1025.600 0.000 1026.400 1.000 ;
  RECT 1025.900 1.000 1026.100 5.200 ;
  RECT 1025.850 5.200 1026.100 5.400 ;
  RECT 1025.850 5.400 1026.050 7.020 ;
  RECT 1020.400 0.000 1021.200 1.000 ;
  RECT 1020.700 1.000 1020.900 5.200 ;
  RECT 1020.640 5.200 1020.900 5.400 ;
  RECT 1020.640 5.400 1020.840 7.020 ;
  RECT 1005.600 0.000 1006.400 1.000 ;
  RECT 1005.900 1.000 1006.100 5.200 ;
  RECT 1005.900 5.200 1006.210 5.400 ;
  RECT 1006.010 5.400 1006.210 7.020 ;
  RECT 999.200 0.000 1000.000 1.000 ;
  RECT 999.500 1.000 999.700 5.200 ;
  RECT 999.500 5.200 999.760 5.400 ;
  RECT 999.560 5.400 999.760 7.020 ;
  RECT 984.800 0.000 985.600 1.000 ;
  RECT 985.100 1.000 985.300 5.200 ;
  RECT 984.930 5.200 985.300 5.400 ;
  RECT 984.930 5.400 985.130 7.020 ;
  RECT 979.600 0.000 980.400 1.000 ;
  RECT 979.900 1.000 980.100 5.200 ;
  RECT 979.720 5.200 980.100 5.400 ;
  RECT 979.720 5.400 979.920 7.020 ;
  RECT 964.800 0.000 965.600 1.000 ;
  RECT 965.100 1.000 965.300 5.200 ;
  RECT 965.090 5.200 965.300 5.400 ;
  RECT 965.090 5.400 965.290 7.020 ;
  RECT 958.400 0.000 959.200 1.000 ;
  RECT 958.700 1.000 958.900 5.200 ;
  RECT 958.640 5.200 958.900 5.400 ;
  RECT 958.640 5.400 958.840 7.020 ;
  RECT 943.600 0.000 944.400 1.000 ;
  RECT 943.900 1.000 944.100 5.200 ;
  RECT 943.900 5.200 944.210 5.400 ;
  RECT 944.010 5.400 944.210 7.020 ;
  RECT 938.400 0.000 939.200 1.000 ;
  RECT 938.700 1.000 938.900 5.200 ;
  RECT 938.700 5.200 939.000 5.400 ;
  RECT 938.800 5.400 939.000 7.020 ;
  RECT 924.000 0.000 924.800 1.000 ;
  RECT 924.300 1.000 924.500 5.200 ;
  RECT 924.170 5.200 924.500 5.400 ;
  RECT 924.170 5.400 924.370 7.020 ;
  RECT 917.600 0.000 918.400 1.000 ;
  RECT 917.900 1.000 918.100 5.200 ;
  RECT 917.720 5.200 918.100 5.400 ;
  RECT 917.720 5.400 917.920 7.020 ;
  RECT 902.800 0.000 903.600 1.000 ;
  RECT 903.100 1.000 903.300 5.200 ;
  RECT 903.090 5.200 903.300 5.400 ;
  RECT 903.090 5.400 903.290 7.020 ;
  RECT 897.600 0.000 898.400 1.000 ;
  RECT 897.900 1.000 898.100 5.200 ;
  RECT 897.880 5.200 898.100 5.400 ;
  RECT 897.880 5.400 898.080 7.020 ;
  RECT 884.800 0.000 885.600 1.000 ;
  RECT 885.100 1.000 885.300 5.200 ;
  RECT 884.970 5.200 885.300 5.400 ;
  RECT 884.970 5.400 885.170 7.020 ;
  RECT 882.800 0.000 883.600 1.000 ;
  RECT 883.100 1.000 883.300 5.200 ;
  RECT 883.100 5.200 883.450 5.400 ;
  RECT 883.250 5.400 883.450 7.020 ;
  RECT 876.400 0.000 877.200 1.000 ;
  RECT 876.700 1.000 876.900 5.200 ;
  RECT 876.700 5.200 877.000 5.400 ;
  RECT 876.800 5.400 877.000 7.020 ;
  RECT 862.000 0.000 862.800 1.000 ;
  RECT 862.300 1.000 862.500 5.200 ;
  RECT 862.170 5.200 862.500 5.400 ;
  RECT 862.170 5.400 862.370 7.020 ;
  RECT 856.800 0.000 857.600 1.000 ;
  RECT 857.100 1.000 857.300 5.200 ;
  RECT 856.960 5.200 857.300 5.400 ;
  RECT 856.960 5.400 857.160 7.020 ;
  RECT 842.000 0.000 842.800 1.000 ;
  RECT 842.300 1.000 842.500 5.200 ;
  RECT 842.300 5.200 842.530 5.400 ;
  RECT 842.330 5.400 842.530 7.020 ;
  RECT 835.600 0.000 836.400 1.000 ;
  RECT 835.900 1.000 836.100 5.200 ;
  RECT 835.880 5.200 836.100 5.400 ;
  RECT 835.880 5.400 836.080 7.020 ;
  RECT 820.800 0.000 821.600 1.000 ;
  RECT 821.100 1.000 821.300 5.200 ;
  RECT 821.100 5.200 821.450 5.400 ;
  RECT 821.250 5.400 821.450 7.020 ;
  RECT 815.600 0.000 816.400 1.000 ;
  RECT 815.900 1.000 816.100 5.200 ;
  RECT 815.900 5.200 816.240 5.400 ;
  RECT 816.040 5.400 816.240 7.020 ;
  RECT 801.200 0.000 802.000 1.000 ;
  RECT 801.500 1.000 801.700 5.200 ;
  RECT 801.410 5.200 801.700 5.400 ;
  RECT 801.410 5.400 801.610 7.020 ;
  RECT 794.800 0.000 795.600 1.000 ;
  RECT 795.100 1.000 795.300 5.200 ;
  RECT 794.960 5.200 795.300 5.400 ;
  RECT 794.960 5.400 795.160 7.020 ;
  RECT 780.000 0.000 780.800 1.000 ;
  RECT 780.300 1.000 780.500 5.200 ;
  RECT 780.300 5.200 780.530 5.400 ;
  RECT 780.330 5.400 780.530 7.020 ;
  RECT 774.800 0.000 775.600 1.000 ;
  RECT 775.100 1.000 775.300 5.200 ;
  RECT 775.100 5.200 775.320 5.400 ;
  RECT 775.120 5.400 775.320 7.020 ;
  RECT 760.000 0.000 760.800 1.000 ;
  RECT 760.300 1.000 760.500 5.200 ;
  RECT 760.300 5.200 760.690 5.400 ;
  RECT 760.490 5.400 760.690 7.020 ;
  RECT 753.600 0.000 754.400 1.000 ;
  RECT 753.900 1.000 754.100 5.200 ;
  RECT 753.900 5.200 754.240 5.400 ;
  RECT 754.040 5.400 754.240 7.020 ;
  RECT 739.200 0.000 740.000 1.000 ;
  RECT 739.500 1.000 739.700 5.200 ;
  RECT 739.410 5.200 739.700 5.400 ;
  RECT 739.410 5.400 739.610 7.020 ;
  RECT 734.000 0.000 734.800 1.000 ;
  RECT 734.300 1.000 734.500 5.200 ;
  RECT 734.200 5.200 734.500 5.400 ;
  RECT 734.200 5.400 734.400 7.020 ;
  RECT 720.800 0.000 721.600 1.000 ;
  RECT 721.100 1.000 721.300 5.200 ;
  RECT 721.100 5.200 721.490 5.400 ;
  RECT 721.290 5.400 721.490 7.020 ;
  RECT 719.200 0.000 720.000 1.000 ;
  RECT 719.500 1.000 719.700 5.200 ;
  RECT 719.500 5.200 719.770 5.400 ;
  RECT 719.570 5.400 719.770 7.020 ;
  RECT 698.400 0.000 699.200 1.000 ;
  RECT 698.700 1.000 698.900 5.200 ;
  RECT 698.700 5.200 699.000 5.400 ;
  RECT 698.800 5.400 699.000 7.020 ;
  RECT 697.200 0.000 698.000 1.000 ;
  RECT 697.500 1.000 697.700 5.200 ;
  RECT 697.500 5.200 697.850 5.400 ;
  RECT 697.650 5.400 697.850 7.020 ;
  RECT 696.000 0.000 696.800 1.000 ;
  RECT 696.300 1.000 696.500 5.200 ;
  RECT 696.300 5.200 696.680 5.400 ;
  RECT 696.480 5.400 696.680 7.020 ;
  RECT 694.800 0.000 695.600 1.000 ;
  RECT 695.100 1.000 695.300 5.200 ;
  RECT 695.100 5.200 695.430 5.400 ;
  RECT 695.230 5.400 695.430 7.020 ;
  RECT 693.600 0.000 694.400 1.000 ;
  RECT 693.900 1.000 694.100 5.200 ;
  RECT 693.900 5.200 694.180 5.400 ;
  RECT 693.980 5.400 694.180 7.020 ;
  RECT 692.400 0.000 693.200 1.000 ;
  RECT 692.700 1.000 692.900 5.200 ;
  RECT 692.700 5.200 692.930 5.400 ;
  RECT 692.730 5.400 692.930 7.020 ;
  RECT 686.400 0.000 687.200 1.000 ;
  RECT 686.700 1.000 686.900 5.200 ;
  RECT 686.700 5.200 686.960 5.400 ;
  RECT 686.760 5.400 686.960 7.020 ;
  RECT 679.200 0.000 680.000 1.000 ;
  RECT 679.500 1.000 679.700 5.200 ;
  RECT 679.460 5.200 679.700 5.400 ;
  RECT 679.460 5.400 679.660 7.020 ;
  RECT 676.800 0.000 677.600 1.000 ;
  RECT 677.100 1.000 677.300 5.200 ;
  RECT 676.980 5.200 677.300 5.400 ;
  RECT 676.980 5.400 677.180 7.020 ;
  RECT 674.000 0.000 674.800 1.000 ;
  RECT 674.300 1.000 674.500 5.200 ;
  RECT 674.120 5.200 674.500 5.400 ;
  RECT 674.120 5.400 674.320 7.020 ;
  RECT 671.200 0.000 672.000 1.000 ;
  RECT 671.500 1.000 671.700 5.200 ;
  RECT 671.500 5.200 671.840 5.400 ;
  RECT 671.640 5.400 671.840 7.020 ;
  RECT 670.000 0.000 670.800 1.000 ;
  RECT 670.300 1.000 670.500 5.200 ;
  RECT 670.120 5.200 670.500 5.400 ;
  RECT 670.120 5.400 670.320 7.020 ;
  RECT 667.200 0.000 668.000 1.000 ;
  RECT 667.500 1.000 667.700 5.200 ;
  RECT 667.500 5.200 667.840 5.400 ;
  RECT 667.640 5.400 667.840 7.020 ;
  RECT 666.000 0.000 666.800 1.000 ;
  RECT 666.300 1.000 666.500 5.200 ;
  RECT 666.120 5.200 666.500 5.400 ;
  RECT 666.120 5.400 666.320 7.020 ;
  RECT 663.200 0.000 664.000 1.000 ;
  RECT 663.500 1.000 663.700 5.200 ;
  RECT 663.500 5.200 663.840 5.400 ;
  RECT 663.640 5.400 663.840 7.020 ;
  RECT 656.400 0.000 657.200 1.000 ;
  RECT 656.700 1.000 656.900 5.200 ;
  RECT 656.700 5.200 656.940 5.400 ;
  RECT 656.740 5.400 656.940 7.020 ;
  RECT 642.000 0.000 642.800 1.000 ;
  RECT 642.300 1.000 642.500 5.200 ;
  RECT 642.110 5.200 642.500 5.400 ;
  RECT 642.110 5.400 642.310 7.020 ;
  RECT 636.400 0.000 637.200 1.000 ;
  RECT 636.700 1.000 636.900 5.200 ;
  RECT 636.700 5.200 637.100 5.400 ;
  RECT 636.900 5.400 637.100 7.020 ;
  RECT 622.000 0.000 622.800 1.000 ;
  RECT 622.300 1.000 622.500 5.200 ;
  RECT 622.270 5.200 622.500 5.400 ;
  RECT 622.270 5.400 622.470 7.020 ;
  RECT 615.600 0.000 616.400 1.000 ;
  RECT 615.900 1.000 616.100 5.200 ;
  RECT 615.820 5.200 616.100 5.400 ;
  RECT 615.820 5.400 616.020 7.020 ;
  RECT 600.800 0.000 601.600 1.000 ;
  RECT 601.100 1.000 601.300 5.200 ;
  RECT 601.100 5.200 601.390 5.400 ;
  RECT 601.190 5.400 601.390 7.020 ;
  RECT 595.600 0.000 596.400 1.000 ;
  RECT 595.900 1.000 596.100 5.200 ;
  RECT 595.900 5.200 596.180 5.400 ;
  RECT 595.980 5.400 596.180 7.020 ;
  RECT 581.200 0.000 582.000 1.000 ;
  RECT 581.500 1.000 581.700 5.200 ;
  RECT 581.350 5.200 581.700 5.400 ;
  RECT 581.350 5.400 581.550 7.020 ;
  RECT 574.400 0.000 575.200 1.000 ;
  RECT 574.700 1.000 574.900 5.200 ;
  RECT 574.700 5.200 575.100 5.400 ;
  RECT 574.900 5.400 575.100 7.020 ;
  RECT 560.000 0.000 560.800 1.000 ;
  RECT 560.300 1.000 560.500 5.200 ;
  RECT 560.270 5.200 560.500 5.400 ;
  RECT 560.270 5.400 560.470 7.020 ;
  RECT 554.800 0.000 555.600 1.000 ;
  RECT 555.100 1.000 555.300 5.200 ;
  RECT 555.060 5.200 555.300 5.400 ;
  RECT 555.060 5.400 555.260 7.020 ;
  RECT 540.000 0.000 540.800 1.000 ;
  RECT 540.300 1.000 540.500 5.200 ;
  RECT 540.300 5.200 540.630 5.400 ;
  RECT 540.430 5.400 540.630 7.020 ;
  RECT 533.600 0.000 534.400 1.000 ;
  RECT 533.900 1.000 534.100 5.200 ;
  RECT 533.900 5.200 534.180 5.400 ;
  RECT 533.980 5.400 534.180 7.020 ;
  RECT 519.200 0.000 520.000 1.000 ;
  RECT 519.500 1.000 519.700 5.200 ;
  RECT 519.350 5.200 519.700 5.400 ;
  RECT 519.350 5.400 519.550 7.020 ;
  RECT 514.000 0.000 514.800 1.000 ;
  RECT 514.300 1.000 514.500 5.200 ;
  RECT 514.140 5.200 514.500 5.400 ;
  RECT 514.140 5.400 514.340 7.020 ;
  RECT 500.800 0.000 501.600 1.000 ;
  RECT 501.100 1.000 501.300 5.200 ;
  RECT 501.100 5.200 501.430 5.400 ;
  RECT 501.230 5.400 501.430 7.020 ;
  RECT 499.200 0.000 500.000 1.000 ;
  RECT 499.500 1.000 499.700 5.200 ;
  RECT 499.500 5.200 499.710 5.400 ;
  RECT 499.510 5.400 499.710 7.020 ;
  RECT 492.800 0.000 493.600 1.000 ;
  RECT 493.100 1.000 493.300 5.200 ;
  RECT 493.060 5.200 493.300 5.400 ;
  RECT 493.060 5.400 493.260 7.020 ;
  RECT 478.000 0.000 478.800 1.000 ;
  RECT 478.300 1.000 478.500 5.200 ;
  RECT 478.300 5.200 478.630 5.400 ;
  RECT 478.430 5.400 478.630 7.020 ;
  RECT 472.800 0.000 473.600 1.000 ;
  RECT 473.100 1.000 473.300 5.200 ;
  RECT 473.100 5.200 473.420 5.400 ;
  RECT 473.220 5.400 473.420 7.020 ;
  RECT 458.400 0.000 459.200 1.000 ;
  RECT 458.700 1.000 458.900 5.200 ;
  RECT 458.590 5.200 458.900 5.400 ;
  RECT 458.590 5.400 458.790 7.020 ;
  RECT 452.000 0.000 452.800 1.000 ;
  RECT 452.300 1.000 452.500 5.200 ;
  RECT 452.140 5.200 452.500 5.400 ;
  RECT 452.140 5.400 452.340 7.020 ;
  RECT 437.200 0.000 438.000 1.000 ;
  RECT 437.500 1.000 437.700 5.200 ;
  RECT 437.500 5.200 437.710 5.400 ;
  RECT 437.510 5.400 437.710 7.020 ;
  RECT 432.000 0.000 432.800 1.000 ;
  RECT 432.300 1.000 432.500 5.200 ;
  RECT 432.300 5.200 432.500 5.400 ;
  RECT 432.300 5.400 432.500 7.020 ;
  RECT 417.200 0.000 418.000 1.000 ;
  RECT 417.500 1.000 417.700 5.200 ;
  RECT 417.500 5.200 417.870 5.400 ;
  RECT 417.670 5.400 417.870 7.020 ;
  RECT 410.800 0.000 411.600 1.000 ;
  RECT 411.100 1.000 411.300 5.200 ;
  RECT 411.100 5.200 411.420 5.400 ;
  RECT 411.220 5.400 411.420 7.020 ;
  RECT 396.400 0.000 397.200 1.000 ;
  RECT 396.700 1.000 396.900 5.200 ;
  RECT 396.590 5.200 396.900 5.400 ;
  RECT 396.590 5.400 396.790 7.020 ;
  RECT 391.200 0.000 392.000 1.000 ;
  RECT 391.500 1.000 391.700 5.200 ;
  RECT 391.380 5.200 391.700 5.400 ;
  RECT 391.380 5.400 391.580 7.020 ;
  RECT 376.400 0.000 377.200 1.000 ;
  RECT 376.700 1.000 376.900 5.200 ;
  RECT 376.700 5.200 376.950 5.400 ;
  RECT 376.750 5.400 376.950 7.020 ;
  RECT 370.000 0.000 370.800 1.000 ;
  RECT 370.300 1.000 370.500 5.200 ;
  RECT 370.300 5.200 370.500 5.400 ;
  RECT 370.300 5.400 370.500 7.020 ;
  RECT 355.200 0.000 356.000 1.000 ;
  RECT 355.500 1.000 355.700 5.200 ;
  RECT 355.500 5.200 355.870 5.400 ;
  RECT 355.670 5.400 355.870 7.020 ;
  RECT 350.000 0.000 350.800 1.000 ;
  RECT 350.300 1.000 350.500 5.200 ;
  RECT 350.300 5.200 350.660 5.400 ;
  RECT 350.460 5.400 350.660 7.020 ;
  RECT 337.200 0.000 338.000 1.000 ;
  RECT 337.500 1.000 337.700 5.200 ;
  RECT 337.500 5.200 337.750 5.400 ;
  RECT 337.550 5.400 337.750 7.020 ;
  RECT 335.600 0.000 336.400 1.000 ;
  RECT 335.900 1.000 336.100 5.200 ;
  RECT 335.830 5.200 336.100 5.400 ;
  RECT 335.830 5.400 336.030 7.020 ;
  RECT 329.200 0.000 330.000 1.000 ;
  RECT 329.500 1.000 329.700 5.200 ;
  RECT 329.380 5.200 329.700 5.400 ;
  RECT 329.380 5.400 329.580 7.020 ;
  RECT 314.400 0.000 315.200 1.000 ;
  RECT 314.700 1.000 314.900 5.200 ;
  RECT 314.700 5.200 314.950 5.400 ;
  RECT 314.750 5.400 314.950 7.020 ;
  RECT 309.200 0.000 310.000 1.000 ;
  RECT 309.500 1.000 309.700 5.200 ;
  RECT 309.500 5.200 309.740 5.400 ;
  RECT 309.540 5.400 309.740 7.020 ;
  RECT 294.800 0.000 295.600 1.000 ;
  RECT 295.100 1.000 295.300 5.200 ;
  RECT 294.910 5.200 295.300 5.400 ;
  RECT 294.910 5.400 295.110 7.020 ;
  RECT 288.000 0.000 288.800 1.000 ;
  RECT 288.300 1.000 288.500 5.200 ;
  RECT 288.300 5.200 288.660 5.400 ;
  RECT 288.460 5.400 288.660 7.020 ;
  RECT 273.600 0.000 274.400 1.000 ;
  RECT 273.900 1.000 274.100 5.200 ;
  RECT 273.830 5.200 274.100 5.400 ;
  RECT 273.830 5.400 274.030 7.020 ;
  RECT 268.400 0.000 269.200 1.000 ;
  RECT 268.700 1.000 268.900 5.200 ;
  RECT 268.620 5.200 268.900 5.400 ;
  RECT 268.620 5.400 268.820 7.020 ;
  RECT 253.600 0.000 254.400 1.000 ;
  RECT 253.900 1.000 254.100 5.200 ;
  RECT 253.900 5.200 254.190 5.400 ;
  RECT 253.990 5.400 254.190 7.020 ;
  RECT 247.200 0.000 248.000 1.000 ;
  RECT 247.500 1.000 247.700 5.200 ;
  RECT 247.500 5.200 247.740 5.400 ;
  RECT 247.540 5.400 247.740 7.020 ;
  RECT 232.800 0.000 233.600 1.000 ;
  RECT 233.100 1.000 233.300 5.200 ;
  RECT 232.910 5.200 233.300 5.400 ;
  RECT 232.910 5.400 233.110 7.020 ;
  RECT 227.200 0.000 228.000 1.000 ;
  RECT 227.500 1.000 227.700 5.200 ;
  RECT 227.500 5.200 227.900 5.400 ;
  RECT 227.700 5.400 227.900 7.020 ;
  RECT 212.800 0.000 213.600 1.000 ;
  RECT 213.100 1.000 213.300 5.200 ;
  RECT 213.070 5.200 213.300 5.400 ;
  RECT 213.070 5.400 213.270 7.020 ;
  RECT 206.400 0.000 207.200 1.000 ;
  RECT 206.700 1.000 206.900 5.200 ;
  RECT 206.620 5.200 206.900 5.400 ;
  RECT 206.620 5.400 206.820 7.020 ;
  RECT 191.600 0.000 192.400 1.000 ;
  RECT 191.900 1.000 192.100 5.200 ;
  RECT 191.900 5.200 192.190 5.400 ;
  RECT 191.990 5.400 192.190 7.020 ;
  RECT 186.400 0.000 187.200 1.000 ;
  RECT 186.700 1.000 186.900 5.200 ;
  RECT 186.700 5.200 186.980 5.400 ;
  RECT 186.780 5.400 186.980 7.020 ;
  RECT 173.600 0.000 174.400 1.000 ;
  RECT 173.900 1.000 174.100 5.200 ;
  RECT 173.870 5.200 174.100 5.400 ;
  RECT 173.870 5.400 174.070 7.020 ;
  RECT 172.000 0.000 172.800 1.000 ;
  RECT 172.300 1.000 172.500 5.200 ;
  RECT 172.150 5.200 172.500 5.400 ;
  RECT 172.150 5.400 172.350 7.020 ;
  RECT 165.200 0.000 166.000 1.000 ;
  RECT 165.500 1.000 165.700 5.200 ;
  RECT 165.500 5.200 165.900 5.400 ;
  RECT 165.700 5.400 165.900 7.020 ;
  RECT 150.800 0.000 151.600 1.000 ;
  RECT 151.100 1.000 151.300 5.200 ;
  RECT 151.070 5.200 151.300 5.400 ;
  RECT 151.070 5.400 151.270 7.020 ;
  RECT 145.600 0.000 146.400 1.000 ;
  RECT 145.900 1.000 146.100 5.200 ;
  RECT 145.860 5.200 146.100 5.400 ;
  RECT 145.860 5.400 146.060 7.020 ;
  RECT 130.800 0.000 131.600 1.000 ;
  RECT 131.100 1.000 131.300 5.200 ;
  RECT 131.100 5.200 131.430 5.400 ;
  RECT 131.230 5.400 131.430 7.020 ;
  RECT 124.400 0.000 125.200 1.000 ;
  RECT 124.700 1.000 124.900 5.200 ;
  RECT 124.700 5.200 124.980 5.400 ;
  RECT 124.780 5.400 124.980 7.020 ;
  RECT 110.000 0.000 110.800 1.000 ;
  RECT 110.300 1.000 110.500 5.200 ;
  RECT 110.150 5.200 110.500 5.400 ;
  RECT 110.150 5.400 110.350 7.020 ;
  RECT 104.800 0.000 105.600 1.000 ;
  RECT 105.100 1.000 105.300 5.200 ;
  RECT 104.940 5.200 105.300 5.400 ;
  RECT 104.940 5.400 105.140 7.020 ;
  RECT 90.000 0.000 90.800 1.000 ;
  RECT 90.300 1.000 90.500 5.200 ;
  RECT 90.300 5.200 90.510 5.400 ;
  RECT 90.310 5.400 90.510 7.020 ;
  RECT 83.600 0.000 84.400 1.000 ;
  RECT 83.900 1.000 84.100 5.200 ;
  RECT 83.860 5.200 84.100 5.400 ;
  RECT 83.860 5.400 84.060 7.020 ;
  RECT 68.800 0.000 69.600 1.000 ;
  RECT 69.100 1.000 69.300 5.200 ;
  RECT 69.100 5.200 69.430 5.400 ;
  RECT 69.230 5.400 69.430 7.020 ;
  RECT 63.600 0.000 64.400 1.000 ;
  RECT 63.900 1.000 64.100 5.200 ;
  RECT 63.900 5.200 64.220 5.400 ;
  RECT 64.020 5.400 64.220 7.020 ;
  RECT 49.200 0.000 50.000 1.000 ;
  RECT 49.500 1.000 49.700 5.200 ;
  RECT 49.390 5.200 49.700 5.400 ;
  RECT 49.390 5.400 49.590 7.020 ;
  RECT 42.800 0.000 43.600 1.000 ;
  RECT 43.100 1.000 43.300 5.200 ;
  RECT 42.940 5.200 43.300 5.400 ;
  RECT 42.940 5.400 43.140 7.020 ;
  RECT 28.000 0.000 28.800 1.000 ;
  RECT 28.300 1.000 28.500 5.200 ;
  RECT 28.300 5.200 28.510 5.400 ;
  RECT 28.310 5.400 28.510 7.020 ;
  RECT 22.800 0.000 23.600 1.000 ;
  RECT 23.100 1.000 23.300 5.200 ;
  RECT 23.100 5.200 23.300 5.400 ;
  RECT 23.100 5.400 23.300 7.020 ;
  RECT 10.000 0.000 10.800 1.000 ;
  RECT 10.300 1.000 10.500 5.200 ;
  RECT 10.190 5.200 10.500 5.400 ;
  RECT 10.190 5.400 10.390 7.020 ;
  RECT 8.000 0.000 8.800 1.000 ;
  RECT 8.300 1.000 8.500 5.200 ;
  RECT 8.300 5.200 8.670 5.400 ;
  RECT 8.470 5.400 8.670 7.020 ;
  RECT 1374.080 9.570 1375.220 11.170 ;
  RECT 1374.080 14.200 1375.220 15.200 ;
  RECT 1374.080 18.730 1375.220 19.730 ;
  RECT 1374.080 21.230 1375.220 22.070 ;
  RECT 1374.080 24.170 1375.220 25.170 ;
  RECT 1374.080 36.320 1375.220 37.320 ;
  RECT 1374.080 39.480 1375.220 40.080 ;
  RECT 1374.080 45.560 1375.220 46.160 ;
  RECT 1374.080 57.100 1375.220 61.420 ;
  RECT 4.280 57.100 5.420 61.420 ;
  RECT 4.280 45.560 5.420 46.160 ;
  RECT 4.280 39.480 5.420 40.080 ;
  RECT 4.280 36.320 5.420 37.320 ;
  RECT 4.280 24.170 5.420 25.170 ;
  RECT 4.280 21.230 5.420 22.070 ;
  RECT 4.280 18.730 5.420 19.730 ;
  RECT 4.280 14.200 5.420 15.200 ;
  RECT 4.280 9.570 5.420 11.170 ;
  RECT 1374.080 545.220 1375.220 545.600 ;
  RECT 1374.080 537.300 1375.220 537.580 ;
  RECT 1374.080 533.620 1375.220 533.900 ;
  RECT 1374.080 529.940 1375.220 530.220 ;
  RECT 1374.080 526.260 1375.220 526.540 ;
  RECT 1374.080 522.580 1375.220 522.860 ;
  RECT 1374.080 518.900 1375.220 519.180 ;
  RECT 1374.080 515.220 1375.220 515.500 ;
  RECT 1374.080 511.540 1375.220 511.820 ;
  RECT 1374.080 507.860 1375.220 508.140 ;
  RECT 1374.080 504.180 1375.220 504.460 ;
  RECT 1374.080 500.500 1375.220 500.780 ;
  RECT 1374.080 496.820 1375.220 497.100 ;
  RECT 1374.080 493.140 1375.220 493.420 ;
  RECT 1374.080 489.460 1375.220 489.740 ;
  RECT 1374.080 485.780 1375.220 486.060 ;
  RECT 1374.080 482.100 1375.220 482.380 ;
  RECT 1374.080 478.420 1375.220 478.700 ;
  RECT 1374.080 474.740 1375.220 475.020 ;
  RECT 1374.080 471.060 1375.220 471.340 ;
  RECT 1374.080 467.380 1375.220 467.660 ;
  RECT 1374.080 463.700 1375.220 463.980 ;
  RECT 1374.080 460.020 1375.220 460.300 ;
  RECT 1374.080 456.340 1375.220 456.620 ;
  RECT 1374.080 452.660 1375.220 452.940 ;
  RECT 1374.080 448.980 1375.220 449.260 ;
  RECT 1374.080 445.300 1375.220 445.580 ;
  RECT 1374.080 441.620 1375.220 441.900 ;
  RECT 1374.080 437.940 1375.220 438.220 ;
  RECT 1374.080 434.260 1375.220 434.540 ;
  RECT 1374.080 430.580 1375.220 430.860 ;
  RECT 1374.080 426.900 1375.220 427.180 ;
  RECT 1374.080 423.220 1375.220 423.500 ;
  RECT 1374.080 419.540 1375.220 419.820 ;
  RECT 1374.080 415.860 1375.220 416.140 ;
  RECT 1374.080 412.180 1375.220 412.460 ;
  RECT 1374.080 408.500 1375.220 408.780 ;
  RECT 1374.080 404.820 1375.220 405.100 ;
  RECT 1374.080 401.140 1375.220 401.420 ;
  RECT 1374.080 397.460 1375.220 397.740 ;
  RECT 1374.080 393.780 1375.220 394.060 ;
  RECT 1374.080 390.100 1375.220 390.380 ;
  RECT 1374.080 386.420 1375.220 386.700 ;
  RECT 1374.080 382.740 1375.220 383.020 ;
  RECT 1374.080 379.060 1375.220 379.340 ;
  RECT 1374.080 375.380 1375.220 375.660 ;
  RECT 1374.080 371.700 1375.220 371.980 ;
  RECT 1374.080 368.020 1375.220 368.300 ;
  RECT 1374.080 364.340 1375.220 364.620 ;
  RECT 1374.080 360.660 1375.220 360.940 ;
  RECT 1374.080 356.980 1375.220 357.260 ;
  RECT 1374.080 353.300 1375.220 353.580 ;
  RECT 1374.080 349.620 1375.220 349.900 ;
  RECT 1374.080 345.940 1375.220 346.220 ;
  RECT 1374.080 342.260 1375.220 342.540 ;
  RECT 1374.080 338.580 1375.220 338.860 ;
  RECT 1374.080 334.900 1375.220 335.180 ;
  RECT 1374.080 331.220 1375.220 331.500 ;
  RECT 1374.080 327.540 1375.220 327.820 ;
  RECT 1374.080 323.860 1375.220 324.140 ;
  RECT 1374.080 320.180 1375.220 320.460 ;
  RECT 1374.080 316.500 1375.220 316.780 ;
  RECT 1374.080 312.820 1375.220 313.100 ;
  RECT 1374.080 309.140 1375.220 309.420 ;
  RECT 1374.080 305.460 1375.220 305.740 ;
  RECT 1374.080 301.780 1375.220 302.060 ;
  RECT 1374.080 298.100 1375.220 298.380 ;
  RECT 1374.080 294.420 1375.220 294.700 ;
  RECT 1374.080 290.740 1375.220 291.020 ;
  RECT 1374.080 287.060 1375.220 287.340 ;
  RECT 1374.080 283.380 1375.220 283.660 ;
  RECT 1374.080 279.700 1375.220 279.980 ;
  RECT 1374.080 276.020 1375.220 276.300 ;
  RECT 1374.080 272.340 1375.220 272.620 ;
  RECT 1374.080 268.660 1375.220 268.940 ;
  RECT 1374.080 264.980 1375.220 265.260 ;
  RECT 1374.080 261.300 1375.220 261.580 ;
  RECT 1374.080 257.620 1375.220 257.900 ;
  RECT 1374.080 253.940 1375.220 254.220 ;
  RECT 1374.080 250.260 1375.220 250.540 ;
  RECT 1374.080 246.580 1375.220 246.860 ;
  RECT 1374.080 242.900 1375.220 243.180 ;
  RECT 1374.080 239.220 1375.220 239.500 ;
  RECT 1374.080 235.540 1375.220 235.820 ;
  RECT 1374.080 231.860 1375.220 232.140 ;
  RECT 1374.080 228.180 1375.220 228.460 ;
  RECT 1374.080 224.500 1375.220 224.780 ;
  RECT 1374.080 220.820 1375.220 221.100 ;
  RECT 1374.080 217.140 1375.220 217.420 ;
  RECT 1374.080 213.460 1375.220 213.740 ;
  RECT 1374.080 209.780 1375.220 210.060 ;
  RECT 1374.080 206.100 1375.220 206.380 ;
  RECT 1374.080 202.420 1375.220 202.700 ;
  RECT 1374.080 198.740 1375.220 199.020 ;
  RECT 1374.080 195.060 1375.220 195.340 ;
  RECT 1374.080 191.380 1375.220 191.660 ;
  RECT 1374.080 187.700 1375.220 187.980 ;
  RECT 1374.080 184.020 1375.220 184.300 ;
  RECT 1374.080 180.340 1375.220 180.620 ;
  RECT 1374.080 176.660 1375.220 176.940 ;
  RECT 1374.080 172.980 1375.220 173.260 ;
  RECT 1374.080 169.300 1375.220 169.580 ;
  RECT 1374.080 165.620 1375.220 165.900 ;
  RECT 1374.080 161.940 1375.220 162.220 ;
  RECT 1374.080 158.260 1375.220 158.540 ;
  RECT 1374.080 154.580 1375.220 154.860 ;
  RECT 1374.080 150.900 1375.220 151.180 ;
  RECT 1374.080 147.220 1375.220 147.500 ;
  RECT 1374.080 143.540 1375.220 143.820 ;
  RECT 1374.080 139.860 1375.220 140.140 ;
  RECT 1374.080 136.180 1375.220 136.460 ;
  RECT 1374.080 132.500 1375.220 132.780 ;
  RECT 1374.080 128.820 1375.220 129.100 ;
  RECT 1374.080 125.140 1375.220 125.420 ;
  RECT 1374.080 121.460 1375.220 121.740 ;
  RECT 1374.080 117.780 1375.220 118.060 ;
  RECT 1374.080 114.100 1375.220 114.380 ;
  RECT 1374.080 110.420 1375.220 110.700 ;
  RECT 1374.080 106.740 1375.220 107.020 ;
  RECT 1374.080 103.060 1375.220 103.340 ;
  RECT 1374.080 99.380 1375.220 99.660 ;
  RECT 1374.080 95.700 1375.220 95.980 ;
  RECT 1374.080 92.020 1375.220 92.300 ;
  RECT 1374.080 88.340 1375.220 88.620 ;
  RECT 1374.080 84.660 1375.220 84.940 ;
  RECT 1374.080 80.980 1375.220 81.260 ;
  RECT 1374.080 77.300 1375.220 77.580 ;
  RECT 1374.080 73.620 1375.220 73.900 ;
  RECT 1374.080 69.940 1375.220 70.220 ;
  RECT 1374.080 65.600 1375.220 65.980 ;
  RECT 718.100 545.790 718.350 546.930 ;
  RECT 759.020 545.790 759.270 546.930 ;
  RECT 799.940 545.790 800.190 546.930 ;
  RECT 840.860 545.790 841.110 546.930 ;
  RECT 881.780 545.790 882.030 546.930 ;
  RECT 922.700 545.790 922.950 546.930 ;
  RECT 963.620 545.790 963.870 546.930 ;
  RECT 1004.540 545.790 1004.790 546.930 ;
  RECT 1045.460 545.790 1045.710 546.930 ;
  RECT 1086.380 545.790 1086.630 546.930 ;
  RECT 1127.300 545.790 1127.550 546.930 ;
  RECT 1168.220 545.790 1168.470 546.930 ;
  RECT 1209.140 545.790 1209.390 546.930 ;
  RECT 1250.060 545.790 1250.310 546.930 ;
  RECT 1290.980 545.790 1291.230 546.930 ;
  RECT 1331.900 545.790 1332.150 546.930 ;
  RECT 701.090 545.790 703.600 546.930 ;
  RECT 688.670 545.790 691.060 546.930 ;
  RECT 681.160 545.790 684.220 546.930 ;
  RECT 705.340 545.790 708.190 546.930 ;
  RECT 709.640 545.790 712.890 546.930 ;
  RECT 678.440 545.790 680.200 546.930 ;
  RECT 673.100 545.790 674.860 546.930 ;
  RECT 669.100 545.790 670.860 546.930 ;
  RECT 665.100 545.790 666.860 546.930 ;
  RECT 4.280 65.600 5.420 65.980 ;
  RECT 4.280 69.940 5.420 70.220 ;
  RECT 4.280 73.620 5.420 73.900 ;
  RECT 4.280 77.300 5.420 77.580 ;
  RECT 4.280 80.980 5.420 81.260 ;
  RECT 4.280 84.660 5.420 84.940 ;
  RECT 4.280 88.340 5.420 88.620 ;
  RECT 4.280 92.020 5.420 92.300 ;
  RECT 4.280 95.700 5.420 95.980 ;
  RECT 4.280 99.380 5.420 99.660 ;
  RECT 4.280 103.060 5.420 103.340 ;
  RECT 4.280 106.740 5.420 107.020 ;
  RECT 4.280 110.420 5.420 110.700 ;
  RECT 4.280 114.100 5.420 114.380 ;
  RECT 4.280 117.780 5.420 118.060 ;
  RECT 4.280 121.460 5.420 121.740 ;
  RECT 4.280 125.140 5.420 125.420 ;
  RECT 4.280 128.820 5.420 129.100 ;
  RECT 4.280 132.500 5.420 132.780 ;
  RECT 4.280 136.180 5.420 136.460 ;
  RECT 4.280 139.860 5.420 140.140 ;
  RECT 4.280 143.540 5.420 143.820 ;
  RECT 4.280 147.220 5.420 147.500 ;
  RECT 4.280 150.900 5.420 151.180 ;
  RECT 4.280 154.580 5.420 154.860 ;
  RECT 4.280 158.260 5.420 158.540 ;
  RECT 4.280 161.940 5.420 162.220 ;
  RECT 4.280 165.620 5.420 165.900 ;
  RECT 4.280 169.300 5.420 169.580 ;
  RECT 4.280 172.980 5.420 173.260 ;
  RECT 4.280 176.660 5.420 176.940 ;
  RECT 4.280 180.340 5.420 180.620 ;
  RECT 4.280 184.020 5.420 184.300 ;
  RECT 4.280 187.700 5.420 187.980 ;
  RECT 4.280 191.380 5.420 191.660 ;
  RECT 4.280 195.060 5.420 195.340 ;
  RECT 4.280 198.740 5.420 199.020 ;
  RECT 4.280 202.420 5.420 202.700 ;
  RECT 4.280 206.100 5.420 206.380 ;
  RECT 4.280 209.780 5.420 210.060 ;
  RECT 4.280 213.460 5.420 213.740 ;
  RECT 4.280 217.140 5.420 217.420 ;
  RECT 4.280 220.820 5.420 221.100 ;
  RECT 4.280 224.500 5.420 224.780 ;
  RECT 4.280 228.180 5.420 228.460 ;
  RECT 4.280 231.860 5.420 232.140 ;
  RECT 4.280 235.540 5.420 235.820 ;
  RECT 4.280 239.220 5.420 239.500 ;
  RECT 4.280 242.900 5.420 243.180 ;
  RECT 4.280 246.580 5.420 246.860 ;
  RECT 4.280 250.260 5.420 250.540 ;
  RECT 4.280 253.940 5.420 254.220 ;
  RECT 4.280 257.620 5.420 257.900 ;
  RECT 4.280 261.300 5.420 261.580 ;
  RECT 4.280 264.980 5.420 265.260 ;
  RECT 4.280 268.660 5.420 268.940 ;
  RECT 4.280 272.340 5.420 272.620 ;
  RECT 4.280 276.020 5.420 276.300 ;
  RECT 4.280 279.700 5.420 279.980 ;
  RECT 4.280 283.380 5.420 283.660 ;
  RECT 4.280 287.060 5.420 287.340 ;
  RECT 4.280 290.740 5.420 291.020 ;
  RECT 4.280 294.420 5.420 294.700 ;
  RECT 4.280 298.100 5.420 298.380 ;
  RECT 4.280 301.780 5.420 302.060 ;
  RECT 4.280 305.460 5.420 305.740 ;
  RECT 4.280 309.140 5.420 309.420 ;
  RECT 4.280 312.820 5.420 313.100 ;
  RECT 4.280 316.500 5.420 316.780 ;
  RECT 4.280 320.180 5.420 320.460 ;
  RECT 4.280 323.860 5.420 324.140 ;
  RECT 4.280 327.540 5.420 327.820 ;
  RECT 4.280 331.220 5.420 331.500 ;
  RECT 4.280 334.900 5.420 335.180 ;
  RECT 4.280 338.580 5.420 338.860 ;
  RECT 4.280 342.260 5.420 342.540 ;
  RECT 4.280 345.940 5.420 346.220 ;
  RECT 4.280 349.620 5.420 349.900 ;
  RECT 4.280 353.300 5.420 353.580 ;
  RECT 4.280 356.980 5.420 357.260 ;
  RECT 4.280 360.660 5.420 360.940 ;
  RECT 4.280 364.340 5.420 364.620 ;
  RECT 4.280 368.020 5.420 368.300 ;
  RECT 4.280 371.700 5.420 371.980 ;
  RECT 4.280 375.380 5.420 375.660 ;
  RECT 4.280 379.060 5.420 379.340 ;
  RECT 4.280 382.740 5.420 383.020 ;
  RECT 4.280 386.420 5.420 386.700 ;
  RECT 4.280 390.100 5.420 390.380 ;
  RECT 4.280 393.780 5.420 394.060 ;
  RECT 4.280 397.460 5.420 397.740 ;
  RECT 4.280 401.140 5.420 401.420 ;
  RECT 4.280 404.820 5.420 405.100 ;
  RECT 4.280 408.500 5.420 408.780 ;
  RECT 4.280 412.180 5.420 412.460 ;
  RECT 4.280 415.860 5.420 416.140 ;
  RECT 4.280 419.540 5.420 419.820 ;
  RECT 4.280 423.220 5.420 423.500 ;
  RECT 4.280 426.900 5.420 427.180 ;
  RECT 4.280 430.580 5.420 430.860 ;
  RECT 4.280 434.260 5.420 434.540 ;
  RECT 4.280 437.940 5.420 438.220 ;
  RECT 4.280 441.620 5.420 441.900 ;
  RECT 4.280 445.300 5.420 445.580 ;
  RECT 4.280 448.980 5.420 449.260 ;
  RECT 4.280 452.660 5.420 452.940 ;
  RECT 4.280 456.340 5.420 456.620 ;
  RECT 4.280 460.020 5.420 460.300 ;
  RECT 4.280 463.700 5.420 463.980 ;
  RECT 4.280 467.380 5.420 467.660 ;
  RECT 4.280 471.060 5.420 471.340 ;
  RECT 4.280 474.740 5.420 475.020 ;
  RECT 4.280 478.420 5.420 478.700 ;
  RECT 4.280 482.100 5.420 482.380 ;
  RECT 4.280 485.780 5.420 486.060 ;
  RECT 4.280 489.460 5.420 489.740 ;
  RECT 4.280 493.140 5.420 493.420 ;
  RECT 4.280 496.820 5.420 497.100 ;
  RECT 4.280 500.500 5.420 500.780 ;
  RECT 4.280 504.180 5.420 504.460 ;
  RECT 4.280 507.860 5.420 508.140 ;
  RECT 4.280 511.540 5.420 511.820 ;
  RECT 4.280 515.220 5.420 515.500 ;
  RECT 4.280 518.900 5.420 519.180 ;
  RECT 4.280 522.580 5.420 522.860 ;
  RECT 4.280 526.260 5.420 526.540 ;
  RECT 4.280 529.940 5.420 530.220 ;
  RECT 4.280 533.620 5.420 533.900 ;
  RECT 4.280 537.300 5.420 537.580 ;
  RECT 4.280 545.220 5.420 545.600 ;
  RECT 47.350 545.790 47.600 546.930 ;
  RECT 88.270 545.790 88.520 546.930 ;
  RECT 129.190 545.790 129.440 546.930 ;
  RECT 170.110 545.790 170.360 546.930 ;
  RECT 211.030 545.790 211.280 546.930 ;
  RECT 251.950 545.790 252.200 546.930 ;
  RECT 292.870 545.790 293.120 546.930 ;
  RECT 333.790 545.790 334.040 546.930 ;
  RECT 374.710 545.790 374.960 546.930 ;
  RECT 415.630 545.790 415.880 546.930 ;
  RECT 456.550 545.790 456.800 546.930 ;
  RECT 497.470 545.790 497.720 546.930 ;
  RECT 538.390 545.790 538.640 546.930 ;
  RECT 579.310 545.790 579.560 546.930 ;
  RECT 620.230 545.790 620.480 546.930 ;
  LAYER ME1 ;
  RECT 5.420 7.020 1374.080 545.790 ;
  RECT 1377.640 3.460 1379.500 549.350 ;
  RECT 0.000 3.460 1.860 549.350 ;
  RECT 1.860 549.350 1377.640 551.210 ;
  RECT 1.860 1.600 1377.640 3.460 ;
  RECT 1375.500 5.600 1377.360 547.210 ;
  RECT 2.140 5.600 4.000 547.210 ;
  RECT 4.000 547.210 1375.500 549.070 ;
  RECT 4.000 3.740 1375.500 5.600 ;
  RECT 2.140 547.210 4.000 549.070 ;
  RECT 0.000 549.350 1.860 551.210 ;
  RECT 1375.500 3.740 1377.360 5.600 ;
  RECT 1377.640 1.600 1379.500 3.460 ;
  RECT 1375.500 547.210 1377.360 549.070 ;
  RECT 1377.640 549.350 1379.500 551.210 ;
  RECT 2.140 3.740 4.000 5.600 ;
  RECT 0.000 1.600 1.860 3.460 ;
  RECT 1367.600 0.000 1368.400 1.000 ;
  RECT 1352.800 0.000 1353.600 1.000 ;
  RECT 1347.600 0.000 1348.400 1.000 ;
  RECT 1333.200 0.000 1334.000 1.000 ;
  RECT 1326.800 0.000 1327.600 1.000 ;
  RECT 1312.000 0.000 1312.800 1.000 ;
  RECT 1306.800 0.000 1307.600 1.000 ;
  RECT 1292.000 0.000 1292.800 1.000 ;
  RECT 1285.600 0.000 1286.400 1.000 ;
  RECT 1271.200 0.000 1272.000 1.000 ;
  RECT 1266.000 0.000 1266.800 1.000 ;
  RECT 1251.200 0.000 1252.000 1.000 ;
  RECT 1244.800 0.000 1245.600 1.000 ;
  RECT 1230.000 0.000 1230.800 1.000 ;
  RECT 1224.800 0.000 1225.600 1.000 ;
  RECT 1212.000 0.000 1212.800 1.000 ;
  RECT 1210.400 0.000 1211.200 1.000 ;
  RECT 1204.000 0.000 1204.800 1.000 ;
  RECT 1189.200 0.000 1190.000 1.000 ;
  RECT 1184.000 0.000 1184.800 1.000 ;
  RECT 1169.200 0.000 1170.000 1.000 ;
  RECT 1162.800 0.000 1163.600 1.000 ;
  RECT 1148.400 0.000 1149.200 1.000 ;
  RECT 1143.200 0.000 1144.000 1.000 ;
  RECT 1128.400 0.000 1129.200 1.000 ;
  RECT 1122.000 0.000 1122.800 1.000 ;
  RECT 1107.200 0.000 1108.000 1.000 ;
  RECT 1102.000 0.000 1102.800 1.000 ;
  RECT 1087.600 0.000 1088.400 1.000 ;
  RECT 1081.200 0.000 1082.000 1.000 ;
  RECT 1066.400 0.000 1067.200 1.000 ;
  RECT 1061.200 0.000 1062.000 1.000 ;
  RECT 1048.400 0.000 1049.200 1.000 ;
  RECT 1046.800 0.000 1047.600 1.000 ;
  RECT 1040.000 0.000 1040.800 1.000 ;
  RECT 1025.600 0.000 1026.400 1.000 ;
  RECT 1020.400 0.000 1021.200 1.000 ;
  RECT 1005.600 0.000 1006.400 1.000 ;
  RECT 999.200 0.000 1000.000 1.000 ;
  RECT 984.800 0.000 985.600 1.000 ;
  RECT 979.600 0.000 980.400 1.000 ;
  RECT 964.800 0.000 965.600 1.000 ;
  RECT 958.400 0.000 959.200 1.000 ;
  RECT 943.600 0.000 944.400 1.000 ;
  RECT 938.400 0.000 939.200 1.000 ;
  RECT 924.000 0.000 924.800 1.000 ;
  RECT 917.600 0.000 918.400 1.000 ;
  RECT 902.800 0.000 903.600 1.000 ;
  RECT 897.600 0.000 898.400 1.000 ;
  RECT 884.800 0.000 885.600 1.000 ;
  RECT 882.800 0.000 883.600 1.000 ;
  RECT 876.400 0.000 877.200 1.000 ;
  RECT 862.000 0.000 862.800 1.000 ;
  RECT 856.800 0.000 857.600 1.000 ;
  RECT 842.000 0.000 842.800 1.000 ;
  RECT 835.600 0.000 836.400 1.000 ;
  RECT 820.800 0.000 821.600 1.000 ;
  RECT 815.600 0.000 816.400 1.000 ;
  RECT 801.200 0.000 802.000 1.000 ;
  RECT 794.800 0.000 795.600 1.000 ;
  RECT 780.000 0.000 780.800 1.000 ;
  RECT 774.800 0.000 775.600 1.000 ;
  RECT 760.000 0.000 760.800 1.000 ;
  RECT 753.600 0.000 754.400 1.000 ;
  RECT 739.200 0.000 740.000 1.000 ;
  RECT 734.000 0.000 734.800 1.000 ;
  RECT 720.800 0.000 721.600 1.000 ;
  RECT 719.200 0.000 720.000 1.000 ;
  RECT 698.400 0.000 699.200 1.000 ;
  RECT 697.200 0.000 698.000 1.000 ;
  RECT 696.000 0.000 696.800 1.000 ;
  RECT 694.800 0.000 695.600 1.000 ;
  RECT 693.600 0.000 694.400 1.000 ;
  RECT 692.400 0.000 693.200 1.000 ;
  RECT 686.400 0.000 687.200 1.000 ;
  RECT 679.200 0.000 680.000 1.000 ;
  RECT 676.800 0.000 677.600 1.000 ;
  RECT 674.000 0.000 674.800 1.000 ;
  RECT 671.200 0.000 672.000 1.000 ;
  RECT 670.000 0.000 670.800 1.000 ;
  RECT 667.200 0.000 668.000 1.000 ;
  RECT 666.000 0.000 666.800 1.000 ;
  RECT 663.200 0.000 664.000 1.000 ;
  RECT 656.400 0.000 657.200 1.000 ;
  RECT 642.000 0.000 642.800 1.000 ;
  RECT 636.400 0.000 637.200 1.000 ;
  RECT 622.000 0.000 622.800 1.000 ;
  RECT 615.600 0.000 616.400 1.000 ;
  RECT 600.800 0.000 601.600 1.000 ;
  RECT 595.600 0.000 596.400 1.000 ;
  RECT 581.200 0.000 582.000 1.000 ;
  RECT 574.400 0.000 575.200 1.000 ;
  RECT 560.000 0.000 560.800 1.000 ;
  RECT 554.800 0.000 555.600 1.000 ;
  RECT 540.000 0.000 540.800 1.000 ;
  RECT 533.600 0.000 534.400 1.000 ;
  RECT 519.200 0.000 520.000 1.000 ;
  RECT 514.000 0.000 514.800 1.000 ;
  RECT 500.800 0.000 501.600 1.000 ;
  RECT 499.200 0.000 500.000 1.000 ;
  RECT 492.800 0.000 493.600 1.000 ;
  RECT 478.000 0.000 478.800 1.000 ;
  RECT 472.800 0.000 473.600 1.000 ;
  RECT 458.400 0.000 459.200 1.000 ;
  RECT 452.000 0.000 452.800 1.000 ;
  RECT 437.200 0.000 438.000 1.000 ;
  RECT 432.000 0.000 432.800 1.000 ;
  RECT 417.200 0.000 418.000 1.000 ;
  RECT 410.800 0.000 411.600 1.000 ;
  RECT 396.400 0.000 397.200 1.000 ;
  RECT 391.200 0.000 392.000 1.000 ;
  RECT 376.400 0.000 377.200 1.000 ;
  RECT 370.000 0.000 370.800 1.000 ;
  RECT 355.200 0.000 356.000 1.000 ;
  RECT 350.000 0.000 350.800 1.000 ;
  RECT 337.200 0.000 338.000 1.000 ;
  RECT 335.600 0.000 336.400 1.000 ;
  RECT 329.200 0.000 330.000 1.000 ;
  RECT 314.400 0.000 315.200 1.000 ;
  RECT 309.200 0.000 310.000 1.000 ;
  RECT 294.800 0.000 295.600 1.000 ;
  RECT 288.000 0.000 288.800 1.000 ;
  RECT 273.600 0.000 274.400 1.000 ;
  RECT 268.400 0.000 269.200 1.000 ;
  RECT 253.600 0.000 254.400 1.000 ;
  RECT 247.200 0.000 248.000 1.000 ;
  RECT 232.800 0.000 233.600 1.000 ;
  RECT 227.200 0.000 228.000 1.000 ;
  RECT 212.800 0.000 213.600 1.000 ;
  RECT 206.400 0.000 207.200 1.000 ;
  RECT 191.600 0.000 192.400 1.000 ;
  RECT 186.400 0.000 187.200 1.000 ;
  RECT 173.600 0.000 174.400 1.000 ;
  RECT 172.000 0.000 172.800 1.000 ;
  RECT 165.200 0.000 166.000 1.000 ;
  RECT 150.800 0.000 151.600 1.000 ;
  RECT 145.600 0.000 146.400 1.000 ;
  RECT 130.800 0.000 131.600 1.000 ;
  RECT 124.400 0.000 125.200 1.000 ;
  RECT 110.000 0.000 110.800 1.000 ;
  RECT 104.800 0.000 105.600 1.000 ;
  RECT 90.000 0.000 90.800 1.000 ;
  RECT 83.600 0.000 84.400 1.000 ;
  RECT 68.800 0.000 69.600 1.000 ;
  RECT 63.600 0.000 64.400 1.000 ;
  RECT 49.200 0.000 50.000 1.000 ;
  RECT 42.800 0.000 43.600 1.000 ;
  RECT 28.000 0.000 28.800 1.000 ;
  RECT 22.800 0.000 23.600 1.000 ;
  RECT 10.000 0.000 10.800 1.000 ;
  RECT 8.000 0.000 8.800 1.000 ;
  LAYER VI2 ;
  RECT 1377.640 3.600 1379.500 549.210 ;
  LAYER VI1 ;
  RECT 1377.640 3.460 1379.500 549.350 ;
  LAYER VI2 ;
  RECT 0.000 3.600 1.860 549.210 ;
  LAYER VI1 ;
  RECT 0.000 3.460 1.860 549.350 ;
  LAYER VI2 ;
  RECT 2.000 549.350 1377.500 551.210 ;
  LAYER VI1 ;
  RECT 1.860 549.350 1377.640 551.210 ;
  LAYER VI2 ;
  RECT 1369.400 1.600 1377.500 3.460 ;
  LAYER VI2 ;
  RECT 1354.600 1.600 1366.840 3.460 ;
  LAYER VI2 ;
  RECT 1349.400 1.600 1352.210 3.460 ;
  LAYER VI2 ;
  RECT 1335.000 1.600 1347.000 3.460 ;
  LAYER VI2 ;
  RECT 1328.600 1.600 1332.370 3.460 ;
  LAYER VI2 ;
  RECT 1313.800 1.600 1325.920 3.460 ;
  LAYER VI2 ;
  RECT 1308.600 1.600 1311.290 3.460 ;
  LAYER VI2 ;
  RECT 1293.800 1.600 1306.080 3.460 ;
  LAYER VI2 ;
  RECT 1287.400 1.600 1291.450 3.460 ;
  LAYER VI2 ;
  RECT 1273.000 1.600 1285.000 3.460 ;
  LAYER VI2 ;
  RECT 1267.800 1.600 1270.370 3.460 ;
  LAYER VI2 ;
  RECT 1253.000 1.600 1265.160 3.460 ;
  LAYER VI2 ;
  RECT 1246.600 1.600 1250.530 3.460 ;
  LAYER VI2 ;
  RECT 1231.800 1.600 1244.080 3.460 ;
  LAYER VI2 ;
  RECT 1226.600 1.600 1229.450 3.460 ;
  LAYER VI2 ;
  RECT 1213.800 1.600 1224.240 3.460 ;
  LAYER VI2 ;
  RECT 1205.800 1.600 1209.610 3.460 ;
  LAYER VI2 ;
  RECT 1191.000 1.600 1203.160 3.460 ;
  LAYER VI2 ;
  RECT 1185.800 1.600 1188.530 3.460 ;
  LAYER VI2 ;
  RECT 1171.000 1.600 1183.320 3.460 ;
  LAYER VI2 ;
  RECT 1164.600 1.600 1168.690 3.460 ;
  LAYER VI2 ;
  RECT 1150.200 1.600 1162.240 3.460 ;
  LAYER VI2 ;
  RECT 1145.000 1.600 1147.610 3.460 ;
  LAYER VI2 ;
  RECT 1130.200 1.600 1142.400 3.460 ;
  LAYER VI2 ;
  RECT 1123.800 1.600 1127.770 3.460 ;
  LAYER VI2 ;
  RECT 1109.000 1.600 1121.320 3.460 ;
  LAYER VI2 ;
  RECT 1103.800 1.600 1106.690 3.460 ;
  LAYER VI2 ;
  RECT 1089.400 1.600 1101.480 3.460 ;
  LAYER VI2 ;
  RECT 1083.000 1.600 1086.850 3.460 ;
  LAYER VI2 ;
  RECT 1068.200 1.600 1080.400 3.460 ;
  LAYER VI2 ;
  RECT 1063.000 1.600 1065.770 3.460 ;
  LAYER VI2 ;
  RECT 1050.200 1.600 1060.560 3.460 ;
  LAYER VI2 ;
  RECT 1041.800 1.600 1045.930 3.460 ;
  LAYER VI2 ;
  RECT 1027.400 1.600 1039.480 3.460 ;
  LAYER VI2 ;
  RECT 1022.200 1.600 1024.850 3.460 ;
  LAYER VI2 ;
  RECT 1007.400 1.600 1019.640 3.460 ;
  LAYER VI2 ;
  RECT 1001.000 1.600 1005.010 3.460 ;
  LAYER VI2 ;
  RECT 986.600 1.600 998.560 3.460 ;
  LAYER VI2 ;
  RECT 981.400 1.600 983.930 3.460 ;
  LAYER VI2 ;
  RECT 966.600 1.600 978.720 3.460 ;
  LAYER VI2 ;
  RECT 960.200 1.600 964.090 3.460 ;
  LAYER VI2 ;
  RECT 945.400 1.600 957.640 3.460 ;
  LAYER VI2 ;
  RECT 940.200 1.600 943.010 3.460 ;
  LAYER VI2 ;
  RECT 925.800 1.600 937.800 3.460 ;
  LAYER VI2 ;
  RECT 919.400 1.600 923.170 3.460 ;
  LAYER VI2 ;
  RECT 904.600 1.600 916.720 3.460 ;
  LAYER VI2 ;
  RECT 899.400 1.600 902.090 3.460 ;
  LAYER VI2 ;
  RECT 886.600 1.600 896.880 3.460 ;
  LAYER VI2 ;
  RECT 878.200 1.600 882.250 3.460 ;
  LAYER VI2 ;
  RECT 863.800 1.600 875.800 3.460 ;
  LAYER VI2 ;
  RECT 858.600 1.600 861.170 3.460 ;
  LAYER VI2 ;
  RECT 843.800 1.600 855.960 3.460 ;
  LAYER VI2 ;
  RECT 837.400 1.600 841.330 3.460 ;
  LAYER VI2 ;
  RECT 822.600 1.600 834.880 3.460 ;
  LAYER VI2 ;
  RECT 817.400 1.600 820.250 3.460 ;
  LAYER VI2 ;
  RECT 803.000 1.600 815.040 3.460 ;
  LAYER VI2 ;
  RECT 796.600 1.600 800.410 3.460 ;
  LAYER VI2 ;
  RECT 781.800 1.600 793.960 3.460 ;
  LAYER VI2 ;
  RECT 776.600 1.600 779.330 3.460 ;
  LAYER VI2 ;
  RECT 761.800 1.600 774.120 3.460 ;
  LAYER VI2 ;
  RECT 755.400 1.600 759.490 3.460 ;
  LAYER VI2 ;
  RECT 741.000 1.600 753.040 3.460 ;
  LAYER VI2 ;
  RECT 735.800 1.600 738.410 3.460 ;
  LAYER VI2 ;
  RECT 722.600 1.600 733.200 3.460 ;
  LAYER VI2 ;
  RECT 700.200 1.600 718.570 3.460 ;
  LAYER VI2 ;
  RECT 688.200 1.600 691.730 3.460 ;
  LAYER VI2 ;
  RECT 681.000 1.600 685.760 3.460 ;
  LAYER VI2 ;
  RECT 658.200 1.600 662.640 3.460 ;
  LAYER VI2 ;
  RECT 643.800 1.600 655.740 3.460 ;
  LAYER VI2 ;
  RECT 638.200 1.600 641.110 3.460 ;
  LAYER VI2 ;
  RECT 623.800 1.600 635.900 3.460 ;
  LAYER VI2 ;
  RECT 617.400 1.600 621.270 3.460 ;
  LAYER VI2 ;
  RECT 602.600 1.600 614.820 3.460 ;
  LAYER VI2 ;
  RECT 597.400 1.600 600.190 3.460 ;
  LAYER VI2 ;
  RECT 583.000 1.600 594.980 3.460 ;
  LAYER VI2 ;
  RECT 576.200 1.600 580.350 3.460 ;
  LAYER VI2 ;
  RECT 561.800 1.600 573.900 3.460 ;
  LAYER VI2 ;
  RECT 556.600 1.600 559.270 3.460 ;
  LAYER VI2 ;
  RECT 541.800 1.600 554.060 3.460 ;
  LAYER VI2 ;
  RECT 535.400 1.600 539.430 3.460 ;
  LAYER VI2 ;
  RECT 521.000 1.600 532.980 3.460 ;
  LAYER VI2 ;
  RECT 515.800 1.600 518.350 3.460 ;
  LAYER VI2 ;
  RECT 502.600 1.600 513.140 3.460 ;
  LAYER VI2 ;
  RECT 494.600 1.600 498.510 3.460 ;
  LAYER VI2 ;
  RECT 479.800 1.600 492.060 3.460 ;
  LAYER VI2 ;
  RECT 474.600 1.600 477.430 3.460 ;
  LAYER VI2 ;
  RECT 460.200 1.600 472.220 3.460 ;
  LAYER VI2 ;
  RECT 453.800 1.600 457.590 3.460 ;
  LAYER VI2 ;
  RECT 439.000 1.600 451.140 3.460 ;
  LAYER VI2 ;
  RECT 433.800 1.600 436.510 3.460 ;
  LAYER VI2 ;
  RECT 419.000 1.600 431.300 3.460 ;
  LAYER VI2 ;
  RECT 412.600 1.600 416.670 3.460 ;
  LAYER VI2 ;
  RECT 398.200 1.600 410.220 3.460 ;
  LAYER VI2 ;
  RECT 393.000 1.600 395.590 3.460 ;
  LAYER VI2 ;
  RECT 378.200 1.600 390.380 3.460 ;
  LAYER VI2 ;
  RECT 371.800 1.600 375.750 3.460 ;
  LAYER VI2 ;
  RECT 357.000 1.600 369.300 3.460 ;
  LAYER VI2 ;
  RECT 351.800 1.600 354.670 3.460 ;
  LAYER VI2 ;
  RECT 339.000 1.600 349.460 3.460 ;
  LAYER VI2 ;
  RECT 331.000 1.600 334.830 3.460 ;
  LAYER VI2 ;
  RECT 316.200 1.600 328.380 3.460 ;
  LAYER VI2 ;
  RECT 311.000 1.600 313.750 3.460 ;
  LAYER VI2 ;
  RECT 296.600 1.600 308.540 3.460 ;
  LAYER VI2 ;
  RECT 289.800 1.600 293.910 3.460 ;
  LAYER VI2 ;
  RECT 275.400 1.600 287.460 3.460 ;
  LAYER VI2 ;
  RECT 270.200 1.600 272.830 3.460 ;
  LAYER VI2 ;
  RECT 255.400 1.600 267.620 3.460 ;
  LAYER VI2 ;
  RECT 249.000 1.600 252.990 3.460 ;
  LAYER VI2 ;
  RECT 234.600 1.600 246.540 3.460 ;
  LAYER VI2 ;
  RECT 229.000 1.600 231.910 3.460 ;
  LAYER VI2 ;
  RECT 214.600 1.600 226.700 3.460 ;
  LAYER VI2 ;
  RECT 208.200 1.600 212.070 3.460 ;
  LAYER VI2 ;
  RECT 193.400 1.600 205.620 3.460 ;
  LAYER VI2 ;
  RECT 188.200 1.600 190.990 3.460 ;
  LAYER VI2 ;
  RECT 175.400 1.600 185.780 3.460 ;
  LAYER VI2 ;
  RECT 167.000 1.600 171.150 3.460 ;
  LAYER VI2 ;
  RECT 152.600 1.600 164.700 3.460 ;
  LAYER VI2 ;
  RECT 147.400 1.600 150.070 3.460 ;
  LAYER VI2 ;
  RECT 132.600 1.600 144.860 3.460 ;
  LAYER VI2 ;
  RECT 126.200 1.600 130.230 3.460 ;
  LAYER VI2 ;
  RECT 111.800 1.600 123.780 3.460 ;
  LAYER VI2 ;
  RECT 106.600 1.600 109.150 3.460 ;
  LAYER VI2 ;
  RECT 91.800 1.600 103.940 3.460 ;
  LAYER VI2 ;
  RECT 85.400 1.600 89.310 3.460 ;
  LAYER VI2 ;
  RECT 70.600 1.600 82.860 3.460 ;
  LAYER VI2 ;
  RECT 65.400 1.600 68.230 3.460 ;
  LAYER VI2 ;
  RECT 51.000 1.600 63.020 3.460 ;
  LAYER VI2 ;
  RECT 44.600 1.600 48.390 3.460 ;
  LAYER VI2 ;
  RECT 29.800 1.600 41.940 3.460 ;
  LAYER VI2 ;
  RECT 24.600 1.600 27.310 3.460 ;
  LAYER VI2 ;
  RECT 11.800 1.600 22.100 3.460 ;
  LAYER VI2 ;
  RECT 2.000 1.600 7.470 3.460 ;
  LAYER VI1 ;
  RECT 1369.400 1.600 1377.640 3.460 ;
  LAYER VI1 ;
  RECT 1354.600 1.600 1366.840 3.460 ;
  LAYER VI1 ;
  RECT 1349.400 1.600 1352.210 3.460 ;
  LAYER VI1 ;
  RECT 1335.000 1.600 1347.000 3.460 ;
  LAYER VI1 ;
  RECT 1328.600 1.600 1332.370 3.460 ;
  LAYER VI1 ;
  RECT 1313.800 1.600 1325.920 3.460 ;
  LAYER VI1 ;
  RECT 1308.600 1.600 1311.290 3.460 ;
  LAYER VI1 ;
  RECT 1293.800 1.600 1306.080 3.460 ;
  LAYER VI1 ;
  RECT 1287.400 1.600 1291.450 3.460 ;
  LAYER VI1 ;
  RECT 1273.000 1.600 1285.000 3.460 ;
  LAYER VI1 ;
  RECT 1267.800 1.600 1270.370 3.460 ;
  LAYER VI1 ;
  RECT 1253.000 1.600 1265.160 3.460 ;
  LAYER VI1 ;
  RECT 1246.600 1.600 1250.530 3.460 ;
  LAYER VI1 ;
  RECT 1231.800 1.600 1244.080 3.460 ;
  LAYER VI1 ;
  RECT 1226.600 1.600 1229.450 3.460 ;
  LAYER VI1 ;
  RECT 1213.800 1.600 1224.240 3.460 ;
  LAYER VI1 ;
  RECT 1205.800 1.600 1209.610 3.460 ;
  LAYER VI1 ;
  RECT 1191.000 1.600 1203.160 3.460 ;
  LAYER VI1 ;
  RECT 1185.800 1.600 1188.530 3.460 ;
  LAYER VI1 ;
  RECT 1171.000 1.600 1183.320 3.460 ;
  LAYER VI1 ;
  RECT 1164.600 1.600 1168.690 3.460 ;
  LAYER VI1 ;
  RECT 1150.200 1.600 1162.240 3.460 ;
  LAYER VI1 ;
  RECT 1145.000 1.600 1147.610 3.460 ;
  LAYER VI1 ;
  RECT 1130.200 1.600 1142.400 3.460 ;
  LAYER VI1 ;
  RECT 1123.800 1.600 1127.770 3.460 ;
  LAYER VI1 ;
  RECT 1109.000 1.600 1121.320 3.460 ;
  LAYER VI1 ;
  RECT 1103.800 1.600 1106.690 3.460 ;
  LAYER VI1 ;
  RECT 1089.400 1.600 1101.480 3.460 ;
  LAYER VI1 ;
  RECT 1083.000 1.600 1086.850 3.460 ;
  LAYER VI1 ;
  RECT 1068.200 1.600 1080.400 3.460 ;
  LAYER VI1 ;
  RECT 1063.000 1.600 1065.770 3.460 ;
  LAYER VI1 ;
  RECT 1050.200 1.600 1060.560 3.460 ;
  LAYER VI1 ;
  RECT 1041.800 1.600 1045.930 3.460 ;
  LAYER VI1 ;
  RECT 1027.400 1.600 1039.480 3.460 ;
  LAYER VI1 ;
  RECT 1022.200 1.600 1024.850 3.460 ;
  LAYER VI1 ;
  RECT 1007.400 1.600 1019.640 3.460 ;
  LAYER VI1 ;
  RECT 1001.000 1.600 1005.010 3.460 ;
  LAYER VI1 ;
  RECT 986.600 1.600 998.560 3.460 ;
  LAYER VI1 ;
  RECT 981.400 1.600 983.930 3.460 ;
  LAYER VI1 ;
  RECT 966.600 1.600 978.720 3.460 ;
  LAYER VI1 ;
  RECT 960.200 1.600 964.090 3.460 ;
  LAYER VI1 ;
  RECT 945.400 1.600 957.640 3.460 ;
  LAYER VI1 ;
  RECT 940.200 1.600 943.010 3.460 ;
  LAYER VI1 ;
  RECT 925.800 1.600 937.800 3.460 ;
  LAYER VI1 ;
  RECT 919.400 1.600 923.170 3.460 ;
  LAYER VI1 ;
  RECT 904.600 1.600 916.720 3.460 ;
  LAYER VI1 ;
  RECT 899.400 1.600 902.090 3.460 ;
  LAYER VI1 ;
  RECT 886.600 1.600 896.880 3.460 ;
  LAYER VI1 ;
  RECT 878.200 1.600 882.250 3.460 ;
  LAYER VI1 ;
  RECT 863.800 1.600 875.800 3.460 ;
  LAYER VI1 ;
  RECT 858.600 1.600 861.170 3.460 ;
  LAYER VI1 ;
  RECT 843.800 1.600 855.960 3.460 ;
  LAYER VI1 ;
  RECT 837.400 1.600 841.330 3.460 ;
  LAYER VI1 ;
  RECT 822.600 1.600 834.880 3.460 ;
  LAYER VI1 ;
  RECT 817.400 1.600 820.250 3.460 ;
  LAYER VI1 ;
  RECT 803.000 1.600 815.040 3.460 ;
  LAYER VI1 ;
  RECT 796.600 1.600 800.410 3.460 ;
  LAYER VI1 ;
  RECT 781.800 1.600 793.960 3.460 ;
  LAYER VI1 ;
  RECT 776.600 1.600 779.330 3.460 ;
  LAYER VI1 ;
  RECT 761.800 1.600 774.120 3.460 ;
  LAYER VI1 ;
  RECT 755.400 1.600 759.490 3.460 ;
  LAYER VI1 ;
  RECT 741.000 1.600 753.040 3.460 ;
  LAYER VI1 ;
  RECT 735.800 1.600 738.410 3.460 ;
  LAYER VI1 ;
  RECT 722.600 1.600 733.200 3.460 ;
  LAYER VI1 ;
  RECT 700.200 1.600 718.570 3.460 ;
  LAYER VI1 ;
  RECT 688.200 1.600 691.730 3.460 ;
  LAYER VI1 ;
  RECT 681.000 1.600 685.760 3.460 ;
  LAYER VI1 ;
  RECT 658.200 1.600 662.640 3.460 ;
  LAYER VI1 ;
  RECT 643.800 1.600 655.740 3.460 ;
  LAYER VI1 ;
  RECT 638.200 1.600 641.110 3.460 ;
  LAYER VI1 ;
  RECT 623.800 1.600 635.900 3.460 ;
  LAYER VI1 ;
  RECT 617.400 1.600 621.270 3.460 ;
  LAYER VI1 ;
  RECT 602.600 1.600 614.820 3.460 ;
  LAYER VI1 ;
  RECT 597.400 1.600 600.190 3.460 ;
  LAYER VI1 ;
  RECT 583.000 1.600 594.980 3.460 ;
  LAYER VI1 ;
  RECT 576.200 1.600 580.350 3.460 ;
  LAYER VI1 ;
  RECT 561.800 1.600 573.900 3.460 ;
  LAYER VI1 ;
  RECT 556.600 1.600 559.270 3.460 ;
  LAYER VI1 ;
  RECT 541.800 1.600 554.060 3.460 ;
  LAYER VI1 ;
  RECT 535.400 1.600 539.430 3.460 ;
  LAYER VI1 ;
  RECT 521.000 1.600 532.980 3.460 ;
  LAYER VI1 ;
  RECT 515.800 1.600 518.350 3.460 ;
  LAYER VI1 ;
  RECT 502.600 1.600 513.140 3.460 ;
  LAYER VI1 ;
  RECT 494.600 1.600 498.510 3.460 ;
  LAYER VI1 ;
  RECT 479.800 1.600 492.060 3.460 ;
  LAYER VI1 ;
  RECT 474.600 1.600 477.430 3.460 ;
  LAYER VI1 ;
  RECT 460.200 1.600 472.220 3.460 ;
  LAYER VI1 ;
  RECT 453.800 1.600 457.590 3.460 ;
  LAYER VI1 ;
  RECT 439.000 1.600 451.140 3.460 ;
  LAYER VI1 ;
  RECT 433.800 1.600 436.510 3.460 ;
  LAYER VI1 ;
  RECT 419.000 1.600 431.300 3.460 ;
  LAYER VI1 ;
  RECT 412.600 1.600 416.670 3.460 ;
  LAYER VI1 ;
  RECT 398.200 1.600 410.220 3.460 ;
  LAYER VI1 ;
  RECT 393.000 1.600 395.590 3.460 ;
  LAYER VI1 ;
  RECT 378.200 1.600 390.380 3.460 ;
  LAYER VI1 ;
  RECT 371.800 1.600 375.750 3.460 ;
  LAYER VI1 ;
  RECT 357.000 1.600 369.300 3.460 ;
  LAYER VI1 ;
  RECT 351.800 1.600 354.670 3.460 ;
  LAYER VI1 ;
  RECT 339.000 1.600 349.460 3.460 ;
  LAYER VI1 ;
  RECT 331.000 1.600 334.830 3.460 ;
  LAYER VI1 ;
  RECT 316.200 1.600 328.380 3.460 ;
  LAYER VI1 ;
  RECT 311.000 1.600 313.750 3.460 ;
  LAYER VI1 ;
  RECT 296.600 1.600 308.540 3.460 ;
  LAYER VI1 ;
  RECT 289.800 1.600 293.910 3.460 ;
  LAYER VI1 ;
  RECT 275.400 1.600 287.460 3.460 ;
  LAYER VI1 ;
  RECT 270.200 1.600 272.830 3.460 ;
  LAYER VI1 ;
  RECT 255.400 1.600 267.620 3.460 ;
  LAYER VI1 ;
  RECT 249.000 1.600 252.990 3.460 ;
  LAYER VI1 ;
  RECT 234.600 1.600 246.540 3.460 ;
  LAYER VI1 ;
  RECT 229.000 1.600 231.910 3.460 ;
  LAYER VI1 ;
  RECT 214.600 1.600 226.700 3.460 ;
  LAYER VI1 ;
  RECT 208.200 1.600 212.070 3.460 ;
  LAYER VI1 ;
  RECT 193.400 1.600 205.620 3.460 ;
  LAYER VI1 ;
  RECT 188.200 1.600 190.990 3.460 ;
  LAYER VI1 ;
  RECT 175.400 1.600 185.780 3.460 ;
  LAYER VI1 ;
  RECT 167.000 1.600 171.150 3.460 ;
  LAYER VI1 ;
  RECT 152.600 1.600 164.700 3.460 ;
  LAYER VI1 ;
  RECT 147.400 1.600 150.070 3.460 ;
  LAYER VI1 ;
  RECT 132.600 1.600 144.860 3.460 ;
  LAYER VI1 ;
  RECT 126.200 1.600 130.230 3.460 ;
  LAYER VI1 ;
  RECT 111.800 1.600 123.780 3.460 ;
  LAYER VI1 ;
  RECT 106.600 1.600 109.150 3.460 ;
  LAYER VI1 ;
  RECT 91.800 1.600 103.940 3.460 ;
  LAYER VI1 ;
  RECT 85.400 1.600 89.310 3.460 ;
  LAYER VI1 ;
  RECT 70.600 1.600 82.860 3.460 ;
  LAYER VI1 ;
  RECT 65.400 1.600 68.230 3.460 ;
  LAYER VI1 ;
  RECT 51.000 1.600 63.020 3.460 ;
  LAYER VI1 ;
  RECT 44.600 1.600 48.390 3.460 ;
  LAYER VI1 ;
  RECT 29.800 1.600 41.940 3.460 ;
  LAYER VI1 ;
  RECT 24.600 1.600 27.310 3.460 ;
  LAYER VI1 ;
  RECT 11.800 1.600 22.100 3.460 ;
  LAYER VI1 ;
  RECT 1.860 1.600 7.470 3.460 ;
  LAYER VI3 ;
  RECT 1375.500 540.280 1377.220 547.210 ;
  LAYER VI3 ;
  RECT 1375.500 64.930 1377.220 67.240 ;
  LAYER VI3 ;
  RECT 1375.500 44.080 1377.220 61.260 ;
  LAYER VI3 ;
  RECT 1375.500 39.620 1377.220 41.480 ;
  LAYER VI3 ;
  RECT 1375.500 29.870 1377.220 33.520 ;
  LAYER VI3 ;
  RECT 1375.500 24.270 1377.220 26.870 ;
  LAYER VI3 ;
  RECT 1375.500 18.130 1377.220 21.270 ;
  LAYER VI3 ;
  RECT 1375.500 5.600 1377.220 11.230 ;
  LAYER VI2 ;
  RECT 1375.500 540.280 1377.220 547.210 ;
  LAYER VI2 ;
  RECT 1375.500 64.930 1377.220 67.240 ;
  LAYER VI2 ;
  RECT 1375.500 44.080 1377.220 61.260 ;
  LAYER VI2 ;
  RECT 1375.500 39.620 1377.220 41.480 ;
  LAYER VI2 ;
  RECT 1375.500 29.870 1377.220 33.520 ;
  LAYER VI2 ;
  RECT 1375.500 24.270 1377.220 26.870 ;
  LAYER VI2 ;
  RECT 1375.500 18.130 1377.220 21.270 ;
  LAYER VI2 ;
  RECT 1375.500 5.600 1377.220 11.230 ;
  LAYER VI1 ;
  RECT 1375.500 5.600 1377.360 547.210 ;
  LAYER VI3 ;
  RECT 2.280 540.280 4.000 547.210 ;
  LAYER VI3 ;
  RECT 2.280 64.930 4.000 67.240 ;
  LAYER VI3 ;
  RECT 2.280 44.080 4.000 61.260 ;
  LAYER VI3 ;
  RECT 2.280 39.620 4.000 41.480 ;
  LAYER VI3 ;
  RECT 2.280 29.870 4.000 33.520 ;
  LAYER VI3 ;
  RECT 2.280 24.270 4.000 26.870 ;
  LAYER VI3 ;
  RECT 2.280 18.130 4.000 21.270 ;
  LAYER VI3 ;
  RECT 2.280 5.600 4.000 11.230 ;
  LAYER VI2 ;
  RECT 2.280 540.280 4.000 547.210 ;
  LAYER VI2 ;
  RECT 2.280 64.930 4.000 67.240 ;
  LAYER VI2 ;
  RECT 2.280 44.080 4.000 61.260 ;
  LAYER VI2 ;
  RECT 2.280 39.620 4.000 41.480 ;
  LAYER VI2 ;
  RECT 2.280 29.870 4.000 33.520 ;
  LAYER VI2 ;
  RECT 2.280 24.270 4.000 26.870 ;
  LAYER VI2 ;
  RECT 2.280 18.130 4.000 21.270 ;
  LAYER VI2 ;
  RECT 2.280 5.600 4.000 11.230 ;
  LAYER VI1 ;
  RECT 2.140 5.600 4.000 547.210 ;
  LAYER VI3 ;
  RECT 1332.580 547.210 1375.500 548.930 ;
  LAYER VI3 ;
  RECT 1291.660 547.210 1330.330 548.930 ;
  LAYER VI3 ;
  RECT 1250.740 547.210 1289.410 548.930 ;
  LAYER VI3 ;
  RECT 1209.820 547.210 1248.490 548.930 ;
  LAYER VI3 ;
  RECT 1168.900 547.210 1207.570 548.930 ;
  LAYER VI3 ;
  RECT 1127.980 547.210 1166.650 548.930 ;
  LAYER VI3 ;
  RECT 1087.060 547.210 1125.730 548.930 ;
  LAYER VI3 ;
  RECT 1046.140 547.210 1084.810 548.930 ;
  LAYER VI3 ;
  RECT 1005.220 547.210 1043.890 548.930 ;
  LAYER VI3 ;
  RECT 964.300 547.210 1002.970 548.930 ;
  LAYER VI3 ;
  RECT 923.380 547.210 962.050 548.930 ;
  LAYER VI3 ;
  RECT 882.460 547.210 921.130 548.930 ;
  LAYER VI3 ;
  RECT 841.540 547.210 880.210 548.930 ;
  LAYER VI3 ;
  RECT 800.620 547.210 839.290 548.930 ;
  LAYER VI3 ;
  RECT 759.700 547.210 798.370 548.930 ;
  LAYER VI3 ;
  RECT 718.780 547.210 757.450 548.930 ;
  LAYER VI3 ;
  RECT 700.040 547.210 713.040 548.930 ;
  LAYER VI3 ;
  RECT 688.910 547.210 693.720 548.930 ;
  LAYER VI3 ;
  RECT 679.200 547.210 683.720 548.930 ;
  LAYER VI3 ;
  RECT 673.860 547.210 675.440 548.930 ;
  LAYER VI3 ;
  RECT 622.050 547.210 661.080 548.930 ;
  LAYER VI3 ;
  RECT 581.130 547.210 619.800 548.930 ;
  LAYER VI3 ;
  RECT 540.210 547.210 578.880 548.930 ;
  LAYER VI3 ;
  RECT 499.290 547.210 537.960 548.930 ;
  LAYER VI3 ;
  RECT 458.370 547.210 497.040 548.930 ;
  LAYER VI3 ;
  RECT 417.450 547.210 456.120 548.930 ;
  LAYER VI3 ;
  RECT 376.530 547.210 415.200 548.930 ;
  LAYER VI3 ;
  RECT 335.610 547.210 374.280 548.930 ;
  LAYER VI3 ;
  RECT 294.690 547.210 333.360 548.930 ;
  LAYER VI3 ;
  RECT 253.770 547.210 292.440 548.930 ;
  LAYER VI3 ;
  RECT 212.850 547.210 251.520 548.930 ;
  LAYER VI3 ;
  RECT 171.930 547.210 210.600 548.930 ;
  LAYER VI3 ;
  RECT 131.010 547.210 169.680 548.930 ;
  LAYER VI3 ;
  RECT 90.090 547.210 128.760 548.930 ;
  LAYER VI3 ;
  RECT 49.170 547.210 87.840 548.930 ;
  LAYER VI3 ;
  RECT 4.000 547.210 46.920 548.930 ;
  LAYER VI2 ;
  RECT 1332.580 547.210 1375.500 548.930 ;
  LAYER VI2 ;
  RECT 1291.660 547.210 1330.330 548.930 ;
  LAYER VI2 ;
  RECT 1250.740 547.210 1289.410 548.930 ;
  LAYER VI2 ;
  RECT 1209.820 547.210 1248.490 548.930 ;
  LAYER VI2 ;
  RECT 1168.900 547.210 1207.570 548.930 ;
  LAYER VI2 ;
  RECT 1127.980 547.210 1166.650 548.930 ;
  LAYER VI2 ;
  RECT 1087.060 547.210 1125.730 548.930 ;
  LAYER VI2 ;
  RECT 1046.140 547.210 1084.810 548.930 ;
  LAYER VI2 ;
  RECT 1005.220 547.210 1043.890 548.930 ;
  LAYER VI2 ;
  RECT 964.300 547.210 1002.970 548.930 ;
  LAYER VI2 ;
  RECT 923.380 547.210 962.050 548.930 ;
  LAYER VI2 ;
  RECT 882.460 547.210 921.130 548.930 ;
  LAYER VI2 ;
  RECT 841.540 547.210 880.210 548.930 ;
  LAYER VI2 ;
  RECT 800.620 547.210 839.290 548.930 ;
  LAYER VI2 ;
  RECT 759.700 547.210 798.370 548.930 ;
  LAYER VI2 ;
  RECT 718.780 547.210 757.450 548.930 ;
  LAYER VI2 ;
  RECT 700.040 547.210 713.040 548.930 ;
  LAYER VI2 ;
  RECT 688.910 547.210 693.720 548.930 ;
  LAYER VI2 ;
  RECT 679.200 547.210 683.720 548.930 ;
  LAYER VI2 ;
  RECT 673.860 547.210 675.440 548.930 ;
  LAYER VI2 ;
  RECT 622.050 547.210 661.080 548.930 ;
  LAYER VI2 ;
  RECT 581.130 547.210 619.800 548.930 ;
  LAYER VI2 ;
  RECT 540.210 547.210 578.880 548.930 ;
  LAYER VI2 ;
  RECT 499.290 547.210 537.960 548.930 ;
  LAYER VI2 ;
  RECT 458.370 547.210 497.040 548.930 ;
  LAYER VI2 ;
  RECT 417.450 547.210 456.120 548.930 ;
  LAYER VI2 ;
  RECT 376.530 547.210 415.200 548.930 ;
  LAYER VI2 ;
  RECT 335.610 547.210 374.280 548.930 ;
  LAYER VI2 ;
  RECT 294.690 547.210 333.360 548.930 ;
  LAYER VI2 ;
  RECT 253.770 547.210 292.440 548.930 ;
  LAYER VI2 ;
  RECT 212.850 547.210 251.520 548.930 ;
  LAYER VI2 ;
  RECT 171.930 547.210 210.600 548.930 ;
  LAYER VI2 ;
  RECT 131.010 547.210 169.680 548.930 ;
  LAYER VI2 ;
  RECT 90.090 547.210 128.760 548.930 ;
  LAYER VI2 ;
  RECT 49.170 547.210 87.840 548.930 ;
  LAYER VI2 ;
  RECT 4.000 547.210 46.920 548.930 ;
  LAYER VI1 ;
  RECT 4.000 547.210 1375.500 549.070 ;
  LAYER VI3 ;
  RECT 1362.100 3.880 1371.940 5.600 ;
  LAYER VI3 ;
  RECT 1342.260 3.880 1352.100 5.600 ;
  LAYER VI3 ;
  RECT 1321.180 3.880 1332.260 5.600 ;
  LAYER VI3 ;
  RECT 1301.340 3.880 1311.180 5.600 ;
  LAYER VI3 ;
  RECT 1280.260 3.880 1291.340 5.600 ;
  LAYER VI3 ;
  RECT 1260.420 3.880 1270.260 5.600 ;
  LAYER VI3 ;
  RECT 1239.340 3.880 1250.420 5.600 ;
  LAYER VI3 ;
  RECT 1219.500 3.880 1229.340 5.600 ;
  LAYER VI3 ;
  RECT 1198.420 3.880 1209.500 5.600 ;
  LAYER VI3 ;
  RECT 1178.580 3.880 1188.420 5.600 ;
  LAYER VI3 ;
  RECT 1157.500 3.880 1168.580 5.600 ;
  LAYER VI3 ;
  RECT 1137.660 3.880 1147.500 5.600 ;
  LAYER VI3 ;
  RECT 1116.580 3.880 1127.660 5.600 ;
  LAYER VI3 ;
  RECT 1096.740 3.880 1106.580 5.600 ;
  LAYER VI3 ;
  RECT 1075.660 3.880 1086.740 5.600 ;
  LAYER VI3 ;
  RECT 1055.820 3.880 1065.660 5.600 ;
  LAYER VI3 ;
  RECT 1034.740 3.880 1045.820 5.600 ;
  LAYER VI3 ;
  RECT 1014.900 3.880 1024.740 5.600 ;
  LAYER VI3 ;
  RECT 993.820 3.880 1004.900 5.600 ;
  LAYER VI3 ;
  RECT 973.980 3.880 983.820 5.600 ;
  LAYER VI3 ;
  RECT 952.900 3.880 963.980 5.600 ;
  LAYER VI3 ;
  RECT 933.060 3.880 942.900 5.600 ;
  LAYER VI3 ;
  RECT 911.980 3.880 923.060 5.600 ;
  LAYER VI3 ;
  RECT 892.140 3.880 901.980 5.600 ;
  LAYER VI3 ;
  RECT 871.060 3.880 882.140 5.600 ;
  LAYER VI3 ;
  RECT 851.220 3.880 861.060 5.600 ;
  LAYER VI3 ;
  RECT 830.140 3.880 841.220 5.600 ;
  LAYER VI3 ;
  RECT 810.300 3.880 820.140 5.600 ;
  LAYER VI3 ;
  RECT 789.220 3.880 800.300 5.600 ;
  LAYER VI3 ;
  RECT 769.380 3.880 779.220 5.600 ;
  LAYER VI3 ;
  RECT 748.300 3.880 759.380 5.600 ;
  LAYER VI3 ;
  RECT 728.460 3.880 738.300 5.600 ;
  LAYER VI3 ;
  RECT 700.490 3.880 718.460 5.600 ;
  LAYER VI3 ;
  RECT 689.170 3.880 692.570 5.600 ;
  LAYER VI3 ;
  RECT 679.200 3.880 683.720 5.600 ;
  LAYER VI3 ;
  RECT 673.860 3.880 675.440 5.600 ;
  LAYER VI3 ;
  RECT 651.000 3.880 662.100 5.600 ;
  LAYER VI3 ;
  RECT 631.160 3.880 641.000 5.600 ;
  LAYER VI3 ;
  RECT 610.080 3.880 621.160 5.600 ;
  LAYER VI3 ;
  RECT 590.240 3.880 600.080 5.600 ;
  LAYER VI3 ;
  RECT 569.160 3.880 580.240 5.600 ;
  LAYER VI3 ;
  RECT 549.320 3.880 559.160 5.600 ;
  LAYER VI3 ;
  RECT 528.240 3.880 539.320 5.600 ;
  LAYER VI3 ;
  RECT 508.400 3.880 518.240 5.600 ;
  LAYER VI3 ;
  RECT 487.320 3.880 498.400 5.600 ;
  LAYER VI3 ;
  RECT 467.480 3.880 477.320 5.600 ;
  LAYER VI3 ;
  RECT 446.400 3.880 457.480 5.600 ;
  LAYER VI3 ;
  RECT 426.560 3.880 436.400 5.600 ;
  LAYER VI3 ;
  RECT 405.480 3.880 416.560 5.600 ;
  LAYER VI3 ;
  RECT 385.640 3.880 395.480 5.600 ;
  LAYER VI3 ;
  RECT 364.560 3.880 375.640 5.600 ;
  LAYER VI3 ;
  RECT 344.720 3.880 354.560 5.600 ;
  LAYER VI3 ;
  RECT 323.640 3.880 334.720 5.600 ;
  LAYER VI3 ;
  RECT 303.800 3.880 313.640 5.600 ;
  LAYER VI3 ;
  RECT 282.720 3.880 293.800 5.600 ;
  LAYER VI3 ;
  RECT 262.880 3.880 272.720 5.600 ;
  LAYER VI3 ;
  RECT 241.800 3.880 252.880 5.600 ;
  LAYER VI3 ;
  RECT 221.960 3.880 231.800 5.600 ;
  LAYER VI3 ;
  RECT 200.880 3.880 211.960 5.600 ;
  LAYER VI3 ;
  RECT 181.040 3.880 190.880 5.600 ;
  LAYER VI3 ;
  RECT 159.960 3.880 171.040 5.600 ;
  LAYER VI3 ;
  RECT 140.120 3.880 149.960 5.600 ;
  LAYER VI3 ;
  RECT 119.040 3.880 130.120 5.600 ;
  LAYER VI3 ;
  RECT 99.200 3.880 109.040 5.600 ;
  LAYER VI3 ;
  RECT 78.120 3.880 89.200 5.600 ;
  LAYER VI3 ;
  RECT 58.280 3.880 68.120 5.600 ;
  LAYER VI3 ;
  RECT 37.200 3.880 48.280 5.600 ;
  LAYER VI3 ;
  RECT 17.360 3.880 27.200 5.600 ;
  LAYER VI2 ;
  RECT 1369.400 3.880 1371.940 5.600 ;
  LAYER VI2 ;
  RECT 1362.100 3.880 1366.840 5.600 ;
  LAYER VI2 ;
  RECT 1349.400 3.880 1352.100 5.600 ;
  LAYER VI2 ;
  RECT 1342.260 3.880 1347.000 5.600 ;
  LAYER VI2 ;
  RECT 1328.600 3.880 1332.260 5.600 ;
  LAYER VI2 ;
  RECT 1321.180 3.880 1325.920 5.600 ;
  LAYER VI2 ;
  RECT 1308.600 3.880 1311.180 5.600 ;
  LAYER VI2 ;
  RECT 1301.340 3.880 1306.080 5.600 ;
  LAYER VI2 ;
  RECT 1287.400 3.880 1291.340 5.600 ;
  LAYER VI2 ;
  RECT 1280.260 3.880 1285.000 5.600 ;
  LAYER VI2 ;
  RECT 1267.800 3.880 1270.260 5.600 ;
  LAYER VI2 ;
  RECT 1260.420 3.880 1265.160 5.600 ;
  LAYER VI2 ;
  RECT 1246.600 3.880 1250.420 5.600 ;
  LAYER VI2 ;
  RECT 1239.340 3.880 1244.080 5.600 ;
  LAYER VI2 ;
  RECT 1226.600 3.880 1229.340 5.600 ;
  LAYER VI2 ;
  RECT 1219.500 3.880 1224.240 5.600 ;
  LAYER VI2 ;
  RECT 1205.800 3.880 1209.500 5.600 ;
  LAYER VI2 ;
  RECT 1198.420 3.880 1203.160 5.600 ;
  LAYER VI2 ;
  RECT 1185.800 3.880 1188.420 5.600 ;
  LAYER VI2 ;
  RECT 1178.580 3.880 1183.320 5.600 ;
  LAYER VI2 ;
  RECT 1164.600 3.880 1168.580 5.600 ;
  LAYER VI2 ;
  RECT 1157.500 3.880 1162.240 5.600 ;
  LAYER VI2 ;
  RECT 1145.000 3.880 1147.500 5.600 ;
  LAYER VI2 ;
  RECT 1137.660 3.880 1142.400 5.600 ;
  LAYER VI2 ;
  RECT 1123.800 3.880 1127.660 5.600 ;
  LAYER VI2 ;
  RECT 1116.580 3.880 1121.320 5.600 ;
  LAYER VI2 ;
  RECT 1103.800 3.880 1106.580 5.600 ;
  LAYER VI2 ;
  RECT 1096.740 3.880 1101.480 5.600 ;
  LAYER VI2 ;
  RECT 1083.000 3.880 1086.740 5.600 ;
  LAYER VI2 ;
  RECT 1075.660 3.880 1080.400 5.600 ;
  LAYER VI2 ;
  RECT 1063.000 3.880 1065.660 5.600 ;
  LAYER VI2 ;
  RECT 1055.820 3.880 1060.560 5.600 ;
  LAYER VI2 ;
  RECT 1041.800 3.880 1045.820 5.600 ;
  LAYER VI2 ;
  RECT 1034.740 3.880 1039.480 5.600 ;
  LAYER VI2 ;
  RECT 1022.200 3.880 1024.740 5.600 ;
  LAYER VI2 ;
  RECT 1014.900 3.880 1019.640 5.600 ;
  LAYER VI2 ;
  RECT 1001.000 3.880 1004.900 5.600 ;
  LAYER VI2 ;
  RECT 993.820 3.880 998.560 5.600 ;
  LAYER VI2 ;
  RECT 981.400 3.880 983.820 5.600 ;
  LAYER VI2 ;
  RECT 973.980 3.880 978.720 5.600 ;
  LAYER VI2 ;
  RECT 960.200 3.880 963.980 5.600 ;
  LAYER VI2 ;
  RECT 952.900 3.880 957.640 5.600 ;
  LAYER VI2 ;
  RECT 940.200 3.880 942.900 5.600 ;
  LAYER VI2 ;
  RECT 933.060 3.880 937.800 5.600 ;
  LAYER VI2 ;
  RECT 919.400 3.880 923.060 5.600 ;
  LAYER VI2 ;
  RECT 911.980 3.880 916.720 5.600 ;
  LAYER VI2 ;
  RECT 899.400 3.880 901.980 5.600 ;
  LAYER VI2 ;
  RECT 892.140 3.880 896.880 5.600 ;
  LAYER VI2 ;
  RECT 878.200 3.880 882.140 5.600 ;
  LAYER VI2 ;
  RECT 871.060 3.880 875.800 5.600 ;
  LAYER VI2 ;
  RECT 858.600 3.880 861.060 5.600 ;
  LAYER VI2 ;
  RECT 851.220 3.880 855.960 5.600 ;
  LAYER VI2 ;
  RECT 837.400 3.880 841.220 5.600 ;
  LAYER VI2 ;
  RECT 830.140 3.880 834.880 5.600 ;
  LAYER VI2 ;
  RECT 817.400 3.880 820.140 5.600 ;
  LAYER VI2 ;
  RECT 810.300 3.880 815.040 5.600 ;
  LAYER VI2 ;
  RECT 796.600 3.880 800.300 5.600 ;
  LAYER VI2 ;
  RECT 789.220 3.880 793.960 5.600 ;
  LAYER VI2 ;
  RECT 776.600 3.880 779.220 5.600 ;
  LAYER VI2 ;
  RECT 769.380 3.880 774.120 5.600 ;
  LAYER VI2 ;
  RECT 755.400 3.880 759.380 5.600 ;
  LAYER VI2 ;
  RECT 748.300 3.880 753.040 5.600 ;
  LAYER VI2 ;
  RECT 735.800 3.880 738.300 5.600 ;
  LAYER VI2 ;
  RECT 728.460 3.880 733.200 5.600 ;
  LAYER VI2 ;
  RECT 700.490 3.880 718.460 5.600 ;
  LAYER VI2 ;
  RECT 689.170 3.880 691.730 5.600 ;
  LAYER VI2 ;
  RECT 681.000 3.880 683.720 5.600 ;
  LAYER VI2 ;
  RECT 658.200 3.880 662.100 5.600 ;
  LAYER VI2 ;
  RECT 651.000 3.880 655.740 5.600 ;
  LAYER VI2 ;
  RECT 638.200 3.880 641.000 5.600 ;
  LAYER VI2 ;
  RECT 631.160 3.880 635.900 5.600 ;
  LAYER VI2 ;
  RECT 617.400 3.880 621.160 5.600 ;
  LAYER VI2 ;
  RECT 610.080 3.880 614.820 5.600 ;
  LAYER VI2 ;
  RECT 597.400 3.880 600.080 5.600 ;
  LAYER VI2 ;
  RECT 590.240 3.880 594.980 5.600 ;
  LAYER VI2 ;
  RECT 576.200 3.880 580.240 5.600 ;
  LAYER VI2 ;
  RECT 569.160 3.880 573.900 5.600 ;
  LAYER VI2 ;
  RECT 556.600 3.880 559.160 5.600 ;
  LAYER VI2 ;
  RECT 549.320 3.880 554.060 5.600 ;
  LAYER VI2 ;
  RECT 535.400 3.880 539.320 5.600 ;
  LAYER VI2 ;
  RECT 528.240 3.880 532.980 5.600 ;
  LAYER VI2 ;
  RECT 515.800 3.880 518.240 5.600 ;
  LAYER VI2 ;
  RECT 508.400 3.880 513.140 5.600 ;
  LAYER VI2 ;
  RECT 494.600 3.880 498.400 5.600 ;
  LAYER VI2 ;
  RECT 487.320 3.880 492.060 5.600 ;
  LAYER VI2 ;
  RECT 474.600 3.880 477.320 5.600 ;
  LAYER VI2 ;
  RECT 467.480 3.880 472.220 5.600 ;
  LAYER VI2 ;
  RECT 453.800 3.880 457.480 5.600 ;
  LAYER VI2 ;
  RECT 446.400 3.880 451.140 5.600 ;
  LAYER VI2 ;
  RECT 433.800 3.880 436.400 5.600 ;
  LAYER VI2 ;
  RECT 426.560 3.880 431.300 5.600 ;
  LAYER VI2 ;
  RECT 412.600 3.880 416.560 5.600 ;
  LAYER VI2 ;
  RECT 405.480 3.880 410.220 5.600 ;
  LAYER VI2 ;
  RECT 393.000 3.880 395.480 5.600 ;
  LAYER VI2 ;
  RECT 385.640 3.880 390.380 5.600 ;
  LAYER VI2 ;
  RECT 371.800 3.880 375.640 5.600 ;
  LAYER VI2 ;
  RECT 364.560 3.880 369.300 5.600 ;
  LAYER VI2 ;
  RECT 351.800 3.880 354.560 5.600 ;
  LAYER VI2 ;
  RECT 344.720 3.880 349.460 5.600 ;
  LAYER VI2 ;
  RECT 331.000 3.880 334.720 5.600 ;
  LAYER VI2 ;
  RECT 323.640 3.880 328.380 5.600 ;
  LAYER VI2 ;
  RECT 311.000 3.880 313.640 5.600 ;
  LAYER VI2 ;
  RECT 303.800 3.880 308.540 5.600 ;
  LAYER VI2 ;
  RECT 289.800 3.880 293.800 5.600 ;
  LAYER VI2 ;
  RECT 282.720 3.880 287.460 5.600 ;
  LAYER VI2 ;
  RECT 270.200 3.880 272.720 5.600 ;
  LAYER VI2 ;
  RECT 262.880 3.880 267.620 5.600 ;
  LAYER VI2 ;
  RECT 249.000 3.880 252.880 5.600 ;
  LAYER VI2 ;
  RECT 241.800 3.880 246.540 5.600 ;
  LAYER VI2 ;
  RECT 229.000 3.880 231.800 5.600 ;
  LAYER VI2 ;
  RECT 221.960 3.880 226.700 5.600 ;
  LAYER VI2 ;
  RECT 208.200 3.880 211.960 5.600 ;
  LAYER VI2 ;
  RECT 200.880 3.880 205.620 5.600 ;
  LAYER VI2 ;
  RECT 188.200 3.880 190.880 5.600 ;
  LAYER VI2 ;
  RECT 181.040 3.880 185.780 5.600 ;
  LAYER VI2 ;
  RECT 167.000 3.880 171.040 5.600 ;
  LAYER VI2 ;
  RECT 159.960 3.880 164.700 5.600 ;
  LAYER VI2 ;
  RECT 147.400 3.880 149.960 5.600 ;
  LAYER VI2 ;
  RECT 140.120 3.880 144.860 5.600 ;
  LAYER VI2 ;
  RECT 126.200 3.880 130.120 5.600 ;
  LAYER VI2 ;
  RECT 119.040 3.880 123.780 5.600 ;
  LAYER VI2 ;
  RECT 106.600 3.880 109.040 5.600 ;
  LAYER VI2 ;
  RECT 99.200 3.880 103.940 5.600 ;
  LAYER VI2 ;
  RECT 85.400 3.880 89.200 5.600 ;
  LAYER VI2 ;
  RECT 78.120 3.880 82.860 5.600 ;
  LAYER VI2 ;
  RECT 65.400 3.880 68.120 5.600 ;
  LAYER VI2 ;
  RECT 58.280 3.880 63.020 5.600 ;
  LAYER VI2 ;
  RECT 44.600 3.880 48.280 5.600 ;
  LAYER VI2 ;
  RECT 37.200 3.880 41.940 5.600 ;
  LAYER VI2 ;
  RECT 24.600 3.880 27.200 5.600 ;
  LAYER VI2 ;
  RECT 17.360 3.880 22.100 5.600 ;
  LAYER VI1 ;
  RECT 1369.400 3.740 1375.500 5.600 ;
  LAYER VI1 ;
  RECT 1354.600 3.740 1366.840 5.600 ;
  LAYER VI1 ;
  RECT 1349.400 3.740 1352.210 5.600 ;
  LAYER VI1 ;
  RECT 1335.000 3.740 1347.000 5.600 ;
  LAYER VI1 ;
  RECT 1328.600 3.740 1332.370 5.600 ;
  LAYER VI1 ;
  RECT 1313.800 3.740 1325.920 5.600 ;
  LAYER VI1 ;
  RECT 1308.600 3.740 1311.290 5.600 ;
  LAYER VI1 ;
  RECT 1293.800 3.740 1306.080 5.600 ;
  LAYER VI1 ;
  RECT 1287.400 3.740 1291.450 5.600 ;
  LAYER VI1 ;
  RECT 1273.000 3.740 1285.000 5.600 ;
  LAYER VI1 ;
  RECT 1267.800 3.740 1270.370 5.600 ;
  LAYER VI1 ;
  RECT 1253.000 3.740 1265.160 5.600 ;
  LAYER VI1 ;
  RECT 1246.600 3.740 1250.530 5.600 ;
  LAYER VI1 ;
  RECT 1231.800 3.740 1244.080 5.600 ;
  LAYER VI1 ;
  RECT 1226.600 3.740 1229.450 5.600 ;
  LAYER VI1 ;
  RECT 1213.800 3.740 1224.240 5.600 ;
  LAYER VI1 ;
  RECT 1205.800 3.740 1209.610 5.600 ;
  LAYER VI1 ;
  RECT 1191.000 3.740 1203.160 5.600 ;
  LAYER VI1 ;
  RECT 1185.800 3.740 1188.530 5.600 ;
  LAYER VI1 ;
  RECT 1171.000 3.740 1183.320 5.600 ;
  LAYER VI1 ;
  RECT 1164.600 3.740 1168.690 5.600 ;
  LAYER VI1 ;
  RECT 1150.200 3.740 1162.240 5.600 ;
  LAYER VI1 ;
  RECT 1145.000 3.740 1147.610 5.600 ;
  LAYER VI1 ;
  RECT 1130.200 3.740 1142.400 5.600 ;
  LAYER VI1 ;
  RECT 1123.800 3.740 1127.770 5.600 ;
  LAYER VI1 ;
  RECT 1109.000 3.740 1121.320 5.600 ;
  LAYER VI1 ;
  RECT 1103.800 3.740 1106.690 5.600 ;
  LAYER VI1 ;
  RECT 1089.400 3.740 1101.480 5.600 ;
  LAYER VI1 ;
  RECT 1083.000 3.740 1086.850 5.600 ;
  LAYER VI1 ;
  RECT 1068.200 3.740 1080.400 5.600 ;
  LAYER VI1 ;
  RECT 1063.000 3.740 1065.770 5.600 ;
  LAYER VI1 ;
  RECT 1050.200 3.740 1060.560 5.600 ;
  LAYER VI1 ;
  RECT 1041.800 3.740 1045.930 5.600 ;
  LAYER VI1 ;
  RECT 1027.400 3.740 1039.480 5.600 ;
  LAYER VI1 ;
  RECT 1022.200 3.740 1024.850 5.600 ;
  LAYER VI1 ;
  RECT 1007.400 3.740 1019.640 5.600 ;
  LAYER VI1 ;
  RECT 1001.000 3.740 1005.010 5.600 ;
  LAYER VI1 ;
  RECT 986.600 3.740 998.560 5.600 ;
  LAYER VI1 ;
  RECT 981.400 3.740 983.930 5.600 ;
  LAYER VI1 ;
  RECT 966.600 3.740 978.720 5.600 ;
  LAYER VI1 ;
  RECT 960.200 3.740 964.090 5.600 ;
  LAYER VI1 ;
  RECT 945.400 3.740 957.640 5.600 ;
  LAYER VI1 ;
  RECT 940.200 3.740 943.010 5.600 ;
  LAYER VI1 ;
  RECT 925.800 3.740 937.800 5.600 ;
  LAYER VI1 ;
  RECT 919.400 3.740 923.170 5.600 ;
  LAYER VI1 ;
  RECT 904.600 3.740 916.720 5.600 ;
  LAYER VI1 ;
  RECT 899.400 3.740 902.090 5.600 ;
  LAYER VI1 ;
  RECT 886.600 3.740 896.880 5.600 ;
  LAYER VI1 ;
  RECT 878.200 3.740 882.250 5.600 ;
  LAYER VI1 ;
  RECT 863.800 3.740 875.800 5.600 ;
  LAYER VI1 ;
  RECT 858.600 3.740 861.170 5.600 ;
  LAYER VI1 ;
  RECT 843.800 3.740 855.960 5.600 ;
  LAYER VI1 ;
  RECT 837.400 3.740 841.330 5.600 ;
  LAYER VI1 ;
  RECT 822.600 3.740 834.880 5.600 ;
  LAYER VI1 ;
  RECT 817.400 3.740 820.250 5.600 ;
  LAYER VI1 ;
  RECT 803.000 3.740 815.040 5.600 ;
  LAYER VI1 ;
  RECT 796.600 3.740 800.410 5.600 ;
  LAYER VI1 ;
  RECT 781.800 3.740 793.960 5.600 ;
  LAYER VI1 ;
  RECT 776.600 3.740 779.330 5.600 ;
  LAYER VI1 ;
  RECT 761.800 3.740 774.120 5.600 ;
  LAYER VI1 ;
  RECT 755.400 3.740 759.490 5.600 ;
  LAYER VI1 ;
  RECT 741.000 3.740 753.040 5.600 ;
  LAYER VI1 ;
  RECT 735.800 3.740 738.410 5.600 ;
  LAYER VI1 ;
  RECT 722.600 3.740 733.200 5.600 ;
  LAYER VI1 ;
  RECT 700.200 3.740 718.570 5.600 ;
  LAYER VI1 ;
  RECT 688.200 3.740 691.730 5.600 ;
  LAYER VI1 ;
  RECT 681.000 3.740 685.760 5.600 ;
  LAYER VI1 ;
  RECT 658.200 3.740 662.640 5.600 ;
  LAYER VI1 ;
  RECT 643.800 3.740 655.740 5.600 ;
  LAYER VI1 ;
  RECT 638.200 3.740 641.110 5.600 ;
  LAYER VI1 ;
  RECT 623.800 3.740 635.900 5.600 ;
  LAYER VI1 ;
  RECT 617.400 3.740 621.270 5.600 ;
  LAYER VI1 ;
  RECT 602.600 3.740 614.820 5.600 ;
  LAYER VI1 ;
  RECT 597.400 3.740 600.190 5.600 ;
  LAYER VI1 ;
  RECT 583.000 3.740 594.980 5.600 ;
  LAYER VI1 ;
  RECT 576.200 3.740 580.350 5.600 ;
  LAYER VI1 ;
  RECT 561.800 3.740 573.900 5.600 ;
  LAYER VI1 ;
  RECT 556.600 3.740 559.270 5.600 ;
  LAYER VI1 ;
  RECT 541.800 3.740 554.060 5.600 ;
  LAYER VI1 ;
  RECT 535.400 3.740 539.430 5.600 ;
  LAYER VI1 ;
  RECT 521.000 3.740 532.980 5.600 ;
  LAYER VI1 ;
  RECT 515.800 3.740 518.350 5.600 ;
  LAYER VI1 ;
  RECT 502.600 3.740 513.140 5.600 ;
  LAYER VI1 ;
  RECT 494.600 3.740 498.510 5.600 ;
  LAYER VI1 ;
  RECT 479.800 3.740 492.060 5.600 ;
  LAYER VI1 ;
  RECT 474.600 3.740 477.430 5.600 ;
  LAYER VI1 ;
  RECT 460.200 3.740 472.220 5.600 ;
  LAYER VI1 ;
  RECT 453.800 3.740 457.590 5.600 ;
  LAYER VI1 ;
  RECT 439.000 3.740 451.140 5.600 ;
  LAYER VI1 ;
  RECT 433.800 3.740 436.510 5.600 ;
  LAYER VI1 ;
  RECT 419.000 3.740 431.300 5.600 ;
  LAYER VI1 ;
  RECT 412.600 3.740 416.670 5.600 ;
  LAYER VI1 ;
  RECT 398.200 3.740 410.220 5.600 ;
  LAYER VI1 ;
  RECT 393.000 3.740 395.590 5.600 ;
  LAYER VI1 ;
  RECT 378.200 3.740 390.380 5.600 ;
  LAYER VI1 ;
  RECT 371.800 3.740 375.750 5.600 ;
  LAYER VI1 ;
  RECT 357.000 3.740 369.300 5.600 ;
  LAYER VI1 ;
  RECT 351.800 3.740 354.670 5.600 ;
  LAYER VI1 ;
  RECT 339.000 3.740 349.460 5.600 ;
  LAYER VI1 ;
  RECT 331.000 3.740 334.830 5.600 ;
  LAYER VI1 ;
  RECT 316.200 3.740 328.380 5.600 ;
  LAYER VI1 ;
  RECT 311.000 3.740 313.750 5.600 ;
  LAYER VI1 ;
  RECT 296.600 3.740 308.540 5.600 ;
  LAYER VI1 ;
  RECT 289.800 3.740 293.910 5.600 ;
  LAYER VI1 ;
  RECT 275.400 3.740 287.460 5.600 ;
  LAYER VI1 ;
  RECT 270.200 3.740 272.830 5.600 ;
  LAYER VI1 ;
  RECT 255.400 3.740 267.620 5.600 ;
  LAYER VI1 ;
  RECT 249.000 3.740 252.990 5.600 ;
  LAYER VI1 ;
  RECT 234.600 3.740 246.540 5.600 ;
  LAYER VI1 ;
  RECT 229.000 3.740 231.910 5.600 ;
  LAYER VI1 ;
  RECT 214.600 3.740 226.700 5.600 ;
  LAYER VI1 ;
  RECT 208.200 3.740 212.070 5.600 ;
  LAYER VI1 ;
  RECT 193.400 3.740 205.620 5.600 ;
  LAYER VI1 ;
  RECT 188.200 3.740 190.990 5.600 ;
  LAYER VI1 ;
  RECT 175.400 3.740 185.780 5.600 ;
  LAYER VI1 ;
  RECT 167.000 3.740 171.150 5.600 ;
  LAYER VI1 ;
  RECT 152.600 3.740 164.700 5.600 ;
  LAYER VI1 ;
  RECT 147.400 3.740 150.070 5.600 ;
  LAYER VI1 ;
  RECT 132.600 3.740 144.860 5.600 ;
  LAYER VI1 ;
  RECT 126.200 3.740 130.230 5.600 ;
  LAYER VI1 ;
  RECT 111.800 3.740 123.780 5.600 ;
  LAYER VI1 ;
  RECT 106.600 3.740 109.150 5.600 ;
  LAYER VI1 ;
  RECT 91.800 3.740 103.940 5.600 ;
  LAYER VI1 ;
  RECT 85.400 3.740 89.310 5.600 ;
  LAYER VI1 ;
  RECT 70.600 3.740 82.860 5.600 ;
  LAYER VI1 ;
  RECT 65.400 3.740 68.230 5.600 ;
  LAYER VI1 ;
  RECT 51.000 3.740 63.020 5.600 ;
  LAYER VI1 ;
  RECT 44.600 3.740 48.390 5.600 ;
  LAYER VI1 ;
  RECT 29.800 3.740 41.940 5.600 ;
  LAYER VI1 ;
  RECT 24.600 3.740 27.310 5.600 ;
  LAYER VI1 ;
  RECT 11.800 3.740 22.100 5.600 ;
  LAYER VI1 ;
  RECT 4.000 3.740 7.470 5.600 ;
  LAYER VI3 ;
  RECT 2.280 547.210 4.000 548.930 ;
  LAYER VI2 ;
  RECT 2.280 547.210 4.000 548.930 ;
  LAYER VI1 ;
  RECT 2.140 547.210 4.000 549.070 ;
  LAYER VI2 ;
  RECT 0.000 549.350 1.860 551.210 ;
  LAYER VI1 ;
  RECT 0.000 549.350 1.860 551.210 ;
  LAYER VI3 ;
  RECT 1375.500 3.880 1377.220 5.600 ;
  LAYER VI2 ;
  RECT 1375.500 3.880 1377.220 5.600 ;
  LAYER VI1 ;
  RECT 1375.500 3.740 1377.360 5.600 ;
  LAYER VI2 ;
  RECT 1377.640 1.600 1379.500 3.460 ;
  LAYER VI1 ;
  RECT 1377.640 1.600 1379.500 3.460 ;
  LAYER VI3 ;
  RECT 1375.500 547.210 1377.220 548.930 ;
  LAYER VI2 ;
  RECT 1375.500 547.210 1377.220 548.930 ;
  LAYER VI1 ;
  RECT 1375.500 547.210 1377.360 549.070 ;
  LAYER VI2 ;
  RECT 1377.640 549.350 1379.500 551.210 ;
  LAYER VI1 ;
  RECT 1377.640 549.350 1379.500 551.210 ;
  LAYER VI3 ;
  RECT 2.280 3.880 4.000 5.600 ;
  LAYER VI2 ;
  RECT 2.280 3.880 4.000 5.600 ;
  LAYER VI1 ;
  RECT 2.140 3.740 4.000 5.600 ;
  LAYER VI2 ;
  RECT 0.000 1.600 1.860 3.460 ;
  LAYER VI1 ;
  RECT 0.000 1.600 1.860 3.460 ;
  LAYER VI1 ;
  RECT 1367.600 0.200 1368.400 1.000 ;
  LAYER VI2 ;
  RECT 1367.600 0.200 1368.400 1.000 ;
  LAYER VI3 ;
  RECT 1367.600 0.200 1368.400 1.000 ;
  LAYER VI1 ;
  RECT 1352.800 0.200 1353.600 1.000 ;
  LAYER VI2 ;
  RECT 1352.800 0.200 1353.600 1.000 ;
  LAYER VI3 ;
  RECT 1352.800 0.200 1353.600 1.000 ;
  LAYER VI1 ;
  RECT 1347.600 0.200 1348.400 1.000 ;
  LAYER VI2 ;
  RECT 1347.600 0.200 1348.400 1.000 ;
  LAYER VI3 ;
  RECT 1347.600 0.200 1348.400 1.000 ;
  LAYER VI1 ;
  RECT 1333.200 0.200 1334.000 1.000 ;
  LAYER VI2 ;
  RECT 1333.200 0.200 1334.000 1.000 ;
  LAYER VI3 ;
  RECT 1333.200 0.200 1334.000 1.000 ;
  LAYER VI1 ;
  RECT 1326.800 0.200 1327.600 1.000 ;
  LAYER VI2 ;
  RECT 1326.800 0.200 1327.600 1.000 ;
  LAYER VI3 ;
  RECT 1326.800 0.200 1327.600 1.000 ;
  LAYER VI1 ;
  RECT 1312.000 0.200 1312.800 1.000 ;
  LAYER VI2 ;
  RECT 1312.000 0.200 1312.800 1.000 ;
  LAYER VI3 ;
  RECT 1312.000 0.200 1312.800 1.000 ;
  LAYER VI1 ;
  RECT 1306.800 0.200 1307.600 1.000 ;
  LAYER VI2 ;
  RECT 1306.800 0.200 1307.600 1.000 ;
  LAYER VI3 ;
  RECT 1306.800 0.200 1307.600 1.000 ;
  LAYER VI1 ;
  RECT 1292.000 0.200 1292.800 1.000 ;
  LAYER VI2 ;
  RECT 1292.000 0.200 1292.800 1.000 ;
  LAYER VI3 ;
  RECT 1292.000 0.200 1292.800 1.000 ;
  LAYER VI1 ;
  RECT 1285.600 0.200 1286.400 1.000 ;
  LAYER VI2 ;
  RECT 1285.600 0.200 1286.400 1.000 ;
  LAYER VI3 ;
  RECT 1285.600 0.200 1286.400 1.000 ;
  LAYER VI1 ;
  RECT 1271.200 0.200 1272.000 1.000 ;
  LAYER VI2 ;
  RECT 1271.200 0.200 1272.000 1.000 ;
  LAYER VI3 ;
  RECT 1271.200 0.200 1272.000 1.000 ;
  LAYER VI1 ;
  RECT 1266.000 0.200 1266.800 1.000 ;
  LAYER VI2 ;
  RECT 1266.000 0.200 1266.800 1.000 ;
  LAYER VI3 ;
  RECT 1266.000 0.200 1266.800 1.000 ;
  LAYER VI1 ;
  RECT 1251.200 0.200 1252.000 1.000 ;
  LAYER VI2 ;
  RECT 1251.200 0.200 1252.000 1.000 ;
  LAYER VI3 ;
  RECT 1251.200 0.200 1252.000 1.000 ;
  LAYER VI1 ;
  RECT 1244.800 0.200 1245.600 1.000 ;
  LAYER VI2 ;
  RECT 1244.800 0.200 1245.600 1.000 ;
  LAYER VI3 ;
  RECT 1244.800 0.200 1245.600 1.000 ;
  LAYER VI1 ;
  RECT 1230.000 0.200 1230.800 1.000 ;
  LAYER VI2 ;
  RECT 1230.000 0.200 1230.800 1.000 ;
  LAYER VI3 ;
  RECT 1230.000 0.200 1230.800 1.000 ;
  LAYER VI1 ;
  RECT 1224.800 0.200 1225.600 1.000 ;
  LAYER VI2 ;
  RECT 1224.800 0.200 1225.600 1.000 ;
  LAYER VI3 ;
  RECT 1224.800 0.200 1225.600 1.000 ;
  LAYER VI1 ;
  RECT 1212.000 0.200 1212.800 1.000 ;
  LAYER VI2 ;
  RECT 1212.000 0.200 1212.800 1.000 ;
  LAYER VI3 ;
  RECT 1212.000 0.200 1212.800 1.000 ;
  LAYER VI1 ;
  RECT 1210.400 0.200 1211.200 1.000 ;
  LAYER VI2 ;
  RECT 1210.400 0.200 1211.200 1.000 ;
  LAYER VI3 ;
  RECT 1210.400 0.200 1211.200 1.000 ;
  LAYER VI1 ;
  RECT 1204.000 0.200 1204.800 1.000 ;
  LAYER VI2 ;
  RECT 1204.000 0.200 1204.800 1.000 ;
  LAYER VI3 ;
  RECT 1204.000 0.200 1204.800 1.000 ;
  LAYER VI1 ;
  RECT 1189.200 0.200 1190.000 1.000 ;
  LAYER VI2 ;
  RECT 1189.200 0.200 1190.000 1.000 ;
  LAYER VI3 ;
  RECT 1189.200 0.200 1190.000 1.000 ;
  LAYER VI1 ;
  RECT 1184.000 0.200 1184.800 1.000 ;
  LAYER VI2 ;
  RECT 1184.000 0.200 1184.800 1.000 ;
  LAYER VI3 ;
  RECT 1184.000 0.200 1184.800 1.000 ;
  LAYER VI1 ;
  RECT 1169.200 0.200 1170.000 1.000 ;
  LAYER VI2 ;
  RECT 1169.200 0.200 1170.000 1.000 ;
  LAYER VI3 ;
  RECT 1169.200 0.200 1170.000 1.000 ;
  LAYER VI1 ;
  RECT 1162.800 0.200 1163.600 1.000 ;
  LAYER VI2 ;
  RECT 1162.800 0.200 1163.600 1.000 ;
  LAYER VI3 ;
  RECT 1162.800 0.200 1163.600 1.000 ;
  LAYER VI1 ;
  RECT 1148.400 0.200 1149.200 1.000 ;
  LAYER VI2 ;
  RECT 1148.400 0.200 1149.200 1.000 ;
  LAYER VI3 ;
  RECT 1148.400 0.200 1149.200 1.000 ;
  LAYER VI1 ;
  RECT 1143.200 0.200 1144.000 1.000 ;
  LAYER VI2 ;
  RECT 1143.200 0.200 1144.000 1.000 ;
  LAYER VI3 ;
  RECT 1143.200 0.200 1144.000 1.000 ;
  LAYER VI1 ;
  RECT 1128.400 0.200 1129.200 1.000 ;
  LAYER VI2 ;
  RECT 1128.400 0.200 1129.200 1.000 ;
  LAYER VI3 ;
  RECT 1128.400 0.200 1129.200 1.000 ;
  LAYER VI1 ;
  RECT 1122.000 0.200 1122.800 1.000 ;
  LAYER VI2 ;
  RECT 1122.000 0.200 1122.800 1.000 ;
  LAYER VI3 ;
  RECT 1122.000 0.200 1122.800 1.000 ;
  LAYER VI1 ;
  RECT 1107.200 0.200 1108.000 1.000 ;
  LAYER VI2 ;
  RECT 1107.200 0.200 1108.000 1.000 ;
  LAYER VI3 ;
  RECT 1107.200 0.200 1108.000 1.000 ;
  LAYER VI1 ;
  RECT 1102.000 0.200 1102.800 1.000 ;
  LAYER VI2 ;
  RECT 1102.000 0.200 1102.800 1.000 ;
  LAYER VI3 ;
  RECT 1102.000 0.200 1102.800 1.000 ;
  LAYER VI1 ;
  RECT 1087.600 0.200 1088.400 1.000 ;
  LAYER VI2 ;
  RECT 1087.600 0.200 1088.400 1.000 ;
  LAYER VI3 ;
  RECT 1087.600 0.200 1088.400 1.000 ;
  LAYER VI1 ;
  RECT 1081.200 0.200 1082.000 1.000 ;
  LAYER VI2 ;
  RECT 1081.200 0.200 1082.000 1.000 ;
  LAYER VI3 ;
  RECT 1081.200 0.200 1082.000 1.000 ;
  LAYER VI1 ;
  RECT 1066.400 0.200 1067.200 1.000 ;
  LAYER VI2 ;
  RECT 1066.400 0.200 1067.200 1.000 ;
  LAYER VI3 ;
  RECT 1066.400 0.200 1067.200 1.000 ;
  LAYER VI1 ;
  RECT 1061.200 0.200 1062.000 1.000 ;
  LAYER VI2 ;
  RECT 1061.200 0.200 1062.000 1.000 ;
  LAYER VI3 ;
  RECT 1061.200 0.200 1062.000 1.000 ;
  LAYER VI1 ;
  RECT 1048.400 0.200 1049.200 1.000 ;
  LAYER VI2 ;
  RECT 1048.400 0.200 1049.200 1.000 ;
  LAYER VI3 ;
  RECT 1048.400 0.200 1049.200 1.000 ;
  LAYER VI1 ;
  RECT 1046.800 0.200 1047.600 1.000 ;
  LAYER VI2 ;
  RECT 1046.800 0.200 1047.600 1.000 ;
  LAYER VI3 ;
  RECT 1046.800 0.200 1047.600 1.000 ;
  LAYER VI1 ;
  RECT 1040.000 0.200 1040.800 1.000 ;
  LAYER VI2 ;
  RECT 1040.000 0.200 1040.800 1.000 ;
  LAYER VI3 ;
  RECT 1040.000 0.200 1040.800 1.000 ;
  LAYER VI1 ;
  RECT 1025.600 0.200 1026.400 1.000 ;
  LAYER VI2 ;
  RECT 1025.600 0.200 1026.400 1.000 ;
  LAYER VI3 ;
  RECT 1025.600 0.200 1026.400 1.000 ;
  LAYER VI1 ;
  RECT 1020.400 0.200 1021.200 1.000 ;
  LAYER VI2 ;
  RECT 1020.400 0.200 1021.200 1.000 ;
  LAYER VI3 ;
  RECT 1020.400 0.200 1021.200 1.000 ;
  LAYER VI1 ;
  RECT 1005.600 0.200 1006.400 1.000 ;
  LAYER VI2 ;
  RECT 1005.600 0.200 1006.400 1.000 ;
  LAYER VI3 ;
  RECT 1005.600 0.200 1006.400 1.000 ;
  LAYER VI1 ;
  RECT 999.200 0.200 1000.000 1.000 ;
  LAYER VI2 ;
  RECT 999.200 0.200 1000.000 1.000 ;
  LAYER VI3 ;
  RECT 999.200 0.200 1000.000 1.000 ;
  LAYER VI1 ;
  RECT 984.800 0.200 985.600 1.000 ;
  LAYER VI2 ;
  RECT 984.800 0.200 985.600 1.000 ;
  LAYER VI3 ;
  RECT 984.800 0.200 985.600 1.000 ;
  LAYER VI1 ;
  RECT 979.600 0.200 980.400 1.000 ;
  LAYER VI2 ;
  RECT 979.600 0.200 980.400 1.000 ;
  LAYER VI3 ;
  RECT 979.600 0.200 980.400 1.000 ;
  LAYER VI1 ;
  RECT 964.800 0.200 965.600 1.000 ;
  LAYER VI2 ;
  RECT 964.800 0.200 965.600 1.000 ;
  LAYER VI3 ;
  RECT 964.800 0.200 965.600 1.000 ;
  LAYER VI1 ;
  RECT 958.400 0.200 959.200 1.000 ;
  LAYER VI2 ;
  RECT 958.400 0.200 959.200 1.000 ;
  LAYER VI3 ;
  RECT 958.400 0.200 959.200 1.000 ;
  LAYER VI1 ;
  RECT 943.600 0.200 944.400 1.000 ;
  LAYER VI2 ;
  RECT 943.600 0.200 944.400 1.000 ;
  LAYER VI3 ;
  RECT 943.600 0.200 944.400 1.000 ;
  LAYER VI1 ;
  RECT 938.400 0.200 939.200 1.000 ;
  LAYER VI2 ;
  RECT 938.400 0.200 939.200 1.000 ;
  LAYER VI3 ;
  RECT 938.400 0.200 939.200 1.000 ;
  LAYER VI1 ;
  RECT 924.000 0.200 924.800 1.000 ;
  LAYER VI2 ;
  RECT 924.000 0.200 924.800 1.000 ;
  LAYER VI3 ;
  RECT 924.000 0.200 924.800 1.000 ;
  LAYER VI1 ;
  RECT 917.600 0.200 918.400 1.000 ;
  LAYER VI2 ;
  RECT 917.600 0.200 918.400 1.000 ;
  LAYER VI3 ;
  RECT 917.600 0.200 918.400 1.000 ;
  LAYER VI1 ;
  RECT 902.800 0.200 903.600 1.000 ;
  LAYER VI2 ;
  RECT 902.800 0.200 903.600 1.000 ;
  LAYER VI3 ;
  RECT 902.800 0.200 903.600 1.000 ;
  LAYER VI1 ;
  RECT 897.600 0.200 898.400 1.000 ;
  LAYER VI2 ;
  RECT 897.600 0.200 898.400 1.000 ;
  LAYER VI3 ;
  RECT 897.600 0.200 898.400 1.000 ;
  LAYER VI1 ;
  RECT 884.800 0.200 885.600 1.000 ;
  LAYER VI2 ;
  RECT 884.800 0.200 885.600 1.000 ;
  LAYER VI3 ;
  RECT 884.800 0.200 885.600 1.000 ;
  LAYER VI1 ;
  RECT 882.800 0.200 883.600 1.000 ;
  LAYER VI2 ;
  RECT 882.800 0.200 883.600 1.000 ;
  LAYER VI3 ;
  RECT 882.800 0.200 883.600 1.000 ;
  LAYER VI1 ;
  RECT 876.400 0.200 877.200 1.000 ;
  LAYER VI2 ;
  RECT 876.400 0.200 877.200 1.000 ;
  LAYER VI3 ;
  RECT 876.400 0.200 877.200 1.000 ;
  LAYER VI1 ;
  RECT 862.000 0.200 862.800 1.000 ;
  LAYER VI2 ;
  RECT 862.000 0.200 862.800 1.000 ;
  LAYER VI3 ;
  RECT 862.000 0.200 862.800 1.000 ;
  LAYER VI1 ;
  RECT 856.800 0.200 857.600 1.000 ;
  LAYER VI2 ;
  RECT 856.800 0.200 857.600 1.000 ;
  LAYER VI3 ;
  RECT 856.800 0.200 857.600 1.000 ;
  LAYER VI1 ;
  RECT 842.000 0.200 842.800 1.000 ;
  LAYER VI2 ;
  RECT 842.000 0.200 842.800 1.000 ;
  LAYER VI3 ;
  RECT 842.000 0.200 842.800 1.000 ;
  LAYER VI1 ;
  RECT 835.600 0.200 836.400 1.000 ;
  LAYER VI2 ;
  RECT 835.600 0.200 836.400 1.000 ;
  LAYER VI3 ;
  RECT 835.600 0.200 836.400 1.000 ;
  LAYER VI1 ;
  RECT 820.800 0.200 821.600 1.000 ;
  LAYER VI2 ;
  RECT 820.800 0.200 821.600 1.000 ;
  LAYER VI3 ;
  RECT 820.800 0.200 821.600 1.000 ;
  LAYER VI1 ;
  RECT 815.600 0.200 816.400 1.000 ;
  LAYER VI2 ;
  RECT 815.600 0.200 816.400 1.000 ;
  LAYER VI3 ;
  RECT 815.600 0.200 816.400 1.000 ;
  LAYER VI1 ;
  RECT 801.200 0.200 802.000 1.000 ;
  LAYER VI2 ;
  RECT 801.200 0.200 802.000 1.000 ;
  LAYER VI3 ;
  RECT 801.200 0.200 802.000 1.000 ;
  LAYER VI1 ;
  RECT 794.800 0.200 795.600 1.000 ;
  LAYER VI2 ;
  RECT 794.800 0.200 795.600 1.000 ;
  LAYER VI3 ;
  RECT 794.800 0.200 795.600 1.000 ;
  LAYER VI1 ;
  RECT 780.000 0.200 780.800 1.000 ;
  LAYER VI2 ;
  RECT 780.000 0.200 780.800 1.000 ;
  LAYER VI3 ;
  RECT 780.000 0.200 780.800 1.000 ;
  LAYER VI1 ;
  RECT 774.800 0.200 775.600 1.000 ;
  LAYER VI2 ;
  RECT 774.800 0.200 775.600 1.000 ;
  LAYER VI3 ;
  RECT 774.800 0.200 775.600 1.000 ;
  LAYER VI1 ;
  RECT 760.000 0.200 760.800 1.000 ;
  LAYER VI2 ;
  RECT 760.000 0.200 760.800 1.000 ;
  LAYER VI3 ;
  RECT 760.000 0.200 760.800 1.000 ;
  LAYER VI1 ;
  RECT 753.600 0.200 754.400 1.000 ;
  LAYER VI2 ;
  RECT 753.600 0.200 754.400 1.000 ;
  LAYER VI3 ;
  RECT 753.600 0.200 754.400 1.000 ;
  LAYER VI1 ;
  RECT 739.200 0.200 740.000 1.000 ;
  LAYER VI2 ;
  RECT 739.200 0.200 740.000 1.000 ;
  LAYER VI3 ;
  RECT 739.200 0.200 740.000 1.000 ;
  LAYER VI1 ;
  RECT 734.000 0.200 734.800 1.000 ;
  LAYER VI2 ;
  RECT 734.000 0.200 734.800 1.000 ;
  LAYER VI3 ;
  RECT 734.000 0.200 734.800 1.000 ;
  LAYER VI1 ;
  RECT 720.800 0.200 721.600 1.000 ;
  LAYER VI2 ;
  RECT 720.800 0.200 721.600 1.000 ;
  LAYER VI3 ;
  RECT 720.800 0.200 721.600 1.000 ;
  LAYER VI1 ;
  RECT 719.200 0.200 720.000 1.000 ;
  LAYER VI2 ;
  RECT 719.200 0.200 720.000 1.000 ;
  LAYER VI3 ;
  RECT 719.200 0.200 720.000 1.000 ;
  LAYER VI1 ;
  RECT 698.400 0.200 699.200 1.000 ;
  LAYER VI2 ;
  RECT 698.400 0.200 699.200 1.000 ;
  LAYER VI3 ;
  RECT 698.400 0.200 699.200 1.000 ;
  LAYER VI1 ;
  RECT 697.200 0.200 698.000 1.000 ;
  LAYER VI2 ;
  RECT 697.200 0.200 698.000 1.000 ;
  LAYER VI3 ;
  RECT 697.200 0.200 698.000 1.000 ;
  LAYER VI1 ;
  RECT 696.000 0.200 696.800 1.000 ;
  LAYER VI2 ;
  RECT 696.000 0.200 696.800 1.000 ;
  LAYER VI3 ;
  RECT 696.000 0.200 696.800 1.000 ;
  LAYER VI1 ;
  RECT 694.800 0.200 695.600 1.000 ;
  LAYER VI2 ;
  RECT 694.800 0.200 695.600 1.000 ;
  LAYER VI3 ;
  RECT 694.800 0.200 695.600 1.000 ;
  LAYER VI1 ;
  RECT 693.600 0.200 694.400 1.000 ;
  LAYER VI2 ;
  RECT 693.600 0.200 694.400 1.000 ;
  LAYER VI3 ;
  RECT 693.600 0.200 694.400 1.000 ;
  LAYER VI1 ;
  RECT 692.400 0.200 693.200 1.000 ;
  LAYER VI2 ;
  RECT 692.400 0.200 693.200 1.000 ;
  LAYER VI3 ;
  RECT 692.400 0.200 693.200 1.000 ;
  LAYER VI1 ;
  RECT 686.400 0.200 687.200 1.000 ;
  LAYER VI2 ;
  RECT 686.400 0.200 687.200 1.000 ;
  LAYER VI3 ;
  RECT 686.400 0.200 687.200 1.000 ;
  LAYER VI1 ;
  RECT 679.200 0.200 680.000 1.000 ;
  LAYER VI2 ;
  RECT 679.200 0.200 680.000 1.000 ;
  LAYER VI3 ;
  RECT 679.200 0.200 680.000 1.000 ;
  LAYER VI1 ;
  RECT 676.800 0.200 677.600 1.000 ;
  LAYER VI2 ;
  RECT 676.800 0.200 677.600 1.000 ;
  LAYER VI3 ;
  RECT 676.800 0.200 677.600 1.000 ;
  LAYER VI1 ;
  RECT 674.000 0.200 674.800 1.000 ;
  LAYER VI2 ;
  RECT 674.000 0.200 674.800 1.000 ;
  LAYER VI3 ;
  RECT 674.000 0.200 674.800 1.000 ;
  LAYER VI1 ;
  RECT 671.200 0.200 672.000 1.000 ;
  LAYER VI2 ;
  RECT 671.200 0.200 672.000 1.000 ;
  LAYER VI3 ;
  RECT 671.200 0.200 672.000 1.000 ;
  LAYER VI1 ;
  RECT 670.000 0.200 670.800 1.000 ;
  LAYER VI2 ;
  RECT 670.000 0.200 670.800 1.000 ;
  LAYER VI3 ;
  RECT 670.000 0.200 670.800 1.000 ;
  LAYER VI1 ;
  RECT 667.200 0.200 668.000 1.000 ;
  LAYER VI2 ;
  RECT 667.200 0.200 668.000 1.000 ;
  LAYER VI3 ;
  RECT 667.200 0.200 668.000 1.000 ;
  LAYER VI1 ;
  RECT 666.000 0.200 666.800 1.000 ;
  LAYER VI2 ;
  RECT 666.000 0.200 666.800 1.000 ;
  LAYER VI3 ;
  RECT 666.000 0.200 666.800 1.000 ;
  LAYER VI1 ;
  RECT 663.200 0.200 664.000 1.000 ;
  LAYER VI2 ;
  RECT 663.200 0.200 664.000 1.000 ;
  LAYER VI3 ;
  RECT 663.200 0.200 664.000 1.000 ;
  LAYER VI1 ;
  RECT 656.400 0.200 657.200 1.000 ;
  LAYER VI2 ;
  RECT 656.400 0.200 657.200 1.000 ;
  LAYER VI3 ;
  RECT 656.400 0.200 657.200 1.000 ;
  LAYER VI1 ;
  RECT 642.000 0.200 642.800 1.000 ;
  LAYER VI2 ;
  RECT 642.000 0.200 642.800 1.000 ;
  LAYER VI3 ;
  RECT 642.000 0.200 642.800 1.000 ;
  LAYER VI1 ;
  RECT 636.400 0.200 637.200 1.000 ;
  LAYER VI2 ;
  RECT 636.400 0.200 637.200 1.000 ;
  LAYER VI3 ;
  RECT 636.400 0.200 637.200 1.000 ;
  LAYER VI1 ;
  RECT 622.000 0.200 622.800 1.000 ;
  LAYER VI2 ;
  RECT 622.000 0.200 622.800 1.000 ;
  LAYER VI3 ;
  RECT 622.000 0.200 622.800 1.000 ;
  LAYER VI1 ;
  RECT 615.600 0.200 616.400 1.000 ;
  LAYER VI2 ;
  RECT 615.600 0.200 616.400 1.000 ;
  LAYER VI3 ;
  RECT 615.600 0.200 616.400 1.000 ;
  LAYER VI1 ;
  RECT 600.800 0.200 601.600 1.000 ;
  LAYER VI2 ;
  RECT 600.800 0.200 601.600 1.000 ;
  LAYER VI3 ;
  RECT 600.800 0.200 601.600 1.000 ;
  LAYER VI1 ;
  RECT 595.600 0.200 596.400 1.000 ;
  LAYER VI2 ;
  RECT 595.600 0.200 596.400 1.000 ;
  LAYER VI3 ;
  RECT 595.600 0.200 596.400 1.000 ;
  LAYER VI1 ;
  RECT 581.200 0.200 582.000 1.000 ;
  LAYER VI2 ;
  RECT 581.200 0.200 582.000 1.000 ;
  LAYER VI3 ;
  RECT 581.200 0.200 582.000 1.000 ;
  LAYER VI1 ;
  RECT 574.400 0.200 575.200 1.000 ;
  LAYER VI2 ;
  RECT 574.400 0.200 575.200 1.000 ;
  LAYER VI3 ;
  RECT 574.400 0.200 575.200 1.000 ;
  LAYER VI1 ;
  RECT 560.000 0.200 560.800 1.000 ;
  LAYER VI2 ;
  RECT 560.000 0.200 560.800 1.000 ;
  LAYER VI3 ;
  RECT 560.000 0.200 560.800 1.000 ;
  LAYER VI1 ;
  RECT 554.800 0.200 555.600 1.000 ;
  LAYER VI2 ;
  RECT 554.800 0.200 555.600 1.000 ;
  LAYER VI3 ;
  RECT 554.800 0.200 555.600 1.000 ;
  LAYER VI1 ;
  RECT 540.000 0.200 540.800 1.000 ;
  LAYER VI2 ;
  RECT 540.000 0.200 540.800 1.000 ;
  LAYER VI3 ;
  RECT 540.000 0.200 540.800 1.000 ;
  LAYER VI1 ;
  RECT 533.600 0.200 534.400 1.000 ;
  LAYER VI2 ;
  RECT 533.600 0.200 534.400 1.000 ;
  LAYER VI3 ;
  RECT 533.600 0.200 534.400 1.000 ;
  LAYER VI1 ;
  RECT 519.200 0.200 520.000 1.000 ;
  LAYER VI2 ;
  RECT 519.200 0.200 520.000 1.000 ;
  LAYER VI3 ;
  RECT 519.200 0.200 520.000 1.000 ;
  LAYER VI1 ;
  RECT 514.000 0.200 514.800 1.000 ;
  LAYER VI2 ;
  RECT 514.000 0.200 514.800 1.000 ;
  LAYER VI3 ;
  RECT 514.000 0.200 514.800 1.000 ;
  LAYER VI1 ;
  RECT 500.800 0.200 501.600 1.000 ;
  LAYER VI2 ;
  RECT 500.800 0.200 501.600 1.000 ;
  LAYER VI3 ;
  RECT 500.800 0.200 501.600 1.000 ;
  LAYER VI1 ;
  RECT 499.200 0.200 500.000 1.000 ;
  LAYER VI2 ;
  RECT 499.200 0.200 500.000 1.000 ;
  LAYER VI3 ;
  RECT 499.200 0.200 500.000 1.000 ;
  LAYER VI1 ;
  RECT 492.800 0.200 493.600 1.000 ;
  LAYER VI2 ;
  RECT 492.800 0.200 493.600 1.000 ;
  LAYER VI3 ;
  RECT 492.800 0.200 493.600 1.000 ;
  LAYER VI1 ;
  RECT 478.000 0.200 478.800 1.000 ;
  LAYER VI2 ;
  RECT 478.000 0.200 478.800 1.000 ;
  LAYER VI3 ;
  RECT 478.000 0.200 478.800 1.000 ;
  LAYER VI1 ;
  RECT 472.800 0.200 473.600 1.000 ;
  LAYER VI2 ;
  RECT 472.800 0.200 473.600 1.000 ;
  LAYER VI3 ;
  RECT 472.800 0.200 473.600 1.000 ;
  LAYER VI1 ;
  RECT 458.400 0.200 459.200 1.000 ;
  LAYER VI2 ;
  RECT 458.400 0.200 459.200 1.000 ;
  LAYER VI3 ;
  RECT 458.400 0.200 459.200 1.000 ;
  LAYER VI1 ;
  RECT 452.000 0.200 452.800 1.000 ;
  LAYER VI2 ;
  RECT 452.000 0.200 452.800 1.000 ;
  LAYER VI3 ;
  RECT 452.000 0.200 452.800 1.000 ;
  LAYER VI1 ;
  RECT 437.200 0.200 438.000 1.000 ;
  LAYER VI2 ;
  RECT 437.200 0.200 438.000 1.000 ;
  LAYER VI3 ;
  RECT 437.200 0.200 438.000 1.000 ;
  LAYER VI1 ;
  RECT 432.000 0.200 432.800 1.000 ;
  LAYER VI2 ;
  RECT 432.000 0.200 432.800 1.000 ;
  LAYER VI3 ;
  RECT 432.000 0.200 432.800 1.000 ;
  LAYER VI1 ;
  RECT 417.200 0.200 418.000 1.000 ;
  LAYER VI2 ;
  RECT 417.200 0.200 418.000 1.000 ;
  LAYER VI3 ;
  RECT 417.200 0.200 418.000 1.000 ;
  LAYER VI1 ;
  RECT 410.800 0.200 411.600 1.000 ;
  LAYER VI2 ;
  RECT 410.800 0.200 411.600 1.000 ;
  LAYER VI3 ;
  RECT 410.800 0.200 411.600 1.000 ;
  LAYER VI1 ;
  RECT 396.400 0.200 397.200 1.000 ;
  LAYER VI2 ;
  RECT 396.400 0.200 397.200 1.000 ;
  LAYER VI3 ;
  RECT 396.400 0.200 397.200 1.000 ;
  LAYER VI1 ;
  RECT 391.200 0.200 392.000 1.000 ;
  LAYER VI2 ;
  RECT 391.200 0.200 392.000 1.000 ;
  LAYER VI3 ;
  RECT 391.200 0.200 392.000 1.000 ;
  LAYER VI1 ;
  RECT 376.400 0.200 377.200 1.000 ;
  LAYER VI2 ;
  RECT 376.400 0.200 377.200 1.000 ;
  LAYER VI3 ;
  RECT 376.400 0.200 377.200 1.000 ;
  LAYER VI1 ;
  RECT 370.000 0.200 370.800 1.000 ;
  LAYER VI2 ;
  RECT 370.000 0.200 370.800 1.000 ;
  LAYER VI3 ;
  RECT 370.000 0.200 370.800 1.000 ;
  LAYER VI1 ;
  RECT 355.200 0.200 356.000 1.000 ;
  LAYER VI2 ;
  RECT 355.200 0.200 356.000 1.000 ;
  LAYER VI3 ;
  RECT 355.200 0.200 356.000 1.000 ;
  LAYER VI1 ;
  RECT 350.000 0.200 350.800 1.000 ;
  LAYER VI2 ;
  RECT 350.000 0.200 350.800 1.000 ;
  LAYER VI3 ;
  RECT 350.000 0.200 350.800 1.000 ;
  LAYER VI1 ;
  RECT 337.200 0.200 338.000 1.000 ;
  LAYER VI2 ;
  RECT 337.200 0.200 338.000 1.000 ;
  LAYER VI3 ;
  RECT 337.200 0.200 338.000 1.000 ;
  LAYER VI1 ;
  RECT 335.600 0.200 336.400 1.000 ;
  LAYER VI2 ;
  RECT 335.600 0.200 336.400 1.000 ;
  LAYER VI3 ;
  RECT 335.600 0.200 336.400 1.000 ;
  LAYER VI1 ;
  RECT 329.200 0.200 330.000 1.000 ;
  LAYER VI2 ;
  RECT 329.200 0.200 330.000 1.000 ;
  LAYER VI3 ;
  RECT 329.200 0.200 330.000 1.000 ;
  LAYER VI1 ;
  RECT 314.400 0.200 315.200 1.000 ;
  LAYER VI2 ;
  RECT 314.400 0.200 315.200 1.000 ;
  LAYER VI3 ;
  RECT 314.400 0.200 315.200 1.000 ;
  LAYER VI1 ;
  RECT 309.200 0.200 310.000 1.000 ;
  LAYER VI2 ;
  RECT 309.200 0.200 310.000 1.000 ;
  LAYER VI3 ;
  RECT 309.200 0.200 310.000 1.000 ;
  LAYER VI1 ;
  RECT 294.800 0.200 295.600 1.000 ;
  LAYER VI2 ;
  RECT 294.800 0.200 295.600 1.000 ;
  LAYER VI3 ;
  RECT 294.800 0.200 295.600 1.000 ;
  LAYER VI1 ;
  RECT 288.000 0.200 288.800 1.000 ;
  LAYER VI2 ;
  RECT 288.000 0.200 288.800 1.000 ;
  LAYER VI3 ;
  RECT 288.000 0.200 288.800 1.000 ;
  LAYER VI1 ;
  RECT 273.600 0.200 274.400 1.000 ;
  LAYER VI2 ;
  RECT 273.600 0.200 274.400 1.000 ;
  LAYER VI3 ;
  RECT 273.600 0.200 274.400 1.000 ;
  LAYER VI1 ;
  RECT 268.400 0.200 269.200 1.000 ;
  LAYER VI2 ;
  RECT 268.400 0.200 269.200 1.000 ;
  LAYER VI3 ;
  RECT 268.400 0.200 269.200 1.000 ;
  LAYER VI1 ;
  RECT 253.600 0.200 254.400 1.000 ;
  LAYER VI2 ;
  RECT 253.600 0.200 254.400 1.000 ;
  LAYER VI3 ;
  RECT 253.600 0.200 254.400 1.000 ;
  LAYER VI1 ;
  RECT 247.200 0.200 248.000 1.000 ;
  LAYER VI2 ;
  RECT 247.200 0.200 248.000 1.000 ;
  LAYER VI3 ;
  RECT 247.200 0.200 248.000 1.000 ;
  LAYER VI1 ;
  RECT 232.800 0.200 233.600 1.000 ;
  LAYER VI2 ;
  RECT 232.800 0.200 233.600 1.000 ;
  LAYER VI3 ;
  RECT 232.800 0.200 233.600 1.000 ;
  LAYER VI1 ;
  RECT 227.200 0.200 228.000 1.000 ;
  LAYER VI2 ;
  RECT 227.200 0.200 228.000 1.000 ;
  LAYER VI3 ;
  RECT 227.200 0.200 228.000 1.000 ;
  LAYER VI1 ;
  RECT 212.800 0.200 213.600 1.000 ;
  LAYER VI2 ;
  RECT 212.800 0.200 213.600 1.000 ;
  LAYER VI3 ;
  RECT 212.800 0.200 213.600 1.000 ;
  LAYER VI1 ;
  RECT 206.400 0.200 207.200 1.000 ;
  LAYER VI2 ;
  RECT 206.400 0.200 207.200 1.000 ;
  LAYER VI3 ;
  RECT 206.400 0.200 207.200 1.000 ;
  LAYER VI1 ;
  RECT 191.600 0.200 192.400 1.000 ;
  LAYER VI2 ;
  RECT 191.600 0.200 192.400 1.000 ;
  LAYER VI3 ;
  RECT 191.600 0.200 192.400 1.000 ;
  LAYER VI1 ;
  RECT 186.400 0.200 187.200 1.000 ;
  LAYER VI2 ;
  RECT 186.400 0.200 187.200 1.000 ;
  LAYER VI3 ;
  RECT 186.400 0.200 187.200 1.000 ;
  LAYER VI1 ;
  RECT 173.600 0.200 174.400 1.000 ;
  LAYER VI2 ;
  RECT 173.600 0.200 174.400 1.000 ;
  LAYER VI3 ;
  RECT 173.600 0.200 174.400 1.000 ;
  LAYER VI1 ;
  RECT 172.000 0.200 172.800 1.000 ;
  LAYER VI2 ;
  RECT 172.000 0.200 172.800 1.000 ;
  LAYER VI3 ;
  RECT 172.000 0.200 172.800 1.000 ;
  LAYER VI1 ;
  RECT 165.200 0.200 166.000 1.000 ;
  LAYER VI2 ;
  RECT 165.200 0.200 166.000 1.000 ;
  LAYER VI3 ;
  RECT 165.200 0.200 166.000 1.000 ;
  LAYER VI1 ;
  RECT 150.800 0.200 151.600 1.000 ;
  LAYER VI2 ;
  RECT 150.800 0.200 151.600 1.000 ;
  LAYER VI3 ;
  RECT 150.800 0.200 151.600 1.000 ;
  LAYER VI1 ;
  RECT 145.600 0.200 146.400 1.000 ;
  LAYER VI2 ;
  RECT 145.600 0.200 146.400 1.000 ;
  LAYER VI3 ;
  RECT 145.600 0.200 146.400 1.000 ;
  LAYER VI1 ;
  RECT 130.800 0.200 131.600 1.000 ;
  LAYER VI2 ;
  RECT 130.800 0.200 131.600 1.000 ;
  LAYER VI3 ;
  RECT 130.800 0.200 131.600 1.000 ;
  LAYER VI1 ;
  RECT 124.400 0.200 125.200 1.000 ;
  LAYER VI2 ;
  RECT 124.400 0.200 125.200 1.000 ;
  LAYER VI3 ;
  RECT 124.400 0.200 125.200 1.000 ;
  LAYER VI1 ;
  RECT 110.000 0.200 110.800 1.000 ;
  LAYER VI2 ;
  RECT 110.000 0.200 110.800 1.000 ;
  LAYER VI3 ;
  RECT 110.000 0.200 110.800 1.000 ;
  LAYER VI1 ;
  RECT 104.800 0.200 105.600 1.000 ;
  LAYER VI2 ;
  RECT 104.800 0.200 105.600 1.000 ;
  LAYER VI3 ;
  RECT 104.800 0.200 105.600 1.000 ;
  LAYER VI1 ;
  RECT 90.000 0.200 90.800 1.000 ;
  LAYER VI2 ;
  RECT 90.000 0.200 90.800 1.000 ;
  LAYER VI3 ;
  RECT 90.000 0.200 90.800 1.000 ;
  LAYER VI1 ;
  RECT 83.600 0.200 84.400 1.000 ;
  LAYER VI2 ;
  RECT 83.600 0.200 84.400 1.000 ;
  LAYER VI3 ;
  RECT 83.600 0.200 84.400 1.000 ;
  LAYER VI1 ;
  RECT 68.800 0.200 69.600 1.000 ;
  LAYER VI2 ;
  RECT 68.800 0.200 69.600 1.000 ;
  LAYER VI3 ;
  RECT 68.800 0.200 69.600 1.000 ;
  LAYER VI1 ;
  RECT 63.600 0.200 64.400 1.000 ;
  LAYER VI2 ;
  RECT 63.600 0.200 64.400 1.000 ;
  LAYER VI3 ;
  RECT 63.600 0.200 64.400 1.000 ;
  LAYER VI1 ;
  RECT 49.200 0.200 50.000 1.000 ;
  LAYER VI2 ;
  RECT 49.200 0.200 50.000 1.000 ;
  LAYER VI3 ;
  RECT 49.200 0.200 50.000 1.000 ;
  LAYER VI1 ;
  RECT 42.800 0.200 43.600 1.000 ;
  LAYER VI2 ;
  RECT 42.800 0.200 43.600 1.000 ;
  LAYER VI3 ;
  RECT 42.800 0.200 43.600 1.000 ;
  LAYER VI1 ;
  RECT 28.000 0.200 28.800 1.000 ;
  LAYER VI2 ;
  RECT 28.000 0.200 28.800 1.000 ;
  LAYER VI3 ;
  RECT 28.000 0.200 28.800 1.000 ;
  LAYER VI1 ;
  RECT 22.800 0.200 23.600 1.000 ;
  LAYER VI2 ;
  RECT 22.800 0.200 23.600 1.000 ;
  LAYER VI3 ;
  RECT 22.800 0.200 23.600 1.000 ;
  LAYER VI1 ;
  RECT 10.000 0.200 10.800 1.000 ;
  LAYER VI2 ;
  RECT 10.000 0.200 10.800 1.000 ;
  LAYER VI3 ;
  RECT 10.000 0.200 10.800 1.000 ;
  LAYER VI1 ;
  RECT 8.000 0.200 8.800 1.000 ;
  LAYER VI2 ;
  RECT 8.000 0.200 8.800 1.000 ;
  LAYER VI3 ;
  RECT 8.000 0.200 8.800 1.000 ;
  LAYER VI3 ;
  RECT 1374.360 9.570 1375.220 11.170 ;
  LAYER VI3 ;
  RECT 1374.820 10.770 1375.020 10.970 ;
  LAYER VI3 ;
  RECT 1374.820 10.370 1375.020 10.570 ;
  LAYER VI3 ;
  RECT 1374.820 9.970 1375.020 10.170 ;
  LAYER VI3 ;
  RECT 1374.820 9.570 1375.020 9.770 ;
  LAYER VI3 ;
  RECT 1374.420 10.770 1374.620 10.970 ;
  LAYER VI3 ;
  RECT 1374.420 10.370 1374.620 10.570 ;
  LAYER VI3 ;
  RECT 1374.420 9.970 1374.620 10.170 ;
  LAYER VI3 ;
  RECT 1374.420 9.570 1374.620 9.770 ;
  LAYER VI2 ;
  RECT 1374.360 9.570 1375.220 11.170 ;
  LAYER VI2 ;
  RECT 1374.820 10.770 1375.020 10.970 ;
  LAYER VI2 ;
  RECT 1374.820 10.370 1375.020 10.570 ;
  LAYER VI2 ;
  RECT 1374.820 9.970 1375.020 10.170 ;
  LAYER VI2 ;
  RECT 1374.820 9.570 1375.020 9.770 ;
  LAYER VI2 ;
  RECT 1374.420 10.770 1374.620 10.970 ;
  LAYER VI2 ;
  RECT 1374.420 10.370 1374.620 10.570 ;
  LAYER VI2 ;
  RECT 1374.420 9.970 1374.620 10.170 ;
  LAYER VI2 ;
  RECT 1374.420 9.570 1374.620 9.770 ;
  LAYER VI3 ;
  RECT 1374.360 14.200 1375.220 15.200 ;
  LAYER VI3 ;
  RECT 1374.820 14.600 1375.020 14.800 ;
  LAYER VI3 ;
  RECT 1374.820 14.200 1375.020 14.400 ;
  LAYER VI3 ;
  RECT 1374.420 14.600 1374.620 14.800 ;
  LAYER VI3 ;
  RECT 1374.420 14.200 1374.620 14.400 ;
  LAYER VI2 ;
  RECT 1374.360 14.200 1375.220 15.200 ;
  LAYER VI2 ;
  RECT 1374.820 14.600 1375.020 14.800 ;
  LAYER VI2 ;
  RECT 1374.820 14.200 1375.020 14.400 ;
  LAYER VI2 ;
  RECT 1374.420 14.600 1374.620 14.800 ;
  LAYER VI2 ;
  RECT 1374.420 14.200 1374.620 14.400 ;
  LAYER VI3 ;
  RECT 1374.360 18.730 1375.220 19.730 ;
  LAYER VI3 ;
  RECT 1374.820 19.130 1375.020 19.330 ;
  LAYER VI3 ;
  RECT 1374.820 18.730 1375.020 18.930 ;
  LAYER VI3 ;
  RECT 1374.420 19.130 1374.620 19.330 ;
  LAYER VI3 ;
  RECT 1374.420 18.730 1374.620 18.930 ;
  LAYER VI2 ;
  RECT 1374.360 18.730 1375.220 19.730 ;
  LAYER VI2 ;
  RECT 1374.820 19.130 1375.020 19.330 ;
  LAYER VI2 ;
  RECT 1374.820 18.730 1375.020 18.930 ;
  LAYER VI2 ;
  RECT 1374.420 19.130 1374.620 19.330 ;
  LAYER VI2 ;
  RECT 1374.420 18.730 1374.620 18.930 ;
  LAYER VI3 ;
  RECT 1374.360 21.230 1375.220 22.070 ;
  LAYER VI3 ;
  RECT 1374.760 21.690 1374.960 21.890 ;
  LAYER VI3 ;
  RECT 1374.760 21.290 1374.960 21.490 ;
  LAYER VI3 ;
  RECT 1374.360 21.690 1374.560 21.890 ;
  LAYER VI3 ;
  RECT 1374.360 21.290 1374.560 21.490 ;
  LAYER VI2 ;
  RECT 1374.360 21.230 1375.220 22.070 ;
  LAYER VI2 ;
  RECT 1374.760 21.690 1374.960 21.890 ;
  LAYER VI2 ;
  RECT 1374.760 21.290 1374.960 21.490 ;
  LAYER VI2 ;
  RECT 1374.360 21.690 1374.560 21.890 ;
  LAYER VI2 ;
  RECT 1374.360 21.290 1374.560 21.490 ;
  LAYER VI3 ;
  RECT 1374.360 24.170 1375.220 25.170 ;
  LAYER VI3 ;
  RECT 1374.820 24.570 1375.020 24.770 ;
  LAYER VI3 ;
  RECT 1374.820 24.170 1375.020 24.370 ;
  LAYER VI3 ;
  RECT 1374.420 24.570 1374.620 24.770 ;
  LAYER VI3 ;
  RECT 1374.420 24.170 1374.620 24.370 ;
  LAYER VI2 ;
  RECT 1374.360 24.170 1375.220 25.170 ;
  LAYER VI2 ;
  RECT 1374.820 24.570 1375.020 24.770 ;
  LAYER VI2 ;
  RECT 1374.820 24.170 1375.020 24.370 ;
  LAYER VI2 ;
  RECT 1374.420 24.570 1374.620 24.770 ;
  LAYER VI2 ;
  RECT 1374.420 24.170 1374.620 24.370 ;
  LAYER VI3 ;
  RECT 1374.360 36.320 1375.220 37.320 ;
  LAYER VI3 ;
  RECT 1374.820 36.720 1375.020 36.920 ;
  LAYER VI3 ;
  RECT 1374.820 36.320 1375.020 36.520 ;
  LAYER VI3 ;
  RECT 1374.420 36.720 1374.620 36.920 ;
  LAYER VI3 ;
  RECT 1374.420 36.320 1374.620 36.520 ;
  LAYER VI2 ;
  RECT 1374.360 36.320 1375.220 37.320 ;
  LAYER VI2 ;
  RECT 1374.820 36.720 1375.020 36.920 ;
  LAYER VI2 ;
  RECT 1374.820 36.320 1375.020 36.520 ;
  LAYER VI2 ;
  RECT 1374.420 36.720 1374.620 36.920 ;
  LAYER VI2 ;
  RECT 1374.420 36.320 1374.620 36.520 ;
  LAYER VI3 ;
  RECT 1374.360 39.480 1375.220 40.080 ;
  LAYER VI3 ;
  RECT 1374.760 39.540 1374.960 39.740 ;
  LAYER VI3 ;
  RECT 1374.360 39.540 1374.560 39.740 ;
  LAYER VI2 ;
  RECT 1374.360 39.480 1375.220 40.080 ;
  LAYER VI2 ;
  RECT 1374.760 39.540 1374.960 39.740 ;
  LAYER VI2 ;
  RECT 1374.360 39.540 1374.560 39.740 ;
  LAYER VI3 ;
  RECT 1374.360 45.560 1375.220 46.160 ;
  LAYER VI3 ;
  RECT 1374.760 45.620 1374.960 45.820 ;
  LAYER VI3 ;
  RECT 1374.360 45.620 1374.560 45.820 ;
  LAYER VI2 ;
  RECT 1374.360 45.560 1375.220 46.160 ;
  LAYER VI2 ;
  RECT 1374.760 45.620 1374.960 45.820 ;
  LAYER VI2 ;
  RECT 1374.360 45.620 1374.560 45.820 ;
  LAYER VI3 ;
  RECT 1374.360 57.100 1375.220 61.420 ;
  LAYER VI3 ;
  RECT 1374.820 61.100 1375.020 61.300 ;
  LAYER VI3 ;
  RECT 1374.820 60.700 1375.020 60.900 ;
  LAYER VI3 ;
  RECT 1374.820 60.300 1375.020 60.500 ;
  LAYER VI3 ;
  RECT 1374.820 59.900 1375.020 60.100 ;
  LAYER VI3 ;
  RECT 1374.820 59.500 1375.020 59.700 ;
  LAYER VI3 ;
  RECT 1374.820 59.100 1375.020 59.300 ;
  LAYER VI3 ;
  RECT 1374.820 58.700 1375.020 58.900 ;
  LAYER VI3 ;
  RECT 1374.820 58.300 1375.020 58.500 ;
  LAYER VI3 ;
  RECT 1374.820 57.900 1375.020 58.100 ;
  LAYER VI3 ;
  RECT 1374.820 57.500 1375.020 57.700 ;
  LAYER VI3 ;
  RECT 1374.820 57.100 1375.020 57.300 ;
  LAYER VI3 ;
  RECT 1374.420 61.100 1374.620 61.300 ;
  LAYER VI3 ;
  RECT 1374.420 60.700 1374.620 60.900 ;
  LAYER VI3 ;
  RECT 1374.420 60.300 1374.620 60.500 ;
  LAYER VI3 ;
  RECT 1374.420 59.900 1374.620 60.100 ;
  LAYER VI3 ;
  RECT 1374.420 59.500 1374.620 59.700 ;
  LAYER VI3 ;
  RECT 1374.420 59.100 1374.620 59.300 ;
  LAYER VI3 ;
  RECT 1374.420 58.700 1374.620 58.900 ;
  LAYER VI3 ;
  RECT 1374.420 58.300 1374.620 58.500 ;
  LAYER VI3 ;
  RECT 1374.420 57.900 1374.620 58.100 ;
  LAYER VI3 ;
  RECT 1374.420 57.500 1374.620 57.700 ;
  LAYER VI3 ;
  RECT 1374.420 57.100 1374.620 57.300 ;
  LAYER VI2 ;
  RECT 1374.360 57.100 1375.220 61.420 ;
  LAYER VI2 ;
  RECT 1374.820 61.100 1375.020 61.300 ;
  LAYER VI2 ;
  RECT 1374.820 60.700 1375.020 60.900 ;
  LAYER VI2 ;
  RECT 1374.820 60.300 1375.020 60.500 ;
  LAYER VI2 ;
  RECT 1374.820 59.900 1375.020 60.100 ;
  LAYER VI2 ;
  RECT 1374.820 59.500 1375.020 59.700 ;
  LAYER VI2 ;
  RECT 1374.820 59.100 1375.020 59.300 ;
  LAYER VI2 ;
  RECT 1374.820 58.700 1375.020 58.900 ;
  LAYER VI2 ;
  RECT 1374.820 58.300 1375.020 58.500 ;
  LAYER VI2 ;
  RECT 1374.820 57.900 1375.020 58.100 ;
  LAYER VI2 ;
  RECT 1374.820 57.500 1375.020 57.700 ;
  LAYER VI2 ;
  RECT 1374.820 57.100 1375.020 57.300 ;
  LAYER VI2 ;
  RECT 1374.420 61.100 1374.620 61.300 ;
  LAYER VI2 ;
  RECT 1374.420 60.700 1374.620 60.900 ;
  LAYER VI2 ;
  RECT 1374.420 60.300 1374.620 60.500 ;
  LAYER VI2 ;
  RECT 1374.420 59.900 1374.620 60.100 ;
  LAYER VI2 ;
  RECT 1374.420 59.500 1374.620 59.700 ;
  LAYER VI2 ;
  RECT 1374.420 59.100 1374.620 59.300 ;
  LAYER VI2 ;
  RECT 1374.420 58.700 1374.620 58.900 ;
  LAYER VI2 ;
  RECT 1374.420 58.300 1374.620 58.500 ;
  LAYER VI2 ;
  RECT 1374.420 57.900 1374.620 58.100 ;
  LAYER VI2 ;
  RECT 1374.420 57.500 1374.620 57.700 ;
  LAYER VI2 ;
  RECT 1374.420 57.100 1374.620 57.300 ;
  LAYER VI3 ;
  RECT 1372.940 5.880 1374.080 6.740 ;
  LAYER VI3 ;
  RECT 1373.740 6.340 1373.940 6.540 ;
  LAYER VI3 ;
  RECT 1373.740 5.940 1373.940 6.140 ;
  LAYER VI3 ;
  RECT 1373.340 6.340 1373.540 6.540 ;
  LAYER VI3 ;
  RECT 1373.340 5.940 1373.540 6.140 ;
  LAYER VI3 ;
  RECT 1372.940 6.340 1373.140 6.540 ;
  LAYER VI3 ;
  RECT 1372.940 5.940 1373.140 6.140 ;
  LAYER VI3 ;
  RECT 719.460 5.880 727.460 6.740 ;
  LAYER VI3 ;
  RECT 727.060 6.340 727.260 6.540 ;
  LAYER VI3 ;
  RECT 727.060 5.940 727.260 6.140 ;
  LAYER VI3 ;
  RECT 726.660 6.340 726.860 6.540 ;
  LAYER VI3 ;
  RECT 726.660 5.940 726.860 6.140 ;
  LAYER VI3 ;
  RECT 726.260 6.340 726.460 6.540 ;
  LAYER VI3 ;
  RECT 726.260 5.940 726.460 6.140 ;
  LAYER VI3 ;
  RECT 725.860 6.340 726.060 6.540 ;
  LAYER VI3 ;
  RECT 725.860 5.940 726.060 6.140 ;
  LAYER VI3 ;
  RECT 725.460 6.340 725.660 6.540 ;
  LAYER VI3 ;
  RECT 725.460 5.940 725.660 6.140 ;
  LAYER VI3 ;
  RECT 725.060 6.340 725.260 6.540 ;
  LAYER VI3 ;
  RECT 725.060 5.940 725.260 6.140 ;
  LAYER VI3 ;
  RECT 724.660 6.340 724.860 6.540 ;
  LAYER VI3 ;
  RECT 724.660 5.940 724.860 6.140 ;
  LAYER VI3 ;
  RECT 724.260 6.340 724.460 6.540 ;
  LAYER VI3 ;
  RECT 724.260 5.940 724.460 6.140 ;
  LAYER VI3 ;
  RECT 723.860 6.340 724.060 6.540 ;
  LAYER VI3 ;
  RECT 723.860 5.940 724.060 6.140 ;
  LAYER VI3 ;
  RECT 723.460 6.340 723.660 6.540 ;
  LAYER VI3 ;
  RECT 723.460 5.940 723.660 6.140 ;
  LAYER VI3 ;
  RECT 723.060 6.340 723.260 6.540 ;
  LAYER VI3 ;
  RECT 723.060 5.940 723.260 6.140 ;
  LAYER VI3 ;
  RECT 722.660 6.340 722.860 6.540 ;
  LAYER VI3 ;
  RECT 722.660 5.940 722.860 6.140 ;
  LAYER VI3 ;
  RECT 722.260 6.340 722.460 6.540 ;
  LAYER VI3 ;
  RECT 722.260 5.940 722.460 6.140 ;
  LAYER VI3 ;
  RECT 721.860 6.340 722.060 6.540 ;
  LAYER VI3 ;
  RECT 721.860 5.940 722.060 6.140 ;
  LAYER VI3 ;
  RECT 721.460 6.340 721.660 6.540 ;
  LAYER VI3 ;
  RECT 721.460 5.940 721.660 6.140 ;
  LAYER VI3 ;
  RECT 721.060 6.340 721.260 6.540 ;
  LAYER VI3 ;
  RECT 721.060 5.940 721.260 6.140 ;
  LAYER VI3 ;
  RECT 720.660 6.340 720.860 6.540 ;
  LAYER VI3 ;
  RECT 720.660 5.940 720.860 6.140 ;
  LAYER VI3 ;
  RECT 720.260 6.340 720.460 6.540 ;
  LAYER VI3 ;
  RECT 720.260 5.940 720.460 6.140 ;
  LAYER VI3 ;
  RECT 719.860 6.340 720.060 6.540 ;
  LAYER VI3 ;
  RECT 719.860 5.940 720.060 6.140 ;
  LAYER VI3 ;
  RECT 719.460 6.340 719.660 6.540 ;
  LAYER VI3 ;
  RECT 719.460 5.940 719.660 6.140 ;
  LAYER VI3 ;
  RECT 739.300 5.880 747.300 6.740 ;
  LAYER VI3 ;
  RECT 746.900 6.340 747.100 6.540 ;
  LAYER VI3 ;
  RECT 746.900 5.940 747.100 6.140 ;
  LAYER VI3 ;
  RECT 746.500 6.340 746.700 6.540 ;
  LAYER VI3 ;
  RECT 746.500 5.940 746.700 6.140 ;
  LAYER VI3 ;
  RECT 746.100 6.340 746.300 6.540 ;
  LAYER VI3 ;
  RECT 746.100 5.940 746.300 6.140 ;
  LAYER VI3 ;
  RECT 745.700 6.340 745.900 6.540 ;
  LAYER VI3 ;
  RECT 745.700 5.940 745.900 6.140 ;
  LAYER VI3 ;
  RECT 745.300 6.340 745.500 6.540 ;
  LAYER VI3 ;
  RECT 745.300 5.940 745.500 6.140 ;
  LAYER VI3 ;
  RECT 744.900 6.340 745.100 6.540 ;
  LAYER VI3 ;
  RECT 744.900 5.940 745.100 6.140 ;
  LAYER VI3 ;
  RECT 744.500 6.340 744.700 6.540 ;
  LAYER VI3 ;
  RECT 744.500 5.940 744.700 6.140 ;
  LAYER VI3 ;
  RECT 744.100 6.340 744.300 6.540 ;
  LAYER VI3 ;
  RECT 744.100 5.940 744.300 6.140 ;
  LAYER VI3 ;
  RECT 743.700 6.340 743.900 6.540 ;
  LAYER VI3 ;
  RECT 743.700 5.940 743.900 6.140 ;
  LAYER VI3 ;
  RECT 743.300 6.340 743.500 6.540 ;
  LAYER VI3 ;
  RECT 743.300 5.940 743.500 6.140 ;
  LAYER VI3 ;
  RECT 742.900 6.340 743.100 6.540 ;
  LAYER VI3 ;
  RECT 742.900 5.940 743.100 6.140 ;
  LAYER VI3 ;
  RECT 742.500 6.340 742.700 6.540 ;
  LAYER VI3 ;
  RECT 742.500 5.940 742.700 6.140 ;
  LAYER VI3 ;
  RECT 742.100 6.340 742.300 6.540 ;
  LAYER VI3 ;
  RECT 742.100 5.940 742.300 6.140 ;
  LAYER VI3 ;
  RECT 741.700 6.340 741.900 6.540 ;
  LAYER VI3 ;
  RECT 741.700 5.940 741.900 6.140 ;
  LAYER VI3 ;
  RECT 741.300 6.340 741.500 6.540 ;
  LAYER VI3 ;
  RECT 741.300 5.940 741.500 6.140 ;
  LAYER VI3 ;
  RECT 740.900 6.340 741.100 6.540 ;
  LAYER VI3 ;
  RECT 740.900 5.940 741.100 6.140 ;
  LAYER VI3 ;
  RECT 740.500 6.340 740.700 6.540 ;
  LAYER VI3 ;
  RECT 740.500 5.940 740.700 6.140 ;
  LAYER VI3 ;
  RECT 740.100 6.340 740.300 6.540 ;
  LAYER VI3 ;
  RECT 740.100 5.940 740.300 6.140 ;
  LAYER VI3 ;
  RECT 739.700 6.340 739.900 6.540 ;
  LAYER VI3 ;
  RECT 739.700 5.940 739.900 6.140 ;
  LAYER VI3 ;
  RECT 739.300 6.340 739.500 6.540 ;
  LAYER VI3 ;
  RECT 739.300 5.940 739.500 6.140 ;
  LAYER VI3 ;
  RECT 760.380 5.880 768.380 6.740 ;
  LAYER VI3 ;
  RECT 767.980 6.340 768.180 6.540 ;
  LAYER VI3 ;
  RECT 767.980 5.940 768.180 6.140 ;
  LAYER VI3 ;
  RECT 767.580 6.340 767.780 6.540 ;
  LAYER VI3 ;
  RECT 767.580 5.940 767.780 6.140 ;
  LAYER VI3 ;
  RECT 767.180 6.340 767.380 6.540 ;
  LAYER VI3 ;
  RECT 767.180 5.940 767.380 6.140 ;
  LAYER VI3 ;
  RECT 766.780 6.340 766.980 6.540 ;
  LAYER VI3 ;
  RECT 766.780 5.940 766.980 6.140 ;
  LAYER VI3 ;
  RECT 766.380 6.340 766.580 6.540 ;
  LAYER VI3 ;
  RECT 766.380 5.940 766.580 6.140 ;
  LAYER VI3 ;
  RECT 765.980 6.340 766.180 6.540 ;
  LAYER VI3 ;
  RECT 765.980 5.940 766.180 6.140 ;
  LAYER VI3 ;
  RECT 765.580 6.340 765.780 6.540 ;
  LAYER VI3 ;
  RECT 765.580 5.940 765.780 6.140 ;
  LAYER VI3 ;
  RECT 765.180 6.340 765.380 6.540 ;
  LAYER VI3 ;
  RECT 765.180 5.940 765.380 6.140 ;
  LAYER VI3 ;
  RECT 764.780 6.340 764.980 6.540 ;
  LAYER VI3 ;
  RECT 764.780 5.940 764.980 6.140 ;
  LAYER VI3 ;
  RECT 764.380 6.340 764.580 6.540 ;
  LAYER VI3 ;
  RECT 764.380 5.940 764.580 6.140 ;
  LAYER VI3 ;
  RECT 763.980 6.340 764.180 6.540 ;
  LAYER VI3 ;
  RECT 763.980 5.940 764.180 6.140 ;
  LAYER VI3 ;
  RECT 763.580 6.340 763.780 6.540 ;
  LAYER VI3 ;
  RECT 763.580 5.940 763.780 6.140 ;
  LAYER VI3 ;
  RECT 763.180 6.340 763.380 6.540 ;
  LAYER VI3 ;
  RECT 763.180 5.940 763.380 6.140 ;
  LAYER VI3 ;
  RECT 762.780 6.340 762.980 6.540 ;
  LAYER VI3 ;
  RECT 762.780 5.940 762.980 6.140 ;
  LAYER VI3 ;
  RECT 762.380 6.340 762.580 6.540 ;
  LAYER VI3 ;
  RECT 762.380 5.940 762.580 6.140 ;
  LAYER VI3 ;
  RECT 761.980 6.340 762.180 6.540 ;
  LAYER VI3 ;
  RECT 761.980 5.940 762.180 6.140 ;
  LAYER VI3 ;
  RECT 761.580 6.340 761.780 6.540 ;
  LAYER VI3 ;
  RECT 761.580 5.940 761.780 6.140 ;
  LAYER VI3 ;
  RECT 761.180 6.340 761.380 6.540 ;
  LAYER VI3 ;
  RECT 761.180 5.940 761.380 6.140 ;
  LAYER VI3 ;
  RECT 760.780 6.340 760.980 6.540 ;
  LAYER VI3 ;
  RECT 760.780 5.940 760.980 6.140 ;
  LAYER VI3 ;
  RECT 760.380 6.340 760.580 6.540 ;
  LAYER VI3 ;
  RECT 760.380 5.940 760.580 6.140 ;
  LAYER VI3 ;
  RECT 780.220 5.880 788.220 6.740 ;
  LAYER VI3 ;
  RECT 787.820 6.340 788.020 6.540 ;
  LAYER VI3 ;
  RECT 787.820 5.940 788.020 6.140 ;
  LAYER VI3 ;
  RECT 787.420 6.340 787.620 6.540 ;
  LAYER VI3 ;
  RECT 787.420 5.940 787.620 6.140 ;
  LAYER VI3 ;
  RECT 787.020 6.340 787.220 6.540 ;
  LAYER VI3 ;
  RECT 787.020 5.940 787.220 6.140 ;
  LAYER VI3 ;
  RECT 786.620 6.340 786.820 6.540 ;
  LAYER VI3 ;
  RECT 786.620 5.940 786.820 6.140 ;
  LAYER VI3 ;
  RECT 786.220 6.340 786.420 6.540 ;
  LAYER VI3 ;
  RECT 786.220 5.940 786.420 6.140 ;
  LAYER VI3 ;
  RECT 785.820 6.340 786.020 6.540 ;
  LAYER VI3 ;
  RECT 785.820 5.940 786.020 6.140 ;
  LAYER VI3 ;
  RECT 785.420 6.340 785.620 6.540 ;
  LAYER VI3 ;
  RECT 785.420 5.940 785.620 6.140 ;
  LAYER VI3 ;
  RECT 785.020 6.340 785.220 6.540 ;
  LAYER VI3 ;
  RECT 785.020 5.940 785.220 6.140 ;
  LAYER VI3 ;
  RECT 784.620 6.340 784.820 6.540 ;
  LAYER VI3 ;
  RECT 784.620 5.940 784.820 6.140 ;
  LAYER VI3 ;
  RECT 784.220 6.340 784.420 6.540 ;
  LAYER VI3 ;
  RECT 784.220 5.940 784.420 6.140 ;
  LAYER VI3 ;
  RECT 783.820 6.340 784.020 6.540 ;
  LAYER VI3 ;
  RECT 783.820 5.940 784.020 6.140 ;
  LAYER VI3 ;
  RECT 783.420 6.340 783.620 6.540 ;
  LAYER VI3 ;
  RECT 783.420 5.940 783.620 6.140 ;
  LAYER VI3 ;
  RECT 783.020 6.340 783.220 6.540 ;
  LAYER VI3 ;
  RECT 783.020 5.940 783.220 6.140 ;
  LAYER VI3 ;
  RECT 782.620 6.340 782.820 6.540 ;
  LAYER VI3 ;
  RECT 782.620 5.940 782.820 6.140 ;
  LAYER VI3 ;
  RECT 782.220 6.340 782.420 6.540 ;
  LAYER VI3 ;
  RECT 782.220 5.940 782.420 6.140 ;
  LAYER VI3 ;
  RECT 781.820 6.340 782.020 6.540 ;
  LAYER VI3 ;
  RECT 781.820 5.940 782.020 6.140 ;
  LAYER VI3 ;
  RECT 781.420 6.340 781.620 6.540 ;
  LAYER VI3 ;
  RECT 781.420 5.940 781.620 6.140 ;
  LAYER VI3 ;
  RECT 781.020 6.340 781.220 6.540 ;
  LAYER VI3 ;
  RECT 781.020 5.940 781.220 6.140 ;
  LAYER VI3 ;
  RECT 780.620 6.340 780.820 6.540 ;
  LAYER VI3 ;
  RECT 780.620 5.940 780.820 6.140 ;
  LAYER VI3 ;
  RECT 780.220 6.340 780.420 6.540 ;
  LAYER VI3 ;
  RECT 780.220 5.940 780.420 6.140 ;
  LAYER VI3 ;
  RECT 801.300 5.880 809.300 6.740 ;
  LAYER VI3 ;
  RECT 808.900 6.340 809.100 6.540 ;
  LAYER VI3 ;
  RECT 808.900 5.940 809.100 6.140 ;
  LAYER VI3 ;
  RECT 808.500 6.340 808.700 6.540 ;
  LAYER VI3 ;
  RECT 808.500 5.940 808.700 6.140 ;
  LAYER VI3 ;
  RECT 808.100 6.340 808.300 6.540 ;
  LAYER VI3 ;
  RECT 808.100 5.940 808.300 6.140 ;
  LAYER VI3 ;
  RECT 807.700 6.340 807.900 6.540 ;
  LAYER VI3 ;
  RECT 807.700 5.940 807.900 6.140 ;
  LAYER VI3 ;
  RECT 807.300 6.340 807.500 6.540 ;
  LAYER VI3 ;
  RECT 807.300 5.940 807.500 6.140 ;
  LAYER VI3 ;
  RECT 806.900 6.340 807.100 6.540 ;
  LAYER VI3 ;
  RECT 806.900 5.940 807.100 6.140 ;
  LAYER VI3 ;
  RECT 806.500 6.340 806.700 6.540 ;
  LAYER VI3 ;
  RECT 806.500 5.940 806.700 6.140 ;
  LAYER VI3 ;
  RECT 806.100 6.340 806.300 6.540 ;
  LAYER VI3 ;
  RECT 806.100 5.940 806.300 6.140 ;
  LAYER VI3 ;
  RECT 805.700 6.340 805.900 6.540 ;
  LAYER VI3 ;
  RECT 805.700 5.940 805.900 6.140 ;
  LAYER VI3 ;
  RECT 805.300 6.340 805.500 6.540 ;
  LAYER VI3 ;
  RECT 805.300 5.940 805.500 6.140 ;
  LAYER VI3 ;
  RECT 804.900 6.340 805.100 6.540 ;
  LAYER VI3 ;
  RECT 804.900 5.940 805.100 6.140 ;
  LAYER VI3 ;
  RECT 804.500 6.340 804.700 6.540 ;
  LAYER VI3 ;
  RECT 804.500 5.940 804.700 6.140 ;
  LAYER VI3 ;
  RECT 804.100 6.340 804.300 6.540 ;
  LAYER VI3 ;
  RECT 804.100 5.940 804.300 6.140 ;
  LAYER VI3 ;
  RECT 803.700 6.340 803.900 6.540 ;
  LAYER VI3 ;
  RECT 803.700 5.940 803.900 6.140 ;
  LAYER VI3 ;
  RECT 803.300 6.340 803.500 6.540 ;
  LAYER VI3 ;
  RECT 803.300 5.940 803.500 6.140 ;
  LAYER VI3 ;
  RECT 802.900 6.340 803.100 6.540 ;
  LAYER VI3 ;
  RECT 802.900 5.940 803.100 6.140 ;
  LAYER VI3 ;
  RECT 802.500 6.340 802.700 6.540 ;
  LAYER VI3 ;
  RECT 802.500 5.940 802.700 6.140 ;
  LAYER VI3 ;
  RECT 802.100 6.340 802.300 6.540 ;
  LAYER VI3 ;
  RECT 802.100 5.940 802.300 6.140 ;
  LAYER VI3 ;
  RECT 801.700 6.340 801.900 6.540 ;
  LAYER VI3 ;
  RECT 801.700 5.940 801.900 6.140 ;
  LAYER VI3 ;
  RECT 801.300 6.340 801.500 6.540 ;
  LAYER VI3 ;
  RECT 801.300 5.940 801.500 6.140 ;
  LAYER VI3 ;
  RECT 821.140 5.880 829.140 6.740 ;
  LAYER VI3 ;
  RECT 828.740 6.340 828.940 6.540 ;
  LAYER VI3 ;
  RECT 828.740 5.940 828.940 6.140 ;
  LAYER VI3 ;
  RECT 828.340 6.340 828.540 6.540 ;
  LAYER VI3 ;
  RECT 828.340 5.940 828.540 6.140 ;
  LAYER VI3 ;
  RECT 827.940 6.340 828.140 6.540 ;
  LAYER VI3 ;
  RECT 827.940 5.940 828.140 6.140 ;
  LAYER VI3 ;
  RECT 827.540 6.340 827.740 6.540 ;
  LAYER VI3 ;
  RECT 827.540 5.940 827.740 6.140 ;
  LAYER VI3 ;
  RECT 827.140 6.340 827.340 6.540 ;
  LAYER VI3 ;
  RECT 827.140 5.940 827.340 6.140 ;
  LAYER VI3 ;
  RECT 826.740 6.340 826.940 6.540 ;
  LAYER VI3 ;
  RECT 826.740 5.940 826.940 6.140 ;
  LAYER VI3 ;
  RECT 826.340 6.340 826.540 6.540 ;
  LAYER VI3 ;
  RECT 826.340 5.940 826.540 6.140 ;
  LAYER VI3 ;
  RECT 825.940 6.340 826.140 6.540 ;
  LAYER VI3 ;
  RECT 825.940 5.940 826.140 6.140 ;
  LAYER VI3 ;
  RECT 825.540 6.340 825.740 6.540 ;
  LAYER VI3 ;
  RECT 825.540 5.940 825.740 6.140 ;
  LAYER VI3 ;
  RECT 825.140 6.340 825.340 6.540 ;
  LAYER VI3 ;
  RECT 825.140 5.940 825.340 6.140 ;
  LAYER VI3 ;
  RECT 824.740 6.340 824.940 6.540 ;
  LAYER VI3 ;
  RECT 824.740 5.940 824.940 6.140 ;
  LAYER VI3 ;
  RECT 824.340 6.340 824.540 6.540 ;
  LAYER VI3 ;
  RECT 824.340 5.940 824.540 6.140 ;
  LAYER VI3 ;
  RECT 823.940 6.340 824.140 6.540 ;
  LAYER VI3 ;
  RECT 823.940 5.940 824.140 6.140 ;
  LAYER VI3 ;
  RECT 823.540 6.340 823.740 6.540 ;
  LAYER VI3 ;
  RECT 823.540 5.940 823.740 6.140 ;
  LAYER VI3 ;
  RECT 823.140 6.340 823.340 6.540 ;
  LAYER VI3 ;
  RECT 823.140 5.940 823.340 6.140 ;
  LAYER VI3 ;
  RECT 822.740 6.340 822.940 6.540 ;
  LAYER VI3 ;
  RECT 822.740 5.940 822.940 6.140 ;
  LAYER VI3 ;
  RECT 822.340 6.340 822.540 6.540 ;
  LAYER VI3 ;
  RECT 822.340 5.940 822.540 6.140 ;
  LAYER VI3 ;
  RECT 821.940 6.340 822.140 6.540 ;
  LAYER VI3 ;
  RECT 821.940 5.940 822.140 6.140 ;
  LAYER VI3 ;
  RECT 821.540 6.340 821.740 6.540 ;
  LAYER VI3 ;
  RECT 821.540 5.940 821.740 6.140 ;
  LAYER VI3 ;
  RECT 821.140 6.340 821.340 6.540 ;
  LAYER VI3 ;
  RECT 821.140 5.940 821.340 6.140 ;
  LAYER VI3 ;
  RECT 842.220 5.880 850.220 6.740 ;
  LAYER VI3 ;
  RECT 849.820 6.340 850.020 6.540 ;
  LAYER VI3 ;
  RECT 849.820 5.940 850.020 6.140 ;
  LAYER VI3 ;
  RECT 849.420 6.340 849.620 6.540 ;
  LAYER VI3 ;
  RECT 849.420 5.940 849.620 6.140 ;
  LAYER VI3 ;
  RECT 849.020 6.340 849.220 6.540 ;
  LAYER VI3 ;
  RECT 849.020 5.940 849.220 6.140 ;
  LAYER VI3 ;
  RECT 848.620 6.340 848.820 6.540 ;
  LAYER VI3 ;
  RECT 848.620 5.940 848.820 6.140 ;
  LAYER VI3 ;
  RECT 848.220 6.340 848.420 6.540 ;
  LAYER VI3 ;
  RECT 848.220 5.940 848.420 6.140 ;
  LAYER VI3 ;
  RECT 847.820 6.340 848.020 6.540 ;
  LAYER VI3 ;
  RECT 847.820 5.940 848.020 6.140 ;
  LAYER VI3 ;
  RECT 847.420 6.340 847.620 6.540 ;
  LAYER VI3 ;
  RECT 847.420 5.940 847.620 6.140 ;
  LAYER VI3 ;
  RECT 847.020 6.340 847.220 6.540 ;
  LAYER VI3 ;
  RECT 847.020 5.940 847.220 6.140 ;
  LAYER VI3 ;
  RECT 846.620 6.340 846.820 6.540 ;
  LAYER VI3 ;
  RECT 846.620 5.940 846.820 6.140 ;
  LAYER VI3 ;
  RECT 846.220 6.340 846.420 6.540 ;
  LAYER VI3 ;
  RECT 846.220 5.940 846.420 6.140 ;
  LAYER VI3 ;
  RECT 845.820 6.340 846.020 6.540 ;
  LAYER VI3 ;
  RECT 845.820 5.940 846.020 6.140 ;
  LAYER VI3 ;
  RECT 845.420 6.340 845.620 6.540 ;
  LAYER VI3 ;
  RECT 845.420 5.940 845.620 6.140 ;
  LAYER VI3 ;
  RECT 845.020 6.340 845.220 6.540 ;
  LAYER VI3 ;
  RECT 845.020 5.940 845.220 6.140 ;
  LAYER VI3 ;
  RECT 844.620 6.340 844.820 6.540 ;
  LAYER VI3 ;
  RECT 844.620 5.940 844.820 6.140 ;
  LAYER VI3 ;
  RECT 844.220 6.340 844.420 6.540 ;
  LAYER VI3 ;
  RECT 844.220 5.940 844.420 6.140 ;
  LAYER VI3 ;
  RECT 843.820 6.340 844.020 6.540 ;
  LAYER VI3 ;
  RECT 843.820 5.940 844.020 6.140 ;
  LAYER VI3 ;
  RECT 843.420 6.340 843.620 6.540 ;
  LAYER VI3 ;
  RECT 843.420 5.940 843.620 6.140 ;
  LAYER VI3 ;
  RECT 843.020 6.340 843.220 6.540 ;
  LAYER VI3 ;
  RECT 843.020 5.940 843.220 6.140 ;
  LAYER VI3 ;
  RECT 842.620 6.340 842.820 6.540 ;
  LAYER VI3 ;
  RECT 842.620 5.940 842.820 6.140 ;
  LAYER VI3 ;
  RECT 842.220 6.340 842.420 6.540 ;
  LAYER VI3 ;
  RECT 842.220 5.940 842.420 6.140 ;
  LAYER VI3 ;
  RECT 862.060 5.880 870.060 6.740 ;
  LAYER VI3 ;
  RECT 869.660 6.340 869.860 6.540 ;
  LAYER VI3 ;
  RECT 869.660 5.940 869.860 6.140 ;
  LAYER VI3 ;
  RECT 869.260 6.340 869.460 6.540 ;
  LAYER VI3 ;
  RECT 869.260 5.940 869.460 6.140 ;
  LAYER VI3 ;
  RECT 868.860 6.340 869.060 6.540 ;
  LAYER VI3 ;
  RECT 868.860 5.940 869.060 6.140 ;
  LAYER VI3 ;
  RECT 868.460 6.340 868.660 6.540 ;
  LAYER VI3 ;
  RECT 868.460 5.940 868.660 6.140 ;
  LAYER VI3 ;
  RECT 868.060 6.340 868.260 6.540 ;
  LAYER VI3 ;
  RECT 868.060 5.940 868.260 6.140 ;
  LAYER VI3 ;
  RECT 867.660 6.340 867.860 6.540 ;
  LAYER VI3 ;
  RECT 867.660 5.940 867.860 6.140 ;
  LAYER VI3 ;
  RECT 867.260 6.340 867.460 6.540 ;
  LAYER VI3 ;
  RECT 867.260 5.940 867.460 6.140 ;
  LAYER VI3 ;
  RECT 866.860 6.340 867.060 6.540 ;
  LAYER VI3 ;
  RECT 866.860 5.940 867.060 6.140 ;
  LAYER VI3 ;
  RECT 866.460 6.340 866.660 6.540 ;
  LAYER VI3 ;
  RECT 866.460 5.940 866.660 6.140 ;
  LAYER VI3 ;
  RECT 866.060 6.340 866.260 6.540 ;
  LAYER VI3 ;
  RECT 866.060 5.940 866.260 6.140 ;
  LAYER VI3 ;
  RECT 865.660 6.340 865.860 6.540 ;
  LAYER VI3 ;
  RECT 865.660 5.940 865.860 6.140 ;
  LAYER VI3 ;
  RECT 865.260 6.340 865.460 6.540 ;
  LAYER VI3 ;
  RECT 865.260 5.940 865.460 6.140 ;
  LAYER VI3 ;
  RECT 864.860 6.340 865.060 6.540 ;
  LAYER VI3 ;
  RECT 864.860 5.940 865.060 6.140 ;
  LAYER VI3 ;
  RECT 864.460 6.340 864.660 6.540 ;
  LAYER VI3 ;
  RECT 864.460 5.940 864.660 6.140 ;
  LAYER VI3 ;
  RECT 864.060 6.340 864.260 6.540 ;
  LAYER VI3 ;
  RECT 864.060 5.940 864.260 6.140 ;
  LAYER VI3 ;
  RECT 863.660 6.340 863.860 6.540 ;
  LAYER VI3 ;
  RECT 863.660 5.940 863.860 6.140 ;
  LAYER VI3 ;
  RECT 863.260 6.340 863.460 6.540 ;
  LAYER VI3 ;
  RECT 863.260 5.940 863.460 6.140 ;
  LAYER VI3 ;
  RECT 862.860 6.340 863.060 6.540 ;
  LAYER VI3 ;
  RECT 862.860 5.940 863.060 6.140 ;
  LAYER VI3 ;
  RECT 862.460 6.340 862.660 6.540 ;
  LAYER VI3 ;
  RECT 862.460 5.940 862.660 6.140 ;
  LAYER VI3 ;
  RECT 862.060 6.340 862.260 6.540 ;
  LAYER VI3 ;
  RECT 862.060 5.940 862.260 6.140 ;
  LAYER VI3 ;
  RECT 883.140 5.880 891.140 6.740 ;
  LAYER VI3 ;
  RECT 890.740 6.340 890.940 6.540 ;
  LAYER VI3 ;
  RECT 890.740 5.940 890.940 6.140 ;
  LAYER VI3 ;
  RECT 890.340 6.340 890.540 6.540 ;
  LAYER VI3 ;
  RECT 890.340 5.940 890.540 6.140 ;
  LAYER VI3 ;
  RECT 889.940 6.340 890.140 6.540 ;
  LAYER VI3 ;
  RECT 889.940 5.940 890.140 6.140 ;
  LAYER VI3 ;
  RECT 889.540 6.340 889.740 6.540 ;
  LAYER VI3 ;
  RECT 889.540 5.940 889.740 6.140 ;
  LAYER VI3 ;
  RECT 889.140 6.340 889.340 6.540 ;
  LAYER VI3 ;
  RECT 889.140 5.940 889.340 6.140 ;
  LAYER VI3 ;
  RECT 888.740 6.340 888.940 6.540 ;
  LAYER VI3 ;
  RECT 888.740 5.940 888.940 6.140 ;
  LAYER VI3 ;
  RECT 888.340 6.340 888.540 6.540 ;
  LAYER VI3 ;
  RECT 888.340 5.940 888.540 6.140 ;
  LAYER VI3 ;
  RECT 887.940 6.340 888.140 6.540 ;
  LAYER VI3 ;
  RECT 887.940 5.940 888.140 6.140 ;
  LAYER VI3 ;
  RECT 887.540 6.340 887.740 6.540 ;
  LAYER VI3 ;
  RECT 887.540 5.940 887.740 6.140 ;
  LAYER VI3 ;
  RECT 887.140 6.340 887.340 6.540 ;
  LAYER VI3 ;
  RECT 887.140 5.940 887.340 6.140 ;
  LAYER VI3 ;
  RECT 886.740 6.340 886.940 6.540 ;
  LAYER VI3 ;
  RECT 886.740 5.940 886.940 6.140 ;
  LAYER VI3 ;
  RECT 886.340 6.340 886.540 6.540 ;
  LAYER VI3 ;
  RECT 886.340 5.940 886.540 6.140 ;
  LAYER VI3 ;
  RECT 885.940 6.340 886.140 6.540 ;
  LAYER VI3 ;
  RECT 885.940 5.940 886.140 6.140 ;
  LAYER VI3 ;
  RECT 885.540 6.340 885.740 6.540 ;
  LAYER VI3 ;
  RECT 885.540 5.940 885.740 6.140 ;
  LAYER VI3 ;
  RECT 885.140 6.340 885.340 6.540 ;
  LAYER VI3 ;
  RECT 885.140 5.940 885.340 6.140 ;
  LAYER VI3 ;
  RECT 884.740 6.340 884.940 6.540 ;
  LAYER VI3 ;
  RECT 884.740 5.940 884.940 6.140 ;
  LAYER VI3 ;
  RECT 884.340 6.340 884.540 6.540 ;
  LAYER VI3 ;
  RECT 884.340 5.940 884.540 6.140 ;
  LAYER VI3 ;
  RECT 883.940 6.340 884.140 6.540 ;
  LAYER VI3 ;
  RECT 883.940 5.940 884.140 6.140 ;
  LAYER VI3 ;
  RECT 883.540 6.340 883.740 6.540 ;
  LAYER VI3 ;
  RECT 883.540 5.940 883.740 6.140 ;
  LAYER VI3 ;
  RECT 883.140 6.340 883.340 6.540 ;
  LAYER VI3 ;
  RECT 883.140 5.940 883.340 6.140 ;
  LAYER VI3 ;
  RECT 902.980 5.880 910.980 6.740 ;
  LAYER VI3 ;
  RECT 910.580 6.340 910.780 6.540 ;
  LAYER VI3 ;
  RECT 910.580 5.940 910.780 6.140 ;
  LAYER VI3 ;
  RECT 910.180 6.340 910.380 6.540 ;
  LAYER VI3 ;
  RECT 910.180 5.940 910.380 6.140 ;
  LAYER VI3 ;
  RECT 909.780 6.340 909.980 6.540 ;
  LAYER VI3 ;
  RECT 909.780 5.940 909.980 6.140 ;
  LAYER VI3 ;
  RECT 909.380 6.340 909.580 6.540 ;
  LAYER VI3 ;
  RECT 909.380 5.940 909.580 6.140 ;
  LAYER VI3 ;
  RECT 908.980 6.340 909.180 6.540 ;
  LAYER VI3 ;
  RECT 908.980 5.940 909.180 6.140 ;
  LAYER VI3 ;
  RECT 908.580 6.340 908.780 6.540 ;
  LAYER VI3 ;
  RECT 908.580 5.940 908.780 6.140 ;
  LAYER VI3 ;
  RECT 908.180 6.340 908.380 6.540 ;
  LAYER VI3 ;
  RECT 908.180 5.940 908.380 6.140 ;
  LAYER VI3 ;
  RECT 907.780 6.340 907.980 6.540 ;
  LAYER VI3 ;
  RECT 907.780 5.940 907.980 6.140 ;
  LAYER VI3 ;
  RECT 907.380 6.340 907.580 6.540 ;
  LAYER VI3 ;
  RECT 907.380 5.940 907.580 6.140 ;
  LAYER VI3 ;
  RECT 906.980 6.340 907.180 6.540 ;
  LAYER VI3 ;
  RECT 906.980 5.940 907.180 6.140 ;
  LAYER VI3 ;
  RECT 906.580 6.340 906.780 6.540 ;
  LAYER VI3 ;
  RECT 906.580 5.940 906.780 6.140 ;
  LAYER VI3 ;
  RECT 906.180 6.340 906.380 6.540 ;
  LAYER VI3 ;
  RECT 906.180 5.940 906.380 6.140 ;
  LAYER VI3 ;
  RECT 905.780 6.340 905.980 6.540 ;
  LAYER VI3 ;
  RECT 905.780 5.940 905.980 6.140 ;
  LAYER VI3 ;
  RECT 905.380 6.340 905.580 6.540 ;
  LAYER VI3 ;
  RECT 905.380 5.940 905.580 6.140 ;
  LAYER VI3 ;
  RECT 904.980 6.340 905.180 6.540 ;
  LAYER VI3 ;
  RECT 904.980 5.940 905.180 6.140 ;
  LAYER VI3 ;
  RECT 904.580 6.340 904.780 6.540 ;
  LAYER VI3 ;
  RECT 904.580 5.940 904.780 6.140 ;
  LAYER VI3 ;
  RECT 904.180 6.340 904.380 6.540 ;
  LAYER VI3 ;
  RECT 904.180 5.940 904.380 6.140 ;
  LAYER VI3 ;
  RECT 903.780 6.340 903.980 6.540 ;
  LAYER VI3 ;
  RECT 903.780 5.940 903.980 6.140 ;
  LAYER VI3 ;
  RECT 903.380 6.340 903.580 6.540 ;
  LAYER VI3 ;
  RECT 903.380 5.940 903.580 6.140 ;
  LAYER VI3 ;
  RECT 902.980 6.340 903.180 6.540 ;
  LAYER VI3 ;
  RECT 902.980 5.940 903.180 6.140 ;
  LAYER VI3 ;
  RECT 924.060 5.880 932.060 6.740 ;
  LAYER VI3 ;
  RECT 931.660 6.340 931.860 6.540 ;
  LAYER VI3 ;
  RECT 931.660 5.940 931.860 6.140 ;
  LAYER VI3 ;
  RECT 931.260 6.340 931.460 6.540 ;
  LAYER VI3 ;
  RECT 931.260 5.940 931.460 6.140 ;
  LAYER VI3 ;
  RECT 930.860 6.340 931.060 6.540 ;
  LAYER VI3 ;
  RECT 930.860 5.940 931.060 6.140 ;
  LAYER VI3 ;
  RECT 930.460 6.340 930.660 6.540 ;
  LAYER VI3 ;
  RECT 930.460 5.940 930.660 6.140 ;
  LAYER VI3 ;
  RECT 930.060 6.340 930.260 6.540 ;
  LAYER VI3 ;
  RECT 930.060 5.940 930.260 6.140 ;
  LAYER VI3 ;
  RECT 929.660 6.340 929.860 6.540 ;
  LAYER VI3 ;
  RECT 929.660 5.940 929.860 6.140 ;
  LAYER VI3 ;
  RECT 929.260 6.340 929.460 6.540 ;
  LAYER VI3 ;
  RECT 929.260 5.940 929.460 6.140 ;
  LAYER VI3 ;
  RECT 928.860 6.340 929.060 6.540 ;
  LAYER VI3 ;
  RECT 928.860 5.940 929.060 6.140 ;
  LAYER VI3 ;
  RECT 928.460 6.340 928.660 6.540 ;
  LAYER VI3 ;
  RECT 928.460 5.940 928.660 6.140 ;
  LAYER VI3 ;
  RECT 928.060 6.340 928.260 6.540 ;
  LAYER VI3 ;
  RECT 928.060 5.940 928.260 6.140 ;
  LAYER VI3 ;
  RECT 927.660 6.340 927.860 6.540 ;
  LAYER VI3 ;
  RECT 927.660 5.940 927.860 6.140 ;
  LAYER VI3 ;
  RECT 927.260 6.340 927.460 6.540 ;
  LAYER VI3 ;
  RECT 927.260 5.940 927.460 6.140 ;
  LAYER VI3 ;
  RECT 926.860 6.340 927.060 6.540 ;
  LAYER VI3 ;
  RECT 926.860 5.940 927.060 6.140 ;
  LAYER VI3 ;
  RECT 926.460 6.340 926.660 6.540 ;
  LAYER VI3 ;
  RECT 926.460 5.940 926.660 6.140 ;
  LAYER VI3 ;
  RECT 926.060 6.340 926.260 6.540 ;
  LAYER VI3 ;
  RECT 926.060 5.940 926.260 6.140 ;
  LAYER VI3 ;
  RECT 925.660 6.340 925.860 6.540 ;
  LAYER VI3 ;
  RECT 925.660 5.940 925.860 6.140 ;
  LAYER VI3 ;
  RECT 925.260 6.340 925.460 6.540 ;
  LAYER VI3 ;
  RECT 925.260 5.940 925.460 6.140 ;
  LAYER VI3 ;
  RECT 924.860 6.340 925.060 6.540 ;
  LAYER VI3 ;
  RECT 924.860 5.940 925.060 6.140 ;
  LAYER VI3 ;
  RECT 924.460 6.340 924.660 6.540 ;
  LAYER VI3 ;
  RECT 924.460 5.940 924.660 6.140 ;
  LAYER VI3 ;
  RECT 924.060 6.340 924.260 6.540 ;
  LAYER VI3 ;
  RECT 924.060 5.940 924.260 6.140 ;
  LAYER VI3 ;
  RECT 943.900 5.880 951.900 6.740 ;
  LAYER VI3 ;
  RECT 951.500 6.340 951.700 6.540 ;
  LAYER VI3 ;
  RECT 951.500 5.940 951.700 6.140 ;
  LAYER VI3 ;
  RECT 951.100 6.340 951.300 6.540 ;
  LAYER VI3 ;
  RECT 951.100 5.940 951.300 6.140 ;
  LAYER VI3 ;
  RECT 950.700 6.340 950.900 6.540 ;
  LAYER VI3 ;
  RECT 950.700 5.940 950.900 6.140 ;
  LAYER VI3 ;
  RECT 950.300 6.340 950.500 6.540 ;
  LAYER VI3 ;
  RECT 950.300 5.940 950.500 6.140 ;
  LAYER VI3 ;
  RECT 949.900 6.340 950.100 6.540 ;
  LAYER VI3 ;
  RECT 949.900 5.940 950.100 6.140 ;
  LAYER VI3 ;
  RECT 949.500 6.340 949.700 6.540 ;
  LAYER VI3 ;
  RECT 949.500 5.940 949.700 6.140 ;
  LAYER VI3 ;
  RECT 949.100 6.340 949.300 6.540 ;
  LAYER VI3 ;
  RECT 949.100 5.940 949.300 6.140 ;
  LAYER VI3 ;
  RECT 948.700 6.340 948.900 6.540 ;
  LAYER VI3 ;
  RECT 948.700 5.940 948.900 6.140 ;
  LAYER VI3 ;
  RECT 948.300 6.340 948.500 6.540 ;
  LAYER VI3 ;
  RECT 948.300 5.940 948.500 6.140 ;
  LAYER VI3 ;
  RECT 947.900 6.340 948.100 6.540 ;
  LAYER VI3 ;
  RECT 947.900 5.940 948.100 6.140 ;
  LAYER VI3 ;
  RECT 947.500 6.340 947.700 6.540 ;
  LAYER VI3 ;
  RECT 947.500 5.940 947.700 6.140 ;
  LAYER VI3 ;
  RECT 947.100 6.340 947.300 6.540 ;
  LAYER VI3 ;
  RECT 947.100 5.940 947.300 6.140 ;
  LAYER VI3 ;
  RECT 946.700 6.340 946.900 6.540 ;
  LAYER VI3 ;
  RECT 946.700 5.940 946.900 6.140 ;
  LAYER VI3 ;
  RECT 946.300 6.340 946.500 6.540 ;
  LAYER VI3 ;
  RECT 946.300 5.940 946.500 6.140 ;
  LAYER VI3 ;
  RECT 945.900 6.340 946.100 6.540 ;
  LAYER VI3 ;
  RECT 945.900 5.940 946.100 6.140 ;
  LAYER VI3 ;
  RECT 945.500 6.340 945.700 6.540 ;
  LAYER VI3 ;
  RECT 945.500 5.940 945.700 6.140 ;
  LAYER VI3 ;
  RECT 945.100 6.340 945.300 6.540 ;
  LAYER VI3 ;
  RECT 945.100 5.940 945.300 6.140 ;
  LAYER VI3 ;
  RECT 944.700 6.340 944.900 6.540 ;
  LAYER VI3 ;
  RECT 944.700 5.940 944.900 6.140 ;
  LAYER VI3 ;
  RECT 944.300 6.340 944.500 6.540 ;
  LAYER VI3 ;
  RECT 944.300 5.940 944.500 6.140 ;
  LAYER VI3 ;
  RECT 943.900 6.340 944.100 6.540 ;
  LAYER VI3 ;
  RECT 943.900 5.940 944.100 6.140 ;
  LAYER VI3 ;
  RECT 964.980 5.880 972.980 6.740 ;
  LAYER VI3 ;
  RECT 972.580 6.340 972.780 6.540 ;
  LAYER VI3 ;
  RECT 972.580 5.940 972.780 6.140 ;
  LAYER VI3 ;
  RECT 972.180 6.340 972.380 6.540 ;
  LAYER VI3 ;
  RECT 972.180 5.940 972.380 6.140 ;
  LAYER VI3 ;
  RECT 971.780 6.340 971.980 6.540 ;
  LAYER VI3 ;
  RECT 971.780 5.940 971.980 6.140 ;
  LAYER VI3 ;
  RECT 971.380 6.340 971.580 6.540 ;
  LAYER VI3 ;
  RECT 971.380 5.940 971.580 6.140 ;
  LAYER VI3 ;
  RECT 970.980 6.340 971.180 6.540 ;
  LAYER VI3 ;
  RECT 970.980 5.940 971.180 6.140 ;
  LAYER VI3 ;
  RECT 970.580 6.340 970.780 6.540 ;
  LAYER VI3 ;
  RECT 970.580 5.940 970.780 6.140 ;
  LAYER VI3 ;
  RECT 970.180 6.340 970.380 6.540 ;
  LAYER VI3 ;
  RECT 970.180 5.940 970.380 6.140 ;
  LAYER VI3 ;
  RECT 969.780 6.340 969.980 6.540 ;
  LAYER VI3 ;
  RECT 969.780 5.940 969.980 6.140 ;
  LAYER VI3 ;
  RECT 969.380 6.340 969.580 6.540 ;
  LAYER VI3 ;
  RECT 969.380 5.940 969.580 6.140 ;
  LAYER VI3 ;
  RECT 968.980 6.340 969.180 6.540 ;
  LAYER VI3 ;
  RECT 968.980 5.940 969.180 6.140 ;
  LAYER VI3 ;
  RECT 968.580 6.340 968.780 6.540 ;
  LAYER VI3 ;
  RECT 968.580 5.940 968.780 6.140 ;
  LAYER VI3 ;
  RECT 968.180 6.340 968.380 6.540 ;
  LAYER VI3 ;
  RECT 968.180 5.940 968.380 6.140 ;
  LAYER VI3 ;
  RECT 967.780 6.340 967.980 6.540 ;
  LAYER VI3 ;
  RECT 967.780 5.940 967.980 6.140 ;
  LAYER VI3 ;
  RECT 967.380 6.340 967.580 6.540 ;
  LAYER VI3 ;
  RECT 967.380 5.940 967.580 6.140 ;
  LAYER VI3 ;
  RECT 966.980 6.340 967.180 6.540 ;
  LAYER VI3 ;
  RECT 966.980 5.940 967.180 6.140 ;
  LAYER VI3 ;
  RECT 966.580 6.340 966.780 6.540 ;
  LAYER VI3 ;
  RECT 966.580 5.940 966.780 6.140 ;
  LAYER VI3 ;
  RECT 966.180 6.340 966.380 6.540 ;
  LAYER VI3 ;
  RECT 966.180 5.940 966.380 6.140 ;
  LAYER VI3 ;
  RECT 965.780 6.340 965.980 6.540 ;
  LAYER VI3 ;
  RECT 965.780 5.940 965.980 6.140 ;
  LAYER VI3 ;
  RECT 965.380 6.340 965.580 6.540 ;
  LAYER VI3 ;
  RECT 965.380 5.940 965.580 6.140 ;
  LAYER VI3 ;
  RECT 964.980 6.340 965.180 6.540 ;
  LAYER VI3 ;
  RECT 964.980 5.940 965.180 6.140 ;
  LAYER VI3 ;
  RECT 984.820 5.880 992.820 6.740 ;
  LAYER VI3 ;
  RECT 992.420 6.340 992.620 6.540 ;
  LAYER VI3 ;
  RECT 992.420 5.940 992.620 6.140 ;
  LAYER VI3 ;
  RECT 992.020 6.340 992.220 6.540 ;
  LAYER VI3 ;
  RECT 992.020 5.940 992.220 6.140 ;
  LAYER VI3 ;
  RECT 991.620 6.340 991.820 6.540 ;
  LAYER VI3 ;
  RECT 991.620 5.940 991.820 6.140 ;
  LAYER VI3 ;
  RECT 991.220 6.340 991.420 6.540 ;
  LAYER VI3 ;
  RECT 991.220 5.940 991.420 6.140 ;
  LAYER VI3 ;
  RECT 990.820 6.340 991.020 6.540 ;
  LAYER VI3 ;
  RECT 990.820 5.940 991.020 6.140 ;
  LAYER VI3 ;
  RECT 990.420 6.340 990.620 6.540 ;
  LAYER VI3 ;
  RECT 990.420 5.940 990.620 6.140 ;
  LAYER VI3 ;
  RECT 990.020 6.340 990.220 6.540 ;
  LAYER VI3 ;
  RECT 990.020 5.940 990.220 6.140 ;
  LAYER VI3 ;
  RECT 989.620 6.340 989.820 6.540 ;
  LAYER VI3 ;
  RECT 989.620 5.940 989.820 6.140 ;
  LAYER VI3 ;
  RECT 989.220 6.340 989.420 6.540 ;
  LAYER VI3 ;
  RECT 989.220 5.940 989.420 6.140 ;
  LAYER VI3 ;
  RECT 988.820 6.340 989.020 6.540 ;
  LAYER VI3 ;
  RECT 988.820 5.940 989.020 6.140 ;
  LAYER VI3 ;
  RECT 988.420 6.340 988.620 6.540 ;
  LAYER VI3 ;
  RECT 988.420 5.940 988.620 6.140 ;
  LAYER VI3 ;
  RECT 988.020 6.340 988.220 6.540 ;
  LAYER VI3 ;
  RECT 988.020 5.940 988.220 6.140 ;
  LAYER VI3 ;
  RECT 987.620 6.340 987.820 6.540 ;
  LAYER VI3 ;
  RECT 987.620 5.940 987.820 6.140 ;
  LAYER VI3 ;
  RECT 987.220 6.340 987.420 6.540 ;
  LAYER VI3 ;
  RECT 987.220 5.940 987.420 6.140 ;
  LAYER VI3 ;
  RECT 986.820 6.340 987.020 6.540 ;
  LAYER VI3 ;
  RECT 986.820 5.940 987.020 6.140 ;
  LAYER VI3 ;
  RECT 986.420 6.340 986.620 6.540 ;
  LAYER VI3 ;
  RECT 986.420 5.940 986.620 6.140 ;
  LAYER VI3 ;
  RECT 986.020 6.340 986.220 6.540 ;
  LAYER VI3 ;
  RECT 986.020 5.940 986.220 6.140 ;
  LAYER VI3 ;
  RECT 985.620 6.340 985.820 6.540 ;
  LAYER VI3 ;
  RECT 985.620 5.940 985.820 6.140 ;
  LAYER VI3 ;
  RECT 985.220 6.340 985.420 6.540 ;
  LAYER VI3 ;
  RECT 985.220 5.940 985.420 6.140 ;
  LAYER VI3 ;
  RECT 984.820 6.340 985.020 6.540 ;
  LAYER VI3 ;
  RECT 984.820 5.940 985.020 6.140 ;
  LAYER VI3 ;
  RECT 1005.900 5.880 1013.900 6.740 ;
  LAYER VI3 ;
  RECT 1013.500 6.340 1013.700 6.540 ;
  LAYER VI3 ;
  RECT 1013.500 5.940 1013.700 6.140 ;
  LAYER VI3 ;
  RECT 1013.100 6.340 1013.300 6.540 ;
  LAYER VI3 ;
  RECT 1013.100 5.940 1013.300 6.140 ;
  LAYER VI3 ;
  RECT 1012.700 6.340 1012.900 6.540 ;
  LAYER VI3 ;
  RECT 1012.700 5.940 1012.900 6.140 ;
  LAYER VI3 ;
  RECT 1012.300 6.340 1012.500 6.540 ;
  LAYER VI3 ;
  RECT 1012.300 5.940 1012.500 6.140 ;
  LAYER VI3 ;
  RECT 1011.900 6.340 1012.100 6.540 ;
  LAYER VI3 ;
  RECT 1011.900 5.940 1012.100 6.140 ;
  LAYER VI3 ;
  RECT 1011.500 6.340 1011.700 6.540 ;
  LAYER VI3 ;
  RECT 1011.500 5.940 1011.700 6.140 ;
  LAYER VI3 ;
  RECT 1011.100 6.340 1011.300 6.540 ;
  LAYER VI3 ;
  RECT 1011.100 5.940 1011.300 6.140 ;
  LAYER VI3 ;
  RECT 1010.700 6.340 1010.900 6.540 ;
  LAYER VI3 ;
  RECT 1010.700 5.940 1010.900 6.140 ;
  LAYER VI3 ;
  RECT 1010.300 6.340 1010.500 6.540 ;
  LAYER VI3 ;
  RECT 1010.300 5.940 1010.500 6.140 ;
  LAYER VI3 ;
  RECT 1009.900 6.340 1010.100 6.540 ;
  LAYER VI3 ;
  RECT 1009.900 5.940 1010.100 6.140 ;
  LAYER VI3 ;
  RECT 1009.500 6.340 1009.700 6.540 ;
  LAYER VI3 ;
  RECT 1009.500 5.940 1009.700 6.140 ;
  LAYER VI3 ;
  RECT 1009.100 6.340 1009.300 6.540 ;
  LAYER VI3 ;
  RECT 1009.100 5.940 1009.300 6.140 ;
  LAYER VI3 ;
  RECT 1008.700 6.340 1008.900 6.540 ;
  LAYER VI3 ;
  RECT 1008.700 5.940 1008.900 6.140 ;
  LAYER VI3 ;
  RECT 1008.300 6.340 1008.500 6.540 ;
  LAYER VI3 ;
  RECT 1008.300 5.940 1008.500 6.140 ;
  LAYER VI3 ;
  RECT 1007.900 6.340 1008.100 6.540 ;
  LAYER VI3 ;
  RECT 1007.900 5.940 1008.100 6.140 ;
  LAYER VI3 ;
  RECT 1007.500 6.340 1007.700 6.540 ;
  LAYER VI3 ;
  RECT 1007.500 5.940 1007.700 6.140 ;
  LAYER VI3 ;
  RECT 1007.100 6.340 1007.300 6.540 ;
  LAYER VI3 ;
  RECT 1007.100 5.940 1007.300 6.140 ;
  LAYER VI3 ;
  RECT 1006.700 6.340 1006.900 6.540 ;
  LAYER VI3 ;
  RECT 1006.700 5.940 1006.900 6.140 ;
  LAYER VI3 ;
  RECT 1006.300 6.340 1006.500 6.540 ;
  LAYER VI3 ;
  RECT 1006.300 5.940 1006.500 6.140 ;
  LAYER VI3 ;
  RECT 1005.900 6.340 1006.100 6.540 ;
  LAYER VI3 ;
  RECT 1005.900 5.940 1006.100 6.140 ;
  LAYER VI3 ;
  RECT 1025.740 5.880 1033.740 6.740 ;
  LAYER VI3 ;
  RECT 1033.340 6.340 1033.540 6.540 ;
  LAYER VI3 ;
  RECT 1033.340 5.940 1033.540 6.140 ;
  LAYER VI3 ;
  RECT 1032.940 6.340 1033.140 6.540 ;
  LAYER VI3 ;
  RECT 1032.940 5.940 1033.140 6.140 ;
  LAYER VI3 ;
  RECT 1032.540 6.340 1032.740 6.540 ;
  LAYER VI3 ;
  RECT 1032.540 5.940 1032.740 6.140 ;
  LAYER VI3 ;
  RECT 1032.140 6.340 1032.340 6.540 ;
  LAYER VI3 ;
  RECT 1032.140 5.940 1032.340 6.140 ;
  LAYER VI3 ;
  RECT 1031.740 6.340 1031.940 6.540 ;
  LAYER VI3 ;
  RECT 1031.740 5.940 1031.940 6.140 ;
  LAYER VI3 ;
  RECT 1031.340 6.340 1031.540 6.540 ;
  LAYER VI3 ;
  RECT 1031.340 5.940 1031.540 6.140 ;
  LAYER VI3 ;
  RECT 1030.940 6.340 1031.140 6.540 ;
  LAYER VI3 ;
  RECT 1030.940 5.940 1031.140 6.140 ;
  LAYER VI3 ;
  RECT 1030.540 6.340 1030.740 6.540 ;
  LAYER VI3 ;
  RECT 1030.540 5.940 1030.740 6.140 ;
  LAYER VI3 ;
  RECT 1030.140 6.340 1030.340 6.540 ;
  LAYER VI3 ;
  RECT 1030.140 5.940 1030.340 6.140 ;
  LAYER VI3 ;
  RECT 1029.740 6.340 1029.940 6.540 ;
  LAYER VI3 ;
  RECT 1029.740 5.940 1029.940 6.140 ;
  LAYER VI3 ;
  RECT 1029.340 6.340 1029.540 6.540 ;
  LAYER VI3 ;
  RECT 1029.340 5.940 1029.540 6.140 ;
  LAYER VI3 ;
  RECT 1028.940 6.340 1029.140 6.540 ;
  LAYER VI3 ;
  RECT 1028.940 5.940 1029.140 6.140 ;
  LAYER VI3 ;
  RECT 1028.540 6.340 1028.740 6.540 ;
  LAYER VI3 ;
  RECT 1028.540 5.940 1028.740 6.140 ;
  LAYER VI3 ;
  RECT 1028.140 6.340 1028.340 6.540 ;
  LAYER VI3 ;
  RECT 1028.140 5.940 1028.340 6.140 ;
  LAYER VI3 ;
  RECT 1027.740 6.340 1027.940 6.540 ;
  LAYER VI3 ;
  RECT 1027.740 5.940 1027.940 6.140 ;
  LAYER VI3 ;
  RECT 1027.340 6.340 1027.540 6.540 ;
  LAYER VI3 ;
  RECT 1027.340 5.940 1027.540 6.140 ;
  LAYER VI3 ;
  RECT 1026.940 6.340 1027.140 6.540 ;
  LAYER VI3 ;
  RECT 1026.940 5.940 1027.140 6.140 ;
  LAYER VI3 ;
  RECT 1026.540 6.340 1026.740 6.540 ;
  LAYER VI3 ;
  RECT 1026.540 5.940 1026.740 6.140 ;
  LAYER VI3 ;
  RECT 1026.140 6.340 1026.340 6.540 ;
  LAYER VI3 ;
  RECT 1026.140 5.940 1026.340 6.140 ;
  LAYER VI3 ;
  RECT 1025.740 6.340 1025.940 6.540 ;
  LAYER VI3 ;
  RECT 1025.740 5.940 1025.940 6.140 ;
  LAYER VI3 ;
  RECT 1046.820 5.880 1054.820 6.740 ;
  LAYER VI3 ;
  RECT 1054.420 6.340 1054.620 6.540 ;
  LAYER VI3 ;
  RECT 1054.420 5.940 1054.620 6.140 ;
  LAYER VI3 ;
  RECT 1054.020 6.340 1054.220 6.540 ;
  LAYER VI3 ;
  RECT 1054.020 5.940 1054.220 6.140 ;
  LAYER VI3 ;
  RECT 1053.620 6.340 1053.820 6.540 ;
  LAYER VI3 ;
  RECT 1053.620 5.940 1053.820 6.140 ;
  LAYER VI3 ;
  RECT 1053.220 6.340 1053.420 6.540 ;
  LAYER VI3 ;
  RECT 1053.220 5.940 1053.420 6.140 ;
  LAYER VI3 ;
  RECT 1052.820 6.340 1053.020 6.540 ;
  LAYER VI3 ;
  RECT 1052.820 5.940 1053.020 6.140 ;
  LAYER VI3 ;
  RECT 1052.420 6.340 1052.620 6.540 ;
  LAYER VI3 ;
  RECT 1052.420 5.940 1052.620 6.140 ;
  LAYER VI3 ;
  RECT 1052.020 6.340 1052.220 6.540 ;
  LAYER VI3 ;
  RECT 1052.020 5.940 1052.220 6.140 ;
  LAYER VI3 ;
  RECT 1051.620 6.340 1051.820 6.540 ;
  LAYER VI3 ;
  RECT 1051.620 5.940 1051.820 6.140 ;
  LAYER VI3 ;
  RECT 1051.220 6.340 1051.420 6.540 ;
  LAYER VI3 ;
  RECT 1051.220 5.940 1051.420 6.140 ;
  LAYER VI3 ;
  RECT 1050.820 6.340 1051.020 6.540 ;
  LAYER VI3 ;
  RECT 1050.820 5.940 1051.020 6.140 ;
  LAYER VI3 ;
  RECT 1050.420 6.340 1050.620 6.540 ;
  LAYER VI3 ;
  RECT 1050.420 5.940 1050.620 6.140 ;
  LAYER VI3 ;
  RECT 1050.020 6.340 1050.220 6.540 ;
  LAYER VI3 ;
  RECT 1050.020 5.940 1050.220 6.140 ;
  LAYER VI3 ;
  RECT 1049.620 6.340 1049.820 6.540 ;
  LAYER VI3 ;
  RECT 1049.620 5.940 1049.820 6.140 ;
  LAYER VI3 ;
  RECT 1049.220 6.340 1049.420 6.540 ;
  LAYER VI3 ;
  RECT 1049.220 5.940 1049.420 6.140 ;
  LAYER VI3 ;
  RECT 1048.820 6.340 1049.020 6.540 ;
  LAYER VI3 ;
  RECT 1048.820 5.940 1049.020 6.140 ;
  LAYER VI3 ;
  RECT 1048.420 6.340 1048.620 6.540 ;
  LAYER VI3 ;
  RECT 1048.420 5.940 1048.620 6.140 ;
  LAYER VI3 ;
  RECT 1048.020 6.340 1048.220 6.540 ;
  LAYER VI3 ;
  RECT 1048.020 5.940 1048.220 6.140 ;
  LAYER VI3 ;
  RECT 1047.620 6.340 1047.820 6.540 ;
  LAYER VI3 ;
  RECT 1047.620 5.940 1047.820 6.140 ;
  LAYER VI3 ;
  RECT 1047.220 6.340 1047.420 6.540 ;
  LAYER VI3 ;
  RECT 1047.220 5.940 1047.420 6.140 ;
  LAYER VI3 ;
  RECT 1046.820 6.340 1047.020 6.540 ;
  LAYER VI3 ;
  RECT 1046.820 5.940 1047.020 6.140 ;
  LAYER VI3 ;
  RECT 1066.660 5.880 1074.660 6.740 ;
  LAYER VI3 ;
  RECT 1074.260 6.340 1074.460 6.540 ;
  LAYER VI3 ;
  RECT 1074.260 5.940 1074.460 6.140 ;
  LAYER VI3 ;
  RECT 1073.860 6.340 1074.060 6.540 ;
  LAYER VI3 ;
  RECT 1073.860 5.940 1074.060 6.140 ;
  LAYER VI3 ;
  RECT 1073.460 6.340 1073.660 6.540 ;
  LAYER VI3 ;
  RECT 1073.460 5.940 1073.660 6.140 ;
  LAYER VI3 ;
  RECT 1073.060 6.340 1073.260 6.540 ;
  LAYER VI3 ;
  RECT 1073.060 5.940 1073.260 6.140 ;
  LAYER VI3 ;
  RECT 1072.660 6.340 1072.860 6.540 ;
  LAYER VI3 ;
  RECT 1072.660 5.940 1072.860 6.140 ;
  LAYER VI3 ;
  RECT 1072.260 6.340 1072.460 6.540 ;
  LAYER VI3 ;
  RECT 1072.260 5.940 1072.460 6.140 ;
  LAYER VI3 ;
  RECT 1071.860 6.340 1072.060 6.540 ;
  LAYER VI3 ;
  RECT 1071.860 5.940 1072.060 6.140 ;
  LAYER VI3 ;
  RECT 1071.460 6.340 1071.660 6.540 ;
  LAYER VI3 ;
  RECT 1071.460 5.940 1071.660 6.140 ;
  LAYER VI3 ;
  RECT 1071.060 6.340 1071.260 6.540 ;
  LAYER VI3 ;
  RECT 1071.060 5.940 1071.260 6.140 ;
  LAYER VI3 ;
  RECT 1070.660 6.340 1070.860 6.540 ;
  LAYER VI3 ;
  RECT 1070.660 5.940 1070.860 6.140 ;
  LAYER VI3 ;
  RECT 1070.260 6.340 1070.460 6.540 ;
  LAYER VI3 ;
  RECT 1070.260 5.940 1070.460 6.140 ;
  LAYER VI3 ;
  RECT 1069.860 6.340 1070.060 6.540 ;
  LAYER VI3 ;
  RECT 1069.860 5.940 1070.060 6.140 ;
  LAYER VI3 ;
  RECT 1069.460 6.340 1069.660 6.540 ;
  LAYER VI3 ;
  RECT 1069.460 5.940 1069.660 6.140 ;
  LAYER VI3 ;
  RECT 1069.060 6.340 1069.260 6.540 ;
  LAYER VI3 ;
  RECT 1069.060 5.940 1069.260 6.140 ;
  LAYER VI3 ;
  RECT 1068.660 6.340 1068.860 6.540 ;
  LAYER VI3 ;
  RECT 1068.660 5.940 1068.860 6.140 ;
  LAYER VI3 ;
  RECT 1068.260 6.340 1068.460 6.540 ;
  LAYER VI3 ;
  RECT 1068.260 5.940 1068.460 6.140 ;
  LAYER VI3 ;
  RECT 1067.860 6.340 1068.060 6.540 ;
  LAYER VI3 ;
  RECT 1067.860 5.940 1068.060 6.140 ;
  LAYER VI3 ;
  RECT 1067.460 6.340 1067.660 6.540 ;
  LAYER VI3 ;
  RECT 1067.460 5.940 1067.660 6.140 ;
  LAYER VI3 ;
  RECT 1067.060 6.340 1067.260 6.540 ;
  LAYER VI3 ;
  RECT 1067.060 5.940 1067.260 6.140 ;
  LAYER VI3 ;
  RECT 1066.660 6.340 1066.860 6.540 ;
  LAYER VI3 ;
  RECT 1066.660 5.940 1066.860 6.140 ;
  LAYER VI3 ;
  RECT 1087.740 5.880 1095.740 6.740 ;
  LAYER VI3 ;
  RECT 1095.340 6.340 1095.540 6.540 ;
  LAYER VI3 ;
  RECT 1095.340 5.940 1095.540 6.140 ;
  LAYER VI3 ;
  RECT 1094.940 6.340 1095.140 6.540 ;
  LAYER VI3 ;
  RECT 1094.940 5.940 1095.140 6.140 ;
  LAYER VI3 ;
  RECT 1094.540 6.340 1094.740 6.540 ;
  LAYER VI3 ;
  RECT 1094.540 5.940 1094.740 6.140 ;
  LAYER VI3 ;
  RECT 1094.140 6.340 1094.340 6.540 ;
  LAYER VI3 ;
  RECT 1094.140 5.940 1094.340 6.140 ;
  LAYER VI3 ;
  RECT 1093.740 6.340 1093.940 6.540 ;
  LAYER VI3 ;
  RECT 1093.740 5.940 1093.940 6.140 ;
  LAYER VI3 ;
  RECT 1093.340 6.340 1093.540 6.540 ;
  LAYER VI3 ;
  RECT 1093.340 5.940 1093.540 6.140 ;
  LAYER VI3 ;
  RECT 1092.940 6.340 1093.140 6.540 ;
  LAYER VI3 ;
  RECT 1092.940 5.940 1093.140 6.140 ;
  LAYER VI3 ;
  RECT 1092.540 6.340 1092.740 6.540 ;
  LAYER VI3 ;
  RECT 1092.540 5.940 1092.740 6.140 ;
  LAYER VI3 ;
  RECT 1092.140 6.340 1092.340 6.540 ;
  LAYER VI3 ;
  RECT 1092.140 5.940 1092.340 6.140 ;
  LAYER VI3 ;
  RECT 1091.740 6.340 1091.940 6.540 ;
  LAYER VI3 ;
  RECT 1091.740 5.940 1091.940 6.140 ;
  LAYER VI3 ;
  RECT 1091.340 6.340 1091.540 6.540 ;
  LAYER VI3 ;
  RECT 1091.340 5.940 1091.540 6.140 ;
  LAYER VI3 ;
  RECT 1090.940 6.340 1091.140 6.540 ;
  LAYER VI3 ;
  RECT 1090.940 5.940 1091.140 6.140 ;
  LAYER VI3 ;
  RECT 1090.540 6.340 1090.740 6.540 ;
  LAYER VI3 ;
  RECT 1090.540 5.940 1090.740 6.140 ;
  LAYER VI3 ;
  RECT 1090.140 6.340 1090.340 6.540 ;
  LAYER VI3 ;
  RECT 1090.140 5.940 1090.340 6.140 ;
  LAYER VI3 ;
  RECT 1089.740 6.340 1089.940 6.540 ;
  LAYER VI3 ;
  RECT 1089.740 5.940 1089.940 6.140 ;
  LAYER VI3 ;
  RECT 1089.340 6.340 1089.540 6.540 ;
  LAYER VI3 ;
  RECT 1089.340 5.940 1089.540 6.140 ;
  LAYER VI3 ;
  RECT 1088.940 6.340 1089.140 6.540 ;
  LAYER VI3 ;
  RECT 1088.940 5.940 1089.140 6.140 ;
  LAYER VI3 ;
  RECT 1088.540 6.340 1088.740 6.540 ;
  LAYER VI3 ;
  RECT 1088.540 5.940 1088.740 6.140 ;
  LAYER VI3 ;
  RECT 1088.140 6.340 1088.340 6.540 ;
  LAYER VI3 ;
  RECT 1088.140 5.940 1088.340 6.140 ;
  LAYER VI3 ;
  RECT 1087.740 6.340 1087.940 6.540 ;
  LAYER VI3 ;
  RECT 1087.740 5.940 1087.940 6.140 ;
  LAYER VI3 ;
  RECT 1107.580 5.880 1115.580 6.740 ;
  LAYER VI3 ;
  RECT 1115.180 6.340 1115.380 6.540 ;
  LAYER VI3 ;
  RECT 1115.180 5.940 1115.380 6.140 ;
  LAYER VI3 ;
  RECT 1114.780 6.340 1114.980 6.540 ;
  LAYER VI3 ;
  RECT 1114.780 5.940 1114.980 6.140 ;
  LAYER VI3 ;
  RECT 1114.380 6.340 1114.580 6.540 ;
  LAYER VI3 ;
  RECT 1114.380 5.940 1114.580 6.140 ;
  LAYER VI3 ;
  RECT 1113.980 6.340 1114.180 6.540 ;
  LAYER VI3 ;
  RECT 1113.980 5.940 1114.180 6.140 ;
  LAYER VI3 ;
  RECT 1113.580 6.340 1113.780 6.540 ;
  LAYER VI3 ;
  RECT 1113.580 5.940 1113.780 6.140 ;
  LAYER VI3 ;
  RECT 1113.180 6.340 1113.380 6.540 ;
  LAYER VI3 ;
  RECT 1113.180 5.940 1113.380 6.140 ;
  LAYER VI3 ;
  RECT 1112.780 6.340 1112.980 6.540 ;
  LAYER VI3 ;
  RECT 1112.780 5.940 1112.980 6.140 ;
  LAYER VI3 ;
  RECT 1112.380 6.340 1112.580 6.540 ;
  LAYER VI3 ;
  RECT 1112.380 5.940 1112.580 6.140 ;
  LAYER VI3 ;
  RECT 1111.980 6.340 1112.180 6.540 ;
  LAYER VI3 ;
  RECT 1111.980 5.940 1112.180 6.140 ;
  LAYER VI3 ;
  RECT 1111.580 6.340 1111.780 6.540 ;
  LAYER VI3 ;
  RECT 1111.580 5.940 1111.780 6.140 ;
  LAYER VI3 ;
  RECT 1111.180 6.340 1111.380 6.540 ;
  LAYER VI3 ;
  RECT 1111.180 5.940 1111.380 6.140 ;
  LAYER VI3 ;
  RECT 1110.780 6.340 1110.980 6.540 ;
  LAYER VI3 ;
  RECT 1110.780 5.940 1110.980 6.140 ;
  LAYER VI3 ;
  RECT 1110.380 6.340 1110.580 6.540 ;
  LAYER VI3 ;
  RECT 1110.380 5.940 1110.580 6.140 ;
  LAYER VI3 ;
  RECT 1109.980 6.340 1110.180 6.540 ;
  LAYER VI3 ;
  RECT 1109.980 5.940 1110.180 6.140 ;
  LAYER VI3 ;
  RECT 1109.580 6.340 1109.780 6.540 ;
  LAYER VI3 ;
  RECT 1109.580 5.940 1109.780 6.140 ;
  LAYER VI3 ;
  RECT 1109.180 6.340 1109.380 6.540 ;
  LAYER VI3 ;
  RECT 1109.180 5.940 1109.380 6.140 ;
  LAYER VI3 ;
  RECT 1108.780 6.340 1108.980 6.540 ;
  LAYER VI3 ;
  RECT 1108.780 5.940 1108.980 6.140 ;
  LAYER VI3 ;
  RECT 1108.380 6.340 1108.580 6.540 ;
  LAYER VI3 ;
  RECT 1108.380 5.940 1108.580 6.140 ;
  LAYER VI3 ;
  RECT 1107.980 6.340 1108.180 6.540 ;
  LAYER VI3 ;
  RECT 1107.980 5.940 1108.180 6.140 ;
  LAYER VI3 ;
  RECT 1107.580 6.340 1107.780 6.540 ;
  LAYER VI3 ;
  RECT 1107.580 5.940 1107.780 6.140 ;
  LAYER VI3 ;
  RECT 1128.660 5.880 1136.660 6.740 ;
  LAYER VI3 ;
  RECT 1136.260 6.340 1136.460 6.540 ;
  LAYER VI3 ;
  RECT 1136.260 5.940 1136.460 6.140 ;
  LAYER VI3 ;
  RECT 1135.860 6.340 1136.060 6.540 ;
  LAYER VI3 ;
  RECT 1135.860 5.940 1136.060 6.140 ;
  LAYER VI3 ;
  RECT 1135.460 6.340 1135.660 6.540 ;
  LAYER VI3 ;
  RECT 1135.460 5.940 1135.660 6.140 ;
  LAYER VI3 ;
  RECT 1135.060 6.340 1135.260 6.540 ;
  LAYER VI3 ;
  RECT 1135.060 5.940 1135.260 6.140 ;
  LAYER VI3 ;
  RECT 1134.660 6.340 1134.860 6.540 ;
  LAYER VI3 ;
  RECT 1134.660 5.940 1134.860 6.140 ;
  LAYER VI3 ;
  RECT 1134.260 6.340 1134.460 6.540 ;
  LAYER VI3 ;
  RECT 1134.260 5.940 1134.460 6.140 ;
  LAYER VI3 ;
  RECT 1133.860 6.340 1134.060 6.540 ;
  LAYER VI3 ;
  RECT 1133.860 5.940 1134.060 6.140 ;
  LAYER VI3 ;
  RECT 1133.460 6.340 1133.660 6.540 ;
  LAYER VI3 ;
  RECT 1133.460 5.940 1133.660 6.140 ;
  LAYER VI3 ;
  RECT 1133.060 6.340 1133.260 6.540 ;
  LAYER VI3 ;
  RECT 1133.060 5.940 1133.260 6.140 ;
  LAYER VI3 ;
  RECT 1132.660 6.340 1132.860 6.540 ;
  LAYER VI3 ;
  RECT 1132.660 5.940 1132.860 6.140 ;
  LAYER VI3 ;
  RECT 1132.260 6.340 1132.460 6.540 ;
  LAYER VI3 ;
  RECT 1132.260 5.940 1132.460 6.140 ;
  LAYER VI3 ;
  RECT 1131.860 6.340 1132.060 6.540 ;
  LAYER VI3 ;
  RECT 1131.860 5.940 1132.060 6.140 ;
  LAYER VI3 ;
  RECT 1131.460 6.340 1131.660 6.540 ;
  LAYER VI3 ;
  RECT 1131.460 5.940 1131.660 6.140 ;
  LAYER VI3 ;
  RECT 1131.060 6.340 1131.260 6.540 ;
  LAYER VI3 ;
  RECT 1131.060 5.940 1131.260 6.140 ;
  LAYER VI3 ;
  RECT 1130.660 6.340 1130.860 6.540 ;
  LAYER VI3 ;
  RECT 1130.660 5.940 1130.860 6.140 ;
  LAYER VI3 ;
  RECT 1130.260 6.340 1130.460 6.540 ;
  LAYER VI3 ;
  RECT 1130.260 5.940 1130.460 6.140 ;
  LAYER VI3 ;
  RECT 1129.860 6.340 1130.060 6.540 ;
  LAYER VI3 ;
  RECT 1129.860 5.940 1130.060 6.140 ;
  LAYER VI3 ;
  RECT 1129.460 6.340 1129.660 6.540 ;
  LAYER VI3 ;
  RECT 1129.460 5.940 1129.660 6.140 ;
  LAYER VI3 ;
  RECT 1129.060 6.340 1129.260 6.540 ;
  LAYER VI3 ;
  RECT 1129.060 5.940 1129.260 6.140 ;
  LAYER VI3 ;
  RECT 1128.660 6.340 1128.860 6.540 ;
  LAYER VI3 ;
  RECT 1128.660 5.940 1128.860 6.140 ;
  LAYER VI3 ;
  RECT 1148.500 5.880 1156.500 6.740 ;
  LAYER VI3 ;
  RECT 1156.100 6.340 1156.300 6.540 ;
  LAYER VI3 ;
  RECT 1156.100 5.940 1156.300 6.140 ;
  LAYER VI3 ;
  RECT 1155.700 6.340 1155.900 6.540 ;
  LAYER VI3 ;
  RECT 1155.700 5.940 1155.900 6.140 ;
  LAYER VI3 ;
  RECT 1155.300 6.340 1155.500 6.540 ;
  LAYER VI3 ;
  RECT 1155.300 5.940 1155.500 6.140 ;
  LAYER VI3 ;
  RECT 1154.900 6.340 1155.100 6.540 ;
  LAYER VI3 ;
  RECT 1154.900 5.940 1155.100 6.140 ;
  LAYER VI3 ;
  RECT 1154.500 6.340 1154.700 6.540 ;
  LAYER VI3 ;
  RECT 1154.500 5.940 1154.700 6.140 ;
  LAYER VI3 ;
  RECT 1154.100 6.340 1154.300 6.540 ;
  LAYER VI3 ;
  RECT 1154.100 5.940 1154.300 6.140 ;
  LAYER VI3 ;
  RECT 1153.700 6.340 1153.900 6.540 ;
  LAYER VI3 ;
  RECT 1153.700 5.940 1153.900 6.140 ;
  LAYER VI3 ;
  RECT 1153.300 6.340 1153.500 6.540 ;
  LAYER VI3 ;
  RECT 1153.300 5.940 1153.500 6.140 ;
  LAYER VI3 ;
  RECT 1152.900 6.340 1153.100 6.540 ;
  LAYER VI3 ;
  RECT 1152.900 5.940 1153.100 6.140 ;
  LAYER VI3 ;
  RECT 1152.500 6.340 1152.700 6.540 ;
  LAYER VI3 ;
  RECT 1152.500 5.940 1152.700 6.140 ;
  LAYER VI3 ;
  RECT 1152.100 6.340 1152.300 6.540 ;
  LAYER VI3 ;
  RECT 1152.100 5.940 1152.300 6.140 ;
  LAYER VI3 ;
  RECT 1151.700 6.340 1151.900 6.540 ;
  LAYER VI3 ;
  RECT 1151.700 5.940 1151.900 6.140 ;
  LAYER VI3 ;
  RECT 1151.300 6.340 1151.500 6.540 ;
  LAYER VI3 ;
  RECT 1151.300 5.940 1151.500 6.140 ;
  LAYER VI3 ;
  RECT 1150.900 6.340 1151.100 6.540 ;
  LAYER VI3 ;
  RECT 1150.900 5.940 1151.100 6.140 ;
  LAYER VI3 ;
  RECT 1150.500 6.340 1150.700 6.540 ;
  LAYER VI3 ;
  RECT 1150.500 5.940 1150.700 6.140 ;
  LAYER VI3 ;
  RECT 1150.100 6.340 1150.300 6.540 ;
  LAYER VI3 ;
  RECT 1150.100 5.940 1150.300 6.140 ;
  LAYER VI3 ;
  RECT 1149.700 6.340 1149.900 6.540 ;
  LAYER VI3 ;
  RECT 1149.700 5.940 1149.900 6.140 ;
  LAYER VI3 ;
  RECT 1149.300 6.340 1149.500 6.540 ;
  LAYER VI3 ;
  RECT 1149.300 5.940 1149.500 6.140 ;
  LAYER VI3 ;
  RECT 1148.900 6.340 1149.100 6.540 ;
  LAYER VI3 ;
  RECT 1148.900 5.940 1149.100 6.140 ;
  LAYER VI3 ;
  RECT 1148.500 6.340 1148.700 6.540 ;
  LAYER VI3 ;
  RECT 1148.500 5.940 1148.700 6.140 ;
  LAYER VI3 ;
  RECT 1169.580 5.880 1177.580 6.740 ;
  LAYER VI3 ;
  RECT 1177.180 6.340 1177.380 6.540 ;
  LAYER VI3 ;
  RECT 1177.180 5.940 1177.380 6.140 ;
  LAYER VI3 ;
  RECT 1176.780 6.340 1176.980 6.540 ;
  LAYER VI3 ;
  RECT 1176.780 5.940 1176.980 6.140 ;
  LAYER VI3 ;
  RECT 1176.380 6.340 1176.580 6.540 ;
  LAYER VI3 ;
  RECT 1176.380 5.940 1176.580 6.140 ;
  LAYER VI3 ;
  RECT 1175.980 6.340 1176.180 6.540 ;
  LAYER VI3 ;
  RECT 1175.980 5.940 1176.180 6.140 ;
  LAYER VI3 ;
  RECT 1175.580 6.340 1175.780 6.540 ;
  LAYER VI3 ;
  RECT 1175.580 5.940 1175.780 6.140 ;
  LAYER VI3 ;
  RECT 1175.180 6.340 1175.380 6.540 ;
  LAYER VI3 ;
  RECT 1175.180 5.940 1175.380 6.140 ;
  LAYER VI3 ;
  RECT 1174.780 6.340 1174.980 6.540 ;
  LAYER VI3 ;
  RECT 1174.780 5.940 1174.980 6.140 ;
  LAYER VI3 ;
  RECT 1174.380 6.340 1174.580 6.540 ;
  LAYER VI3 ;
  RECT 1174.380 5.940 1174.580 6.140 ;
  LAYER VI3 ;
  RECT 1173.980 6.340 1174.180 6.540 ;
  LAYER VI3 ;
  RECT 1173.980 5.940 1174.180 6.140 ;
  LAYER VI3 ;
  RECT 1173.580 6.340 1173.780 6.540 ;
  LAYER VI3 ;
  RECT 1173.580 5.940 1173.780 6.140 ;
  LAYER VI3 ;
  RECT 1173.180 6.340 1173.380 6.540 ;
  LAYER VI3 ;
  RECT 1173.180 5.940 1173.380 6.140 ;
  LAYER VI3 ;
  RECT 1172.780 6.340 1172.980 6.540 ;
  LAYER VI3 ;
  RECT 1172.780 5.940 1172.980 6.140 ;
  LAYER VI3 ;
  RECT 1172.380 6.340 1172.580 6.540 ;
  LAYER VI3 ;
  RECT 1172.380 5.940 1172.580 6.140 ;
  LAYER VI3 ;
  RECT 1171.980 6.340 1172.180 6.540 ;
  LAYER VI3 ;
  RECT 1171.980 5.940 1172.180 6.140 ;
  LAYER VI3 ;
  RECT 1171.580 6.340 1171.780 6.540 ;
  LAYER VI3 ;
  RECT 1171.580 5.940 1171.780 6.140 ;
  LAYER VI3 ;
  RECT 1171.180 6.340 1171.380 6.540 ;
  LAYER VI3 ;
  RECT 1171.180 5.940 1171.380 6.140 ;
  LAYER VI3 ;
  RECT 1170.780 6.340 1170.980 6.540 ;
  LAYER VI3 ;
  RECT 1170.780 5.940 1170.980 6.140 ;
  LAYER VI3 ;
  RECT 1170.380 6.340 1170.580 6.540 ;
  LAYER VI3 ;
  RECT 1170.380 5.940 1170.580 6.140 ;
  LAYER VI3 ;
  RECT 1169.980 6.340 1170.180 6.540 ;
  LAYER VI3 ;
  RECT 1169.980 5.940 1170.180 6.140 ;
  LAYER VI3 ;
  RECT 1169.580 6.340 1169.780 6.540 ;
  LAYER VI3 ;
  RECT 1169.580 5.940 1169.780 6.140 ;
  LAYER VI3 ;
  RECT 1189.420 5.880 1197.420 6.740 ;
  LAYER VI3 ;
  RECT 1197.020 6.340 1197.220 6.540 ;
  LAYER VI3 ;
  RECT 1197.020 5.940 1197.220 6.140 ;
  LAYER VI3 ;
  RECT 1196.620 6.340 1196.820 6.540 ;
  LAYER VI3 ;
  RECT 1196.620 5.940 1196.820 6.140 ;
  LAYER VI3 ;
  RECT 1196.220 6.340 1196.420 6.540 ;
  LAYER VI3 ;
  RECT 1196.220 5.940 1196.420 6.140 ;
  LAYER VI3 ;
  RECT 1195.820 6.340 1196.020 6.540 ;
  LAYER VI3 ;
  RECT 1195.820 5.940 1196.020 6.140 ;
  LAYER VI3 ;
  RECT 1195.420 6.340 1195.620 6.540 ;
  LAYER VI3 ;
  RECT 1195.420 5.940 1195.620 6.140 ;
  LAYER VI3 ;
  RECT 1195.020 6.340 1195.220 6.540 ;
  LAYER VI3 ;
  RECT 1195.020 5.940 1195.220 6.140 ;
  LAYER VI3 ;
  RECT 1194.620 6.340 1194.820 6.540 ;
  LAYER VI3 ;
  RECT 1194.620 5.940 1194.820 6.140 ;
  LAYER VI3 ;
  RECT 1194.220 6.340 1194.420 6.540 ;
  LAYER VI3 ;
  RECT 1194.220 5.940 1194.420 6.140 ;
  LAYER VI3 ;
  RECT 1193.820 6.340 1194.020 6.540 ;
  LAYER VI3 ;
  RECT 1193.820 5.940 1194.020 6.140 ;
  LAYER VI3 ;
  RECT 1193.420 6.340 1193.620 6.540 ;
  LAYER VI3 ;
  RECT 1193.420 5.940 1193.620 6.140 ;
  LAYER VI3 ;
  RECT 1193.020 6.340 1193.220 6.540 ;
  LAYER VI3 ;
  RECT 1193.020 5.940 1193.220 6.140 ;
  LAYER VI3 ;
  RECT 1192.620 6.340 1192.820 6.540 ;
  LAYER VI3 ;
  RECT 1192.620 5.940 1192.820 6.140 ;
  LAYER VI3 ;
  RECT 1192.220 6.340 1192.420 6.540 ;
  LAYER VI3 ;
  RECT 1192.220 5.940 1192.420 6.140 ;
  LAYER VI3 ;
  RECT 1191.820 6.340 1192.020 6.540 ;
  LAYER VI3 ;
  RECT 1191.820 5.940 1192.020 6.140 ;
  LAYER VI3 ;
  RECT 1191.420 6.340 1191.620 6.540 ;
  LAYER VI3 ;
  RECT 1191.420 5.940 1191.620 6.140 ;
  LAYER VI3 ;
  RECT 1191.020 6.340 1191.220 6.540 ;
  LAYER VI3 ;
  RECT 1191.020 5.940 1191.220 6.140 ;
  LAYER VI3 ;
  RECT 1190.620 6.340 1190.820 6.540 ;
  LAYER VI3 ;
  RECT 1190.620 5.940 1190.820 6.140 ;
  LAYER VI3 ;
  RECT 1190.220 6.340 1190.420 6.540 ;
  LAYER VI3 ;
  RECT 1190.220 5.940 1190.420 6.140 ;
  LAYER VI3 ;
  RECT 1189.820 6.340 1190.020 6.540 ;
  LAYER VI3 ;
  RECT 1189.820 5.940 1190.020 6.140 ;
  LAYER VI3 ;
  RECT 1189.420 6.340 1189.620 6.540 ;
  LAYER VI3 ;
  RECT 1189.420 5.940 1189.620 6.140 ;
  LAYER VI3 ;
  RECT 1210.500 5.880 1218.500 6.740 ;
  LAYER VI3 ;
  RECT 1218.100 6.340 1218.300 6.540 ;
  LAYER VI3 ;
  RECT 1218.100 5.940 1218.300 6.140 ;
  LAYER VI3 ;
  RECT 1217.700 6.340 1217.900 6.540 ;
  LAYER VI3 ;
  RECT 1217.700 5.940 1217.900 6.140 ;
  LAYER VI3 ;
  RECT 1217.300 6.340 1217.500 6.540 ;
  LAYER VI3 ;
  RECT 1217.300 5.940 1217.500 6.140 ;
  LAYER VI3 ;
  RECT 1216.900 6.340 1217.100 6.540 ;
  LAYER VI3 ;
  RECT 1216.900 5.940 1217.100 6.140 ;
  LAYER VI3 ;
  RECT 1216.500 6.340 1216.700 6.540 ;
  LAYER VI3 ;
  RECT 1216.500 5.940 1216.700 6.140 ;
  LAYER VI3 ;
  RECT 1216.100 6.340 1216.300 6.540 ;
  LAYER VI3 ;
  RECT 1216.100 5.940 1216.300 6.140 ;
  LAYER VI3 ;
  RECT 1215.700 6.340 1215.900 6.540 ;
  LAYER VI3 ;
  RECT 1215.700 5.940 1215.900 6.140 ;
  LAYER VI3 ;
  RECT 1215.300 6.340 1215.500 6.540 ;
  LAYER VI3 ;
  RECT 1215.300 5.940 1215.500 6.140 ;
  LAYER VI3 ;
  RECT 1214.900 6.340 1215.100 6.540 ;
  LAYER VI3 ;
  RECT 1214.900 5.940 1215.100 6.140 ;
  LAYER VI3 ;
  RECT 1214.500 6.340 1214.700 6.540 ;
  LAYER VI3 ;
  RECT 1214.500 5.940 1214.700 6.140 ;
  LAYER VI3 ;
  RECT 1214.100 6.340 1214.300 6.540 ;
  LAYER VI3 ;
  RECT 1214.100 5.940 1214.300 6.140 ;
  LAYER VI3 ;
  RECT 1213.700 6.340 1213.900 6.540 ;
  LAYER VI3 ;
  RECT 1213.700 5.940 1213.900 6.140 ;
  LAYER VI3 ;
  RECT 1213.300 6.340 1213.500 6.540 ;
  LAYER VI3 ;
  RECT 1213.300 5.940 1213.500 6.140 ;
  LAYER VI3 ;
  RECT 1212.900 6.340 1213.100 6.540 ;
  LAYER VI3 ;
  RECT 1212.900 5.940 1213.100 6.140 ;
  LAYER VI3 ;
  RECT 1212.500 6.340 1212.700 6.540 ;
  LAYER VI3 ;
  RECT 1212.500 5.940 1212.700 6.140 ;
  LAYER VI3 ;
  RECT 1212.100 6.340 1212.300 6.540 ;
  LAYER VI3 ;
  RECT 1212.100 5.940 1212.300 6.140 ;
  LAYER VI3 ;
  RECT 1211.700 6.340 1211.900 6.540 ;
  LAYER VI3 ;
  RECT 1211.700 5.940 1211.900 6.140 ;
  LAYER VI3 ;
  RECT 1211.300 6.340 1211.500 6.540 ;
  LAYER VI3 ;
  RECT 1211.300 5.940 1211.500 6.140 ;
  LAYER VI3 ;
  RECT 1210.900 6.340 1211.100 6.540 ;
  LAYER VI3 ;
  RECT 1210.900 5.940 1211.100 6.140 ;
  LAYER VI3 ;
  RECT 1210.500 6.340 1210.700 6.540 ;
  LAYER VI3 ;
  RECT 1210.500 5.940 1210.700 6.140 ;
  LAYER VI3 ;
  RECT 1230.340 5.880 1238.340 6.740 ;
  LAYER VI3 ;
  RECT 1237.940 6.340 1238.140 6.540 ;
  LAYER VI3 ;
  RECT 1237.940 5.940 1238.140 6.140 ;
  LAYER VI3 ;
  RECT 1237.540 6.340 1237.740 6.540 ;
  LAYER VI3 ;
  RECT 1237.540 5.940 1237.740 6.140 ;
  LAYER VI3 ;
  RECT 1237.140 6.340 1237.340 6.540 ;
  LAYER VI3 ;
  RECT 1237.140 5.940 1237.340 6.140 ;
  LAYER VI3 ;
  RECT 1236.740 6.340 1236.940 6.540 ;
  LAYER VI3 ;
  RECT 1236.740 5.940 1236.940 6.140 ;
  LAYER VI3 ;
  RECT 1236.340 6.340 1236.540 6.540 ;
  LAYER VI3 ;
  RECT 1236.340 5.940 1236.540 6.140 ;
  LAYER VI3 ;
  RECT 1235.940 6.340 1236.140 6.540 ;
  LAYER VI3 ;
  RECT 1235.940 5.940 1236.140 6.140 ;
  LAYER VI3 ;
  RECT 1235.540 6.340 1235.740 6.540 ;
  LAYER VI3 ;
  RECT 1235.540 5.940 1235.740 6.140 ;
  LAYER VI3 ;
  RECT 1235.140 6.340 1235.340 6.540 ;
  LAYER VI3 ;
  RECT 1235.140 5.940 1235.340 6.140 ;
  LAYER VI3 ;
  RECT 1234.740 6.340 1234.940 6.540 ;
  LAYER VI3 ;
  RECT 1234.740 5.940 1234.940 6.140 ;
  LAYER VI3 ;
  RECT 1234.340 6.340 1234.540 6.540 ;
  LAYER VI3 ;
  RECT 1234.340 5.940 1234.540 6.140 ;
  LAYER VI3 ;
  RECT 1233.940 6.340 1234.140 6.540 ;
  LAYER VI3 ;
  RECT 1233.940 5.940 1234.140 6.140 ;
  LAYER VI3 ;
  RECT 1233.540 6.340 1233.740 6.540 ;
  LAYER VI3 ;
  RECT 1233.540 5.940 1233.740 6.140 ;
  LAYER VI3 ;
  RECT 1233.140 6.340 1233.340 6.540 ;
  LAYER VI3 ;
  RECT 1233.140 5.940 1233.340 6.140 ;
  LAYER VI3 ;
  RECT 1232.740 6.340 1232.940 6.540 ;
  LAYER VI3 ;
  RECT 1232.740 5.940 1232.940 6.140 ;
  LAYER VI3 ;
  RECT 1232.340 6.340 1232.540 6.540 ;
  LAYER VI3 ;
  RECT 1232.340 5.940 1232.540 6.140 ;
  LAYER VI3 ;
  RECT 1231.940 6.340 1232.140 6.540 ;
  LAYER VI3 ;
  RECT 1231.940 5.940 1232.140 6.140 ;
  LAYER VI3 ;
  RECT 1231.540 6.340 1231.740 6.540 ;
  LAYER VI3 ;
  RECT 1231.540 5.940 1231.740 6.140 ;
  LAYER VI3 ;
  RECT 1231.140 6.340 1231.340 6.540 ;
  LAYER VI3 ;
  RECT 1231.140 5.940 1231.340 6.140 ;
  LAYER VI3 ;
  RECT 1230.740 6.340 1230.940 6.540 ;
  LAYER VI3 ;
  RECT 1230.740 5.940 1230.940 6.140 ;
  LAYER VI3 ;
  RECT 1230.340 6.340 1230.540 6.540 ;
  LAYER VI3 ;
  RECT 1230.340 5.940 1230.540 6.140 ;
  LAYER VI3 ;
  RECT 1251.420 5.880 1259.420 6.740 ;
  LAYER VI3 ;
  RECT 1259.020 6.340 1259.220 6.540 ;
  LAYER VI3 ;
  RECT 1259.020 5.940 1259.220 6.140 ;
  LAYER VI3 ;
  RECT 1258.620 6.340 1258.820 6.540 ;
  LAYER VI3 ;
  RECT 1258.620 5.940 1258.820 6.140 ;
  LAYER VI3 ;
  RECT 1258.220 6.340 1258.420 6.540 ;
  LAYER VI3 ;
  RECT 1258.220 5.940 1258.420 6.140 ;
  LAYER VI3 ;
  RECT 1257.820 6.340 1258.020 6.540 ;
  LAYER VI3 ;
  RECT 1257.820 5.940 1258.020 6.140 ;
  LAYER VI3 ;
  RECT 1257.420 6.340 1257.620 6.540 ;
  LAYER VI3 ;
  RECT 1257.420 5.940 1257.620 6.140 ;
  LAYER VI3 ;
  RECT 1257.020 6.340 1257.220 6.540 ;
  LAYER VI3 ;
  RECT 1257.020 5.940 1257.220 6.140 ;
  LAYER VI3 ;
  RECT 1256.620 6.340 1256.820 6.540 ;
  LAYER VI3 ;
  RECT 1256.620 5.940 1256.820 6.140 ;
  LAYER VI3 ;
  RECT 1256.220 6.340 1256.420 6.540 ;
  LAYER VI3 ;
  RECT 1256.220 5.940 1256.420 6.140 ;
  LAYER VI3 ;
  RECT 1255.820 6.340 1256.020 6.540 ;
  LAYER VI3 ;
  RECT 1255.820 5.940 1256.020 6.140 ;
  LAYER VI3 ;
  RECT 1255.420 6.340 1255.620 6.540 ;
  LAYER VI3 ;
  RECT 1255.420 5.940 1255.620 6.140 ;
  LAYER VI3 ;
  RECT 1255.020 6.340 1255.220 6.540 ;
  LAYER VI3 ;
  RECT 1255.020 5.940 1255.220 6.140 ;
  LAYER VI3 ;
  RECT 1254.620 6.340 1254.820 6.540 ;
  LAYER VI3 ;
  RECT 1254.620 5.940 1254.820 6.140 ;
  LAYER VI3 ;
  RECT 1254.220 6.340 1254.420 6.540 ;
  LAYER VI3 ;
  RECT 1254.220 5.940 1254.420 6.140 ;
  LAYER VI3 ;
  RECT 1253.820 6.340 1254.020 6.540 ;
  LAYER VI3 ;
  RECT 1253.820 5.940 1254.020 6.140 ;
  LAYER VI3 ;
  RECT 1253.420 6.340 1253.620 6.540 ;
  LAYER VI3 ;
  RECT 1253.420 5.940 1253.620 6.140 ;
  LAYER VI3 ;
  RECT 1253.020 6.340 1253.220 6.540 ;
  LAYER VI3 ;
  RECT 1253.020 5.940 1253.220 6.140 ;
  LAYER VI3 ;
  RECT 1252.620 6.340 1252.820 6.540 ;
  LAYER VI3 ;
  RECT 1252.620 5.940 1252.820 6.140 ;
  LAYER VI3 ;
  RECT 1252.220 6.340 1252.420 6.540 ;
  LAYER VI3 ;
  RECT 1252.220 5.940 1252.420 6.140 ;
  LAYER VI3 ;
  RECT 1251.820 6.340 1252.020 6.540 ;
  LAYER VI3 ;
  RECT 1251.820 5.940 1252.020 6.140 ;
  LAYER VI3 ;
  RECT 1251.420 6.340 1251.620 6.540 ;
  LAYER VI3 ;
  RECT 1251.420 5.940 1251.620 6.140 ;
  LAYER VI3 ;
  RECT 1271.260 5.880 1279.260 6.740 ;
  LAYER VI3 ;
  RECT 1278.860 6.340 1279.060 6.540 ;
  LAYER VI3 ;
  RECT 1278.860 5.940 1279.060 6.140 ;
  LAYER VI3 ;
  RECT 1278.460 6.340 1278.660 6.540 ;
  LAYER VI3 ;
  RECT 1278.460 5.940 1278.660 6.140 ;
  LAYER VI3 ;
  RECT 1278.060 6.340 1278.260 6.540 ;
  LAYER VI3 ;
  RECT 1278.060 5.940 1278.260 6.140 ;
  LAYER VI3 ;
  RECT 1277.660 6.340 1277.860 6.540 ;
  LAYER VI3 ;
  RECT 1277.660 5.940 1277.860 6.140 ;
  LAYER VI3 ;
  RECT 1277.260 6.340 1277.460 6.540 ;
  LAYER VI3 ;
  RECT 1277.260 5.940 1277.460 6.140 ;
  LAYER VI3 ;
  RECT 1276.860 6.340 1277.060 6.540 ;
  LAYER VI3 ;
  RECT 1276.860 5.940 1277.060 6.140 ;
  LAYER VI3 ;
  RECT 1276.460 6.340 1276.660 6.540 ;
  LAYER VI3 ;
  RECT 1276.460 5.940 1276.660 6.140 ;
  LAYER VI3 ;
  RECT 1276.060 6.340 1276.260 6.540 ;
  LAYER VI3 ;
  RECT 1276.060 5.940 1276.260 6.140 ;
  LAYER VI3 ;
  RECT 1275.660 6.340 1275.860 6.540 ;
  LAYER VI3 ;
  RECT 1275.660 5.940 1275.860 6.140 ;
  LAYER VI3 ;
  RECT 1275.260 6.340 1275.460 6.540 ;
  LAYER VI3 ;
  RECT 1275.260 5.940 1275.460 6.140 ;
  LAYER VI3 ;
  RECT 1274.860 6.340 1275.060 6.540 ;
  LAYER VI3 ;
  RECT 1274.860 5.940 1275.060 6.140 ;
  LAYER VI3 ;
  RECT 1274.460 6.340 1274.660 6.540 ;
  LAYER VI3 ;
  RECT 1274.460 5.940 1274.660 6.140 ;
  LAYER VI3 ;
  RECT 1274.060 6.340 1274.260 6.540 ;
  LAYER VI3 ;
  RECT 1274.060 5.940 1274.260 6.140 ;
  LAYER VI3 ;
  RECT 1273.660 6.340 1273.860 6.540 ;
  LAYER VI3 ;
  RECT 1273.660 5.940 1273.860 6.140 ;
  LAYER VI3 ;
  RECT 1273.260 6.340 1273.460 6.540 ;
  LAYER VI3 ;
  RECT 1273.260 5.940 1273.460 6.140 ;
  LAYER VI3 ;
  RECT 1272.860 6.340 1273.060 6.540 ;
  LAYER VI3 ;
  RECT 1272.860 5.940 1273.060 6.140 ;
  LAYER VI3 ;
  RECT 1272.460 6.340 1272.660 6.540 ;
  LAYER VI3 ;
  RECT 1272.460 5.940 1272.660 6.140 ;
  LAYER VI3 ;
  RECT 1272.060 6.340 1272.260 6.540 ;
  LAYER VI3 ;
  RECT 1272.060 5.940 1272.260 6.140 ;
  LAYER VI3 ;
  RECT 1271.660 6.340 1271.860 6.540 ;
  LAYER VI3 ;
  RECT 1271.660 5.940 1271.860 6.140 ;
  LAYER VI3 ;
  RECT 1271.260 6.340 1271.460 6.540 ;
  LAYER VI3 ;
  RECT 1271.260 5.940 1271.460 6.140 ;
  LAYER VI3 ;
  RECT 1292.340 5.880 1300.340 6.740 ;
  LAYER VI3 ;
  RECT 1299.940 6.340 1300.140 6.540 ;
  LAYER VI3 ;
  RECT 1299.940 5.940 1300.140 6.140 ;
  LAYER VI3 ;
  RECT 1299.540 6.340 1299.740 6.540 ;
  LAYER VI3 ;
  RECT 1299.540 5.940 1299.740 6.140 ;
  LAYER VI3 ;
  RECT 1299.140 6.340 1299.340 6.540 ;
  LAYER VI3 ;
  RECT 1299.140 5.940 1299.340 6.140 ;
  LAYER VI3 ;
  RECT 1298.740 6.340 1298.940 6.540 ;
  LAYER VI3 ;
  RECT 1298.740 5.940 1298.940 6.140 ;
  LAYER VI3 ;
  RECT 1298.340 6.340 1298.540 6.540 ;
  LAYER VI3 ;
  RECT 1298.340 5.940 1298.540 6.140 ;
  LAYER VI3 ;
  RECT 1297.940 6.340 1298.140 6.540 ;
  LAYER VI3 ;
  RECT 1297.940 5.940 1298.140 6.140 ;
  LAYER VI3 ;
  RECT 1297.540 6.340 1297.740 6.540 ;
  LAYER VI3 ;
  RECT 1297.540 5.940 1297.740 6.140 ;
  LAYER VI3 ;
  RECT 1297.140 6.340 1297.340 6.540 ;
  LAYER VI3 ;
  RECT 1297.140 5.940 1297.340 6.140 ;
  LAYER VI3 ;
  RECT 1296.740 6.340 1296.940 6.540 ;
  LAYER VI3 ;
  RECT 1296.740 5.940 1296.940 6.140 ;
  LAYER VI3 ;
  RECT 1296.340 6.340 1296.540 6.540 ;
  LAYER VI3 ;
  RECT 1296.340 5.940 1296.540 6.140 ;
  LAYER VI3 ;
  RECT 1295.940 6.340 1296.140 6.540 ;
  LAYER VI3 ;
  RECT 1295.940 5.940 1296.140 6.140 ;
  LAYER VI3 ;
  RECT 1295.540 6.340 1295.740 6.540 ;
  LAYER VI3 ;
  RECT 1295.540 5.940 1295.740 6.140 ;
  LAYER VI3 ;
  RECT 1295.140 6.340 1295.340 6.540 ;
  LAYER VI3 ;
  RECT 1295.140 5.940 1295.340 6.140 ;
  LAYER VI3 ;
  RECT 1294.740 6.340 1294.940 6.540 ;
  LAYER VI3 ;
  RECT 1294.740 5.940 1294.940 6.140 ;
  LAYER VI3 ;
  RECT 1294.340 6.340 1294.540 6.540 ;
  LAYER VI3 ;
  RECT 1294.340 5.940 1294.540 6.140 ;
  LAYER VI3 ;
  RECT 1293.940 6.340 1294.140 6.540 ;
  LAYER VI3 ;
  RECT 1293.940 5.940 1294.140 6.140 ;
  LAYER VI3 ;
  RECT 1293.540 6.340 1293.740 6.540 ;
  LAYER VI3 ;
  RECT 1293.540 5.940 1293.740 6.140 ;
  LAYER VI3 ;
  RECT 1293.140 6.340 1293.340 6.540 ;
  LAYER VI3 ;
  RECT 1293.140 5.940 1293.340 6.140 ;
  LAYER VI3 ;
  RECT 1292.740 6.340 1292.940 6.540 ;
  LAYER VI3 ;
  RECT 1292.740 5.940 1292.940 6.140 ;
  LAYER VI3 ;
  RECT 1292.340 6.340 1292.540 6.540 ;
  LAYER VI3 ;
  RECT 1292.340 5.940 1292.540 6.140 ;
  LAYER VI3 ;
  RECT 1312.180 5.880 1320.180 6.740 ;
  LAYER VI3 ;
  RECT 1319.780 6.340 1319.980 6.540 ;
  LAYER VI3 ;
  RECT 1319.780 5.940 1319.980 6.140 ;
  LAYER VI3 ;
  RECT 1319.380 6.340 1319.580 6.540 ;
  LAYER VI3 ;
  RECT 1319.380 5.940 1319.580 6.140 ;
  LAYER VI3 ;
  RECT 1318.980 6.340 1319.180 6.540 ;
  LAYER VI3 ;
  RECT 1318.980 5.940 1319.180 6.140 ;
  LAYER VI3 ;
  RECT 1318.580 6.340 1318.780 6.540 ;
  LAYER VI3 ;
  RECT 1318.580 5.940 1318.780 6.140 ;
  LAYER VI3 ;
  RECT 1318.180 6.340 1318.380 6.540 ;
  LAYER VI3 ;
  RECT 1318.180 5.940 1318.380 6.140 ;
  LAYER VI3 ;
  RECT 1317.780 6.340 1317.980 6.540 ;
  LAYER VI3 ;
  RECT 1317.780 5.940 1317.980 6.140 ;
  LAYER VI3 ;
  RECT 1317.380 6.340 1317.580 6.540 ;
  LAYER VI3 ;
  RECT 1317.380 5.940 1317.580 6.140 ;
  LAYER VI3 ;
  RECT 1316.980 6.340 1317.180 6.540 ;
  LAYER VI3 ;
  RECT 1316.980 5.940 1317.180 6.140 ;
  LAYER VI3 ;
  RECT 1316.580 6.340 1316.780 6.540 ;
  LAYER VI3 ;
  RECT 1316.580 5.940 1316.780 6.140 ;
  LAYER VI3 ;
  RECT 1316.180 6.340 1316.380 6.540 ;
  LAYER VI3 ;
  RECT 1316.180 5.940 1316.380 6.140 ;
  LAYER VI3 ;
  RECT 1315.780 6.340 1315.980 6.540 ;
  LAYER VI3 ;
  RECT 1315.780 5.940 1315.980 6.140 ;
  LAYER VI3 ;
  RECT 1315.380 6.340 1315.580 6.540 ;
  LAYER VI3 ;
  RECT 1315.380 5.940 1315.580 6.140 ;
  LAYER VI3 ;
  RECT 1314.980 6.340 1315.180 6.540 ;
  LAYER VI3 ;
  RECT 1314.980 5.940 1315.180 6.140 ;
  LAYER VI3 ;
  RECT 1314.580 6.340 1314.780 6.540 ;
  LAYER VI3 ;
  RECT 1314.580 5.940 1314.780 6.140 ;
  LAYER VI3 ;
  RECT 1314.180 6.340 1314.380 6.540 ;
  LAYER VI3 ;
  RECT 1314.180 5.940 1314.380 6.140 ;
  LAYER VI3 ;
  RECT 1313.780 6.340 1313.980 6.540 ;
  LAYER VI3 ;
  RECT 1313.780 5.940 1313.980 6.140 ;
  LAYER VI3 ;
  RECT 1313.380 6.340 1313.580 6.540 ;
  LAYER VI3 ;
  RECT 1313.380 5.940 1313.580 6.140 ;
  LAYER VI3 ;
  RECT 1312.980 6.340 1313.180 6.540 ;
  LAYER VI3 ;
  RECT 1312.980 5.940 1313.180 6.140 ;
  LAYER VI3 ;
  RECT 1312.580 6.340 1312.780 6.540 ;
  LAYER VI3 ;
  RECT 1312.580 5.940 1312.780 6.140 ;
  LAYER VI3 ;
  RECT 1312.180 6.340 1312.380 6.540 ;
  LAYER VI3 ;
  RECT 1312.180 5.940 1312.380 6.140 ;
  LAYER VI3 ;
  RECT 1333.260 5.880 1341.260 6.740 ;
  LAYER VI3 ;
  RECT 1340.860 6.340 1341.060 6.540 ;
  LAYER VI3 ;
  RECT 1340.860 5.940 1341.060 6.140 ;
  LAYER VI3 ;
  RECT 1340.460 6.340 1340.660 6.540 ;
  LAYER VI3 ;
  RECT 1340.460 5.940 1340.660 6.140 ;
  LAYER VI3 ;
  RECT 1340.060 6.340 1340.260 6.540 ;
  LAYER VI3 ;
  RECT 1340.060 5.940 1340.260 6.140 ;
  LAYER VI3 ;
  RECT 1339.660 6.340 1339.860 6.540 ;
  LAYER VI3 ;
  RECT 1339.660 5.940 1339.860 6.140 ;
  LAYER VI3 ;
  RECT 1339.260 6.340 1339.460 6.540 ;
  LAYER VI3 ;
  RECT 1339.260 5.940 1339.460 6.140 ;
  LAYER VI3 ;
  RECT 1338.860 6.340 1339.060 6.540 ;
  LAYER VI3 ;
  RECT 1338.860 5.940 1339.060 6.140 ;
  LAYER VI3 ;
  RECT 1338.460 6.340 1338.660 6.540 ;
  LAYER VI3 ;
  RECT 1338.460 5.940 1338.660 6.140 ;
  LAYER VI3 ;
  RECT 1338.060 6.340 1338.260 6.540 ;
  LAYER VI3 ;
  RECT 1338.060 5.940 1338.260 6.140 ;
  LAYER VI3 ;
  RECT 1337.660 6.340 1337.860 6.540 ;
  LAYER VI3 ;
  RECT 1337.660 5.940 1337.860 6.140 ;
  LAYER VI3 ;
  RECT 1337.260 6.340 1337.460 6.540 ;
  LAYER VI3 ;
  RECT 1337.260 5.940 1337.460 6.140 ;
  LAYER VI3 ;
  RECT 1336.860 6.340 1337.060 6.540 ;
  LAYER VI3 ;
  RECT 1336.860 5.940 1337.060 6.140 ;
  LAYER VI3 ;
  RECT 1336.460 6.340 1336.660 6.540 ;
  LAYER VI3 ;
  RECT 1336.460 5.940 1336.660 6.140 ;
  LAYER VI3 ;
  RECT 1336.060 6.340 1336.260 6.540 ;
  LAYER VI3 ;
  RECT 1336.060 5.940 1336.260 6.140 ;
  LAYER VI3 ;
  RECT 1335.660 6.340 1335.860 6.540 ;
  LAYER VI3 ;
  RECT 1335.660 5.940 1335.860 6.140 ;
  LAYER VI3 ;
  RECT 1335.260 6.340 1335.460 6.540 ;
  LAYER VI3 ;
  RECT 1335.260 5.940 1335.460 6.140 ;
  LAYER VI3 ;
  RECT 1334.860 6.340 1335.060 6.540 ;
  LAYER VI3 ;
  RECT 1334.860 5.940 1335.060 6.140 ;
  LAYER VI3 ;
  RECT 1334.460 6.340 1334.660 6.540 ;
  LAYER VI3 ;
  RECT 1334.460 5.940 1334.660 6.140 ;
  LAYER VI3 ;
  RECT 1334.060 6.340 1334.260 6.540 ;
  LAYER VI3 ;
  RECT 1334.060 5.940 1334.260 6.140 ;
  LAYER VI3 ;
  RECT 1333.660 6.340 1333.860 6.540 ;
  LAYER VI3 ;
  RECT 1333.660 5.940 1333.860 6.140 ;
  LAYER VI3 ;
  RECT 1333.260 6.340 1333.460 6.540 ;
  LAYER VI3 ;
  RECT 1333.260 5.940 1333.460 6.140 ;
  LAYER VI3 ;
  RECT 1353.100 5.880 1361.100 6.740 ;
  LAYER VI3 ;
  RECT 1360.700 6.340 1360.900 6.540 ;
  LAYER VI3 ;
  RECT 1360.700 5.940 1360.900 6.140 ;
  LAYER VI3 ;
  RECT 1360.300 6.340 1360.500 6.540 ;
  LAYER VI3 ;
  RECT 1360.300 5.940 1360.500 6.140 ;
  LAYER VI3 ;
  RECT 1359.900 6.340 1360.100 6.540 ;
  LAYER VI3 ;
  RECT 1359.900 5.940 1360.100 6.140 ;
  LAYER VI3 ;
  RECT 1359.500 6.340 1359.700 6.540 ;
  LAYER VI3 ;
  RECT 1359.500 5.940 1359.700 6.140 ;
  LAYER VI3 ;
  RECT 1359.100 6.340 1359.300 6.540 ;
  LAYER VI3 ;
  RECT 1359.100 5.940 1359.300 6.140 ;
  LAYER VI3 ;
  RECT 1358.700 6.340 1358.900 6.540 ;
  LAYER VI3 ;
  RECT 1358.700 5.940 1358.900 6.140 ;
  LAYER VI3 ;
  RECT 1358.300 6.340 1358.500 6.540 ;
  LAYER VI3 ;
  RECT 1358.300 5.940 1358.500 6.140 ;
  LAYER VI3 ;
  RECT 1357.900 6.340 1358.100 6.540 ;
  LAYER VI3 ;
  RECT 1357.900 5.940 1358.100 6.140 ;
  LAYER VI3 ;
  RECT 1357.500 6.340 1357.700 6.540 ;
  LAYER VI3 ;
  RECT 1357.500 5.940 1357.700 6.140 ;
  LAYER VI3 ;
  RECT 1357.100 6.340 1357.300 6.540 ;
  LAYER VI3 ;
  RECT 1357.100 5.940 1357.300 6.140 ;
  LAYER VI3 ;
  RECT 1356.700 6.340 1356.900 6.540 ;
  LAYER VI3 ;
  RECT 1356.700 5.940 1356.900 6.140 ;
  LAYER VI3 ;
  RECT 1356.300 6.340 1356.500 6.540 ;
  LAYER VI3 ;
  RECT 1356.300 5.940 1356.500 6.140 ;
  LAYER VI3 ;
  RECT 1355.900 6.340 1356.100 6.540 ;
  LAYER VI3 ;
  RECT 1355.900 5.940 1356.100 6.140 ;
  LAYER VI3 ;
  RECT 1355.500 6.340 1355.700 6.540 ;
  LAYER VI3 ;
  RECT 1355.500 5.940 1355.700 6.140 ;
  LAYER VI3 ;
  RECT 1355.100 6.340 1355.300 6.540 ;
  LAYER VI3 ;
  RECT 1355.100 5.940 1355.300 6.140 ;
  LAYER VI3 ;
  RECT 1354.700 6.340 1354.900 6.540 ;
  LAYER VI3 ;
  RECT 1354.700 5.940 1354.900 6.140 ;
  LAYER VI3 ;
  RECT 1354.300 6.340 1354.500 6.540 ;
  LAYER VI3 ;
  RECT 1354.300 5.940 1354.500 6.140 ;
  LAYER VI3 ;
  RECT 1353.900 6.340 1354.100 6.540 ;
  LAYER VI3 ;
  RECT 1353.900 5.940 1354.100 6.140 ;
  LAYER VI3 ;
  RECT 1353.500 6.340 1353.700 6.540 ;
  LAYER VI3 ;
  RECT 1353.500 5.940 1353.700 6.140 ;
  LAYER VI3 ;
  RECT 1353.100 6.340 1353.300 6.540 ;
  LAYER VI3 ;
  RECT 1353.100 5.940 1353.300 6.140 ;
  LAYER VI3 ;
  RECT 684.720 5.880 688.170 6.740 ;
  LAYER VI3 ;
  RECT 687.920 6.340 688.120 6.540 ;
  LAYER VI3 ;
  RECT 687.920 5.940 688.120 6.140 ;
  LAYER VI3 ;
  RECT 687.520 6.340 687.720 6.540 ;
  LAYER VI3 ;
  RECT 687.520 5.940 687.720 6.140 ;
  LAYER VI3 ;
  RECT 687.120 6.340 687.320 6.540 ;
  LAYER VI3 ;
  RECT 687.120 5.940 687.320 6.140 ;
  LAYER VI3 ;
  RECT 686.720 6.340 686.920 6.540 ;
  LAYER VI3 ;
  RECT 686.720 5.940 686.920 6.140 ;
  LAYER VI3 ;
  RECT 686.320 6.340 686.520 6.540 ;
  LAYER VI3 ;
  RECT 686.320 5.940 686.520 6.140 ;
  LAYER VI3 ;
  RECT 685.920 6.340 686.120 6.540 ;
  LAYER VI3 ;
  RECT 685.920 5.940 686.120 6.140 ;
  LAYER VI3 ;
  RECT 685.520 6.340 685.720 6.540 ;
  LAYER VI3 ;
  RECT 685.520 5.940 685.720 6.140 ;
  LAYER VI3 ;
  RECT 685.120 6.340 685.320 6.540 ;
  LAYER VI3 ;
  RECT 685.120 5.940 685.320 6.140 ;
  LAYER VI3 ;
  RECT 684.720 6.340 684.920 6.540 ;
  LAYER VI3 ;
  RECT 684.720 5.940 684.920 6.140 ;
  LAYER VI3 ;
  RECT 693.570 5.880 699.490 6.740 ;
  LAYER VI3 ;
  RECT 699.170 6.340 699.370 6.540 ;
  LAYER VI3 ;
  RECT 699.170 5.940 699.370 6.140 ;
  LAYER VI3 ;
  RECT 698.770 6.340 698.970 6.540 ;
  LAYER VI3 ;
  RECT 698.770 5.940 698.970 6.140 ;
  LAYER VI3 ;
  RECT 698.370 6.340 698.570 6.540 ;
  LAYER VI3 ;
  RECT 698.370 5.940 698.570 6.140 ;
  LAYER VI3 ;
  RECT 697.970 6.340 698.170 6.540 ;
  LAYER VI3 ;
  RECT 697.970 5.940 698.170 6.140 ;
  LAYER VI3 ;
  RECT 697.570 6.340 697.770 6.540 ;
  LAYER VI3 ;
  RECT 697.570 5.940 697.770 6.140 ;
  LAYER VI3 ;
  RECT 697.170 6.340 697.370 6.540 ;
  LAYER VI3 ;
  RECT 697.170 5.940 697.370 6.140 ;
  LAYER VI3 ;
  RECT 696.770 6.340 696.970 6.540 ;
  LAYER VI3 ;
  RECT 696.770 5.940 696.970 6.140 ;
  LAYER VI3 ;
  RECT 696.370 6.340 696.570 6.540 ;
  LAYER VI3 ;
  RECT 696.370 5.940 696.570 6.140 ;
  LAYER VI3 ;
  RECT 695.970 6.340 696.170 6.540 ;
  LAYER VI3 ;
  RECT 695.970 5.940 696.170 6.140 ;
  LAYER VI3 ;
  RECT 695.570 6.340 695.770 6.540 ;
  LAYER VI3 ;
  RECT 695.570 5.940 695.770 6.140 ;
  LAYER VI3 ;
  RECT 695.170 6.340 695.370 6.540 ;
  LAYER VI3 ;
  RECT 695.170 5.940 695.370 6.140 ;
  LAYER VI3 ;
  RECT 694.770 6.340 694.970 6.540 ;
  LAYER VI3 ;
  RECT 694.770 5.940 694.970 6.140 ;
  LAYER VI3 ;
  RECT 694.370 6.340 694.570 6.540 ;
  LAYER VI3 ;
  RECT 694.370 5.940 694.570 6.140 ;
  LAYER VI3 ;
  RECT 693.970 6.340 694.170 6.540 ;
  LAYER VI3 ;
  RECT 693.970 5.940 694.170 6.140 ;
  LAYER VI3 ;
  RECT 693.570 6.340 693.770 6.540 ;
  LAYER VI3 ;
  RECT 693.570 5.940 693.770 6.140 ;
  LAYER VI3 ;
  RECT 676.440 5.880 678.200 6.740 ;
  LAYER VI3 ;
  RECT 677.640 6.340 677.840 6.540 ;
  LAYER VI3 ;
  RECT 677.640 5.940 677.840 6.140 ;
  LAYER VI3 ;
  RECT 677.240 6.340 677.440 6.540 ;
  LAYER VI3 ;
  RECT 677.240 5.940 677.440 6.140 ;
  LAYER VI3 ;
  RECT 676.840 6.340 677.040 6.540 ;
  LAYER VI3 ;
  RECT 676.840 5.940 677.040 6.140 ;
  LAYER VI3 ;
  RECT 676.440 6.340 676.640 6.540 ;
  LAYER VI3 ;
  RECT 676.440 5.940 676.640 6.140 ;
  LAYER VI3 ;
  RECT 671.100 5.880 672.860 6.740 ;
  LAYER VI3 ;
  RECT 672.300 6.340 672.500 6.540 ;
  LAYER VI3 ;
  RECT 672.300 5.940 672.500 6.140 ;
  LAYER VI3 ;
  RECT 671.900 6.340 672.100 6.540 ;
  LAYER VI3 ;
  RECT 671.900 5.940 672.100 6.140 ;
  LAYER VI3 ;
  RECT 671.500 6.340 671.700 6.540 ;
  LAYER VI3 ;
  RECT 671.500 5.940 671.700 6.140 ;
  LAYER VI3 ;
  RECT 671.100 6.340 671.300 6.540 ;
  LAYER VI3 ;
  RECT 671.100 5.940 671.300 6.140 ;
  LAYER VI3 ;
  RECT 667.100 5.880 668.860 6.740 ;
  LAYER VI3 ;
  RECT 668.300 6.340 668.500 6.540 ;
  LAYER VI3 ;
  RECT 668.300 5.940 668.500 6.140 ;
  LAYER VI3 ;
  RECT 667.900 6.340 668.100 6.540 ;
  LAYER VI3 ;
  RECT 667.900 5.940 668.100 6.140 ;
  LAYER VI3 ;
  RECT 667.500 6.340 667.700 6.540 ;
  LAYER VI3 ;
  RECT 667.500 5.940 667.700 6.140 ;
  LAYER VI3 ;
  RECT 667.100 6.340 667.300 6.540 ;
  LAYER VI3 ;
  RECT 667.100 5.940 667.300 6.140 ;
  LAYER VI3 ;
  RECT 663.100 5.880 664.860 6.740 ;
  LAYER VI3 ;
  RECT 664.300 6.340 664.500 6.540 ;
  LAYER VI3 ;
  RECT 664.300 5.940 664.500 6.140 ;
  LAYER VI3 ;
  RECT 663.900 6.340 664.100 6.540 ;
  LAYER VI3 ;
  RECT 663.900 5.940 664.100 6.140 ;
  LAYER VI3 ;
  RECT 663.500 6.340 663.700 6.540 ;
  LAYER VI3 ;
  RECT 663.500 5.940 663.700 6.140 ;
  LAYER VI3 ;
  RECT 663.100 6.340 663.300 6.540 ;
  LAYER VI3 ;
  RECT 663.100 5.940 663.300 6.140 ;
  LAYER VI3 ;
  RECT 4.280 57.100 5.140 61.420 ;
  LAYER VI3 ;
  RECT 4.740 61.100 4.940 61.300 ;
  LAYER VI3 ;
  RECT 4.740 60.700 4.940 60.900 ;
  LAYER VI3 ;
  RECT 4.740 60.300 4.940 60.500 ;
  LAYER VI3 ;
  RECT 4.740 59.900 4.940 60.100 ;
  LAYER VI3 ;
  RECT 4.740 59.500 4.940 59.700 ;
  LAYER VI3 ;
  RECT 4.740 59.100 4.940 59.300 ;
  LAYER VI3 ;
  RECT 4.740 58.700 4.940 58.900 ;
  LAYER VI3 ;
  RECT 4.740 58.300 4.940 58.500 ;
  LAYER VI3 ;
  RECT 4.740 57.900 4.940 58.100 ;
  LAYER VI3 ;
  RECT 4.740 57.500 4.940 57.700 ;
  LAYER VI3 ;
  RECT 4.740 57.100 4.940 57.300 ;
  LAYER VI3 ;
  RECT 4.340 61.100 4.540 61.300 ;
  LAYER VI3 ;
  RECT 4.340 60.700 4.540 60.900 ;
  LAYER VI3 ;
  RECT 4.340 60.300 4.540 60.500 ;
  LAYER VI3 ;
  RECT 4.340 59.900 4.540 60.100 ;
  LAYER VI3 ;
  RECT 4.340 59.500 4.540 59.700 ;
  LAYER VI3 ;
  RECT 4.340 59.100 4.540 59.300 ;
  LAYER VI3 ;
  RECT 4.340 58.700 4.540 58.900 ;
  LAYER VI3 ;
  RECT 4.340 58.300 4.540 58.500 ;
  LAYER VI3 ;
  RECT 4.340 57.900 4.540 58.100 ;
  LAYER VI3 ;
  RECT 4.340 57.500 4.540 57.700 ;
  LAYER VI3 ;
  RECT 4.340 57.100 4.540 57.300 ;
  LAYER VI2 ;
  RECT 4.280 57.100 5.140 61.420 ;
  LAYER VI2 ;
  RECT 4.740 61.100 4.940 61.300 ;
  LAYER VI2 ;
  RECT 4.740 60.700 4.940 60.900 ;
  LAYER VI2 ;
  RECT 4.740 60.300 4.940 60.500 ;
  LAYER VI2 ;
  RECT 4.740 59.900 4.940 60.100 ;
  LAYER VI2 ;
  RECT 4.740 59.500 4.940 59.700 ;
  LAYER VI2 ;
  RECT 4.740 59.100 4.940 59.300 ;
  LAYER VI2 ;
  RECT 4.740 58.700 4.940 58.900 ;
  LAYER VI2 ;
  RECT 4.740 58.300 4.940 58.500 ;
  LAYER VI2 ;
  RECT 4.740 57.900 4.940 58.100 ;
  LAYER VI2 ;
  RECT 4.740 57.500 4.940 57.700 ;
  LAYER VI2 ;
  RECT 4.740 57.100 4.940 57.300 ;
  LAYER VI2 ;
  RECT 4.340 61.100 4.540 61.300 ;
  LAYER VI2 ;
  RECT 4.340 60.700 4.540 60.900 ;
  LAYER VI2 ;
  RECT 4.340 60.300 4.540 60.500 ;
  LAYER VI2 ;
  RECT 4.340 59.900 4.540 60.100 ;
  LAYER VI2 ;
  RECT 4.340 59.500 4.540 59.700 ;
  LAYER VI2 ;
  RECT 4.340 59.100 4.540 59.300 ;
  LAYER VI2 ;
  RECT 4.340 58.700 4.540 58.900 ;
  LAYER VI2 ;
  RECT 4.340 58.300 4.540 58.500 ;
  LAYER VI2 ;
  RECT 4.340 57.900 4.540 58.100 ;
  LAYER VI2 ;
  RECT 4.340 57.500 4.540 57.700 ;
  LAYER VI2 ;
  RECT 4.340 57.100 4.540 57.300 ;
  LAYER VI3 ;
  RECT 4.280 45.560 5.140 46.160 ;
  LAYER VI3 ;
  RECT 4.680 45.620 4.880 45.820 ;
  LAYER VI3 ;
  RECT 4.280 45.620 4.480 45.820 ;
  LAYER VI2 ;
  RECT 4.280 45.560 5.140 46.160 ;
  LAYER VI2 ;
  RECT 4.680 45.620 4.880 45.820 ;
  LAYER VI2 ;
  RECT 4.280 45.620 4.480 45.820 ;
  LAYER VI3 ;
  RECT 4.280 39.480 5.140 40.080 ;
  LAYER VI3 ;
  RECT 4.680 39.540 4.880 39.740 ;
  LAYER VI3 ;
  RECT 4.280 39.540 4.480 39.740 ;
  LAYER VI2 ;
  RECT 4.280 39.480 5.140 40.080 ;
  LAYER VI2 ;
  RECT 4.680 39.540 4.880 39.740 ;
  LAYER VI2 ;
  RECT 4.280 39.540 4.480 39.740 ;
  LAYER VI3 ;
  RECT 4.280 36.320 5.140 37.320 ;
  LAYER VI3 ;
  RECT 4.740 36.720 4.940 36.920 ;
  LAYER VI3 ;
  RECT 4.740 36.320 4.940 36.520 ;
  LAYER VI3 ;
  RECT 4.340 36.720 4.540 36.920 ;
  LAYER VI3 ;
  RECT 4.340 36.320 4.540 36.520 ;
  LAYER VI2 ;
  RECT 4.280 36.320 5.140 37.320 ;
  LAYER VI2 ;
  RECT 4.740 36.720 4.940 36.920 ;
  LAYER VI2 ;
  RECT 4.740 36.320 4.940 36.520 ;
  LAYER VI2 ;
  RECT 4.340 36.720 4.540 36.920 ;
  LAYER VI2 ;
  RECT 4.340 36.320 4.540 36.520 ;
  LAYER VI3 ;
  RECT 4.280 24.170 5.140 25.170 ;
  LAYER VI3 ;
  RECT 4.740 24.570 4.940 24.770 ;
  LAYER VI3 ;
  RECT 4.740 24.170 4.940 24.370 ;
  LAYER VI3 ;
  RECT 4.340 24.570 4.540 24.770 ;
  LAYER VI3 ;
  RECT 4.340 24.170 4.540 24.370 ;
  LAYER VI2 ;
  RECT 4.280 24.170 5.140 25.170 ;
  LAYER VI2 ;
  RECT 4.740 24.570 4.940 24.770 ;
  LAYER VI2 ;
  RECT 4.740 24.170 4.940 24.370 ;
  LAYER VI2 ;
  RECT 4.340 24.570 4.540 24.770 ;
  LAYER VI2 ;
  RECT 4.340 24.170 4.540 24.370 ;
  LAYER VI3 ;
  RECT 4.280 21.230 5.140 22.070 ;
  LAYER VI3 ;
  RECT 4.680 21.690 4.880 21.890 ;
  LAYER VI3 ;
  RECT 4.680 21.290 4.880 21.490 ;
  LAYER VI3 ;
  RECT 4.280 21.690 4.480 21.890 ;
  LAYER VI3 ;
  RECT 4.280 21.290 4.480 21.490 ;
  LAYER VI2 ;
  RECT 4.280 21.230 5.140 22.070 ;
  LAYER VI2 ;
  RECT 4.680 21.690 4.880 21.890 ;
  LAYER VI2 ;
  RECT 4.680 21.290 4.880 21.490 ;
  LAYER VI2 ;
  RECT 4.280 21.690 4.480 21.890 ;
  LAYER VI2 ;
  RECT 4.280 21.290 4.480 21.490 ;
  LAYER VI3 ;
  RECT 4.280 18.730 5.140 19.730 ;
  LAYER VI3 ;
  RECT 4.740 19.130 4.940 19.330 ;
  LAYER VI3 ;
  RECT 4.740 18.730 4.940 18.930 ;
  LAYER VI3 ;
  RECT 4.340 19.130 4.540 19.330 ;
  LAYER VI3 ;
  RECT 4.340 18.730 4.540 18.930 ;
  LAYER VI2 ;
  RECT 4.280 18.730 5.140 19.730 ;
  LAYER VI2 ;
  RECT 4.740 19.130 4.940 19.330 ;
  LAYER VI2 ;
  RECT 4.740 18.730 4.940 18.930 ;
  LAYER VI2 ;
  RECT 4.340 19.130 4.540 19.330 ;
  LAYER VI2 ;
  RECT 4.340 18.730 4.540 18.930 ;
  LAYER VI3 ;
  RECT 4.280 14.200 5.140 15.200 ;
  LAYER VI3 ;
  RECT 4.740 14.600 4.940 14.800 ;
  LAYER VI3 ;
  RECT 4.740 14.200 4.940 14.400 ;
  LAYER VI3 ;
  RECT 4.340 14.600 4.540 14.800 ;
  LAYER VI3 ;
  RECT 4.340 14.200 4.540 14.400 ;
  LAYER VI2 ;
  RECT 4.280 14.200 5.140 15.200 ;
  LAYER VI2 ;
  RECT 4.740 14.600 4.940 14.800 ;
  LAYER VI2 ;
  RECT 4.740 14.200 4.940 14.400 ;
  LAYER VI2 ;
  RECT 4.340 14.600 4.540 14.800 ;
  LAYER VI2 ;
  RECT 4.340 14.200 4.540 14.400 ;
  LAYER VI3 ;
  RECT 4.280 9.570 5.140 11.170 ;
  LAYER VI3 ;
  RECT 4.740 10.770 4.940 10.970 ;
  LAYER VI3 ;
  RECT 4.740 10.370 4.940 10.570 ;
  LAYER VI3 ;
  RECT 4.740 9.970 4.940 10.170 ;
  LAYER VI3 ;
  RECT 4.740 9.570 4.940 9.770 ;
  LAYER VI3 ;
  RECT 4.340 10.770 4.540 10.970 ;
  LAYER VI3 ;
  RECT 4.340 10.370 4.540 10.570 ;
  LAYER VI3 ;
  RECT 4.340 9.970 4.540 10.170 ;
  LAYER VI3 ;
  RECT 4.340 9.570 4.540 9.770 ;
  LAYER VI2 ;
  RECT 4.280 9.570 5.140 11.170 ;
  LAYER VI2 ;
  RECT 4.740 10.770 4.940 10.970 ;
  LAYER VI2 ;
  RECT 4.740 10.370 4.940 10.570 ;
  LAYER VI2 ;
  RECT 4.740 9.970 4.940 10.170 ;
  LAYER VI2 ;
  RECT 4.740 9.570 4.940 9.770 ;
  LAYER VI2 ;
  RECT 4.340 10.770 4.540 10.970 ;
  LAYER VI2 ;
  RECT 4.340 10.370 4.540 10.570 ;
  LAYER VI2 ;
  RECT 4.340 9.970 4.540 10.170 ;
  LAYER VI2 ;
  RECT 4.340 9.570 4.540 9.770 ;
  LAYER VI3 ;
  RECT 5.420 5.880 6.560 6.740 ;
  LAYER VI3 ;
  RECT 6.220 6.340 6.420 6.540 ;
  LAYER VI3 ;
  RECT 6.220 5.940 6.420 6.140 ;
  LAYER VI3 ;
  RECT 5.820 6.340 6.020 6.540 ;
  LAYER VI3 ;
  RECT 5.820 5.940 6.020 6.140 ;
  LAYER VI3 ;
  RECT 5.420 6.340 5.620 6.540 ;
  LAYER VI3 ;
  RECT 5.420 5.940 5.620 6.140 ;
  LAYER VI3 ;
  RECT 8.360 5.880 16.360 6.740 ;
  LAYER VI3 ;
  RECT 15.960 6.340 16.160 6.540 ;
  LAYER VI3 ;
  RECT 15.960 5.940 16.160 6.140 ;
  LAYER VI3 ;
  RECT 15.560 6.340 15.760 6.540 ;
  LAYER VI3 ;
  RECT 15.560 5.940 15.760 6.140 ;
  LAYER VI3 ;
  RECT 15.160 6.340 15.360 6.540 ;
  LAYER VI3 ;
  RECT 15.160 5.940 15.360 6.140 ;
  LAYER VI3 ;
  RECT 14.760 6.340 14.960 6.540 ;
  LAYER VI3 ;
  RECT 14.760 5.940 14.960 6.140 ;
  LAYER VI3 ;
  RECT 14.360 6.340 14.560 6.540 ;
  LAYER VI3 ;
  RECT 14.360 5.940 14.560 6.140 ;
  LAYER VI3 ;
  RECT 13.960 6.340 14.160 6.540 ;
  LAYER VI3 ;
  RECT 13.960 5.940 14.160 6.140 ;
  LAYER VI3 ;
  RECT 13.560 6.340 13.760 6.540 ;
  LAYER VI3 ;
  RECT 13.560 5.940 13.760 6.140 ;
  LAYER VI3 ;
  RECT 13.160 6.340 13.360 6.540 ;
  LAYER VI3 ;
  RECT 13.160 5.940 13.360 6.140 ;
  LAYER VI3 ;
  RECT 12.760 6.340 12.960 6.540 ;
  LAYER VI3 ;
  RECT 12.760 5.940 12.960 6.140 ;
  LAYER VI3 ;
  RECT 12.360 6.340 12.560 6.540 ;
  LAYER VI3 ;
  RECT 12.360 5.940 12.560 6.140 ;
  LAYER VI3 ;
  RECT 11.960 6.340 12.160 6.540 ;
  LAYER VI3 ;
  RECT 11.960 5.940 12.160 6.140 ;
  LAYER VI3 ;
  RECT 11.560 6.340 11.760 6.540 ;
  LAYER VI3 ;
  RECT 11.560 5.940 11.760 6.140 ;
  LAYER VI3 ;
  RECT 11.160 6.340 11.360 6.540 ;
  LAYER VI3 ;
  RECT 11.160 5.940 11.360 6.140 ;
  LAYER VI3 ;
  RECT 10.760 6.340 10.960 6.540 ;
  LAYER VI3 ;
  RECT 10.760 5.940 10.960 6.140 ;
  LAYER VI3 ;
  RECT 10.360 6.340 10.560 6.540 ;
  LAYER VI3 ;
  RECT 10.360 5.940 10.560 6.140 ;
  LAYER VI3 ;
  RECT 9.960 6.340 10.160 6.540 ;
  LAYER VI3 ;
  RECT 9.960 5.940 10.160 6.140 ;
  LAYER VI3 ;
  RECT 9.560 6.340 9.760 6.540 ;
  LAYER VI3 ;
  RECT 9.560 5.940 9.760 6.140 ;
  LAYER VI3 ;
  RECT 9.160 6.340 9.360 6.540 ;
  LAYER VI3 ;
  RECT 9.160 5.940 9.360 6.140 ;
  LAYER VI3 ;
  RECT 8.760 6.340 8.960 6.540 ;
  LAYER VI3 ;
  RECT 8.760 5.940 8.960 6.140 ;
  LAYER VI3 ;
  RECT 8.360 6.340 8.560 6.540 ;
  LAYER VI3 ;
  RECT 8.360 5.940 8.560 6.140 ;
  LAYER VI3 ;
  RECT 28.200 5.880 36.200 6.740 ;
  LAYER VI3 ;
  RECT 35.800 6.340 36.000 6.540 ;
  LAYER VI3 ;
  RECT 35.800 5.940 36.000 6.140 ;
  LAYER VI3 ;
  RECT 35.400 6.340 35.600 6.540 ;
  LAYER VI3 ;
  RECT 35.400 5.940 35.600 6.140 ;
  LAYER VI3 ;
  RECT 35.000 6.340 35.200 6.540 ;
  LAYER VI3 ;
  RECT 35.000 5.940 35.200 6.140 ;
  LAYER VI3 ;
  RECT 34.600 6.340 34.800 6.540 ;
  LAYER VI3 ;
  RECT 34.600 5.940 34.800 6.140 ;
  LAYER VI3 ;
  RECT 34.200 6.340 34.400 6.540 ;
  LAYER VI3 ;
  RECT 34.200 5.940 34.400 6.140 ;
  LAYER VI3 ;
  RECT 33.800 6.340 34.000 6.540 ;
  LAYER VI3 ;
  RECT 33.800 5.940 34.000 6.140 ;
  LAYER VI3 ;
  RECT 33.400 6.340 33.600 6.540 ;
  LAYER VI3 ;
  RECT 33.400 5.940 33.600 6.140 ;
  LAYER VI3 ;
  RECT 33.000 6.340 33.200 6.540 ;
  LAYER VI3 ;
  RECT 33.000 5.940 33.200 6.140 ;
  LAYER VI3 ;
  RECT 32.600 6.340 32.800 6.540 ;
  LAYER VI3 ;
  RECT 32.600 5.940 32.800 6.140 ;
  LAYER VI3 ;
  RECT 32.200 6.340 32.400 6.540 ;
  LAYER VI3 ;
  RECT 32.200 5.940 32.400 6.140 ;
  LAYER VI3 ;
  RECT 31.800 6.340 32.000 6.540 ;
  LAYER VI3 ;
  RECT 31.800 5.940 32.000 6.140 ;
  LAYER VI3 ;
  RECT 31.400 6.340 31.600 6.540 ;
  LAYER VI3 ;
  RECT 31.400 5.940 31.600 6.140 ;
  LAYER VI3 ;
  RECT 31.000 6.340 31.200 6.540 ;
  LAYER VI3 ;
  RECT 31.000 5.940 31.200 6.140 ;
  LAYER VI3 ;
  RECT 30.600 6.340 30.800 6.540 ;
  LAYER VI3 ;
  RECT 30.600 5.940 30.800 6.140 ;
  LAYER VI3 ;
  RECT 30.200 6.340 30.400 6.540 ;
  LAYER VI3 ;
  RECT 30.200 5.940 30.400 6.140 ;
  LAYER VI3 ;
  RECT 29.800 6.340 30.000 6.540 ;
  LAYER VI3 ;
  RECT 29.800 5.940 30.000 6.140 ;
  LAYER VI3 ;
  RECT 29.400 6.340 29.600 6.540 ;
  LAYER VI3 ;
  RECT 29.400 5.940 29.600 6.140 ;
  LAYER VI3 ;
  RECT 29.000 6.340 29.200 6.540 ;
  LAYER VI3 ;
  RECT 29.000 5.940 29.200 6.140 ;
  LAYER VI3 ;
  RECT 28.600 6.340 28.800 6.540 ;
  LAYER VI3 ;
  RECT 28.600 5.940 28.800 6.140 ;
  LAYER VI3 ;
  RECT 28.200 6.340 28.400 6.540 ;
  LAYER VI3 ;
  RECT 28.200 5.940 28.400 6.140 ;
  LAYER VI3 ;
  RECT 49.280 5.880 57.280 6.740 ;
  LAYER VI3 ;
  RECT 56.880 6.340 57.080 6.540 ;
  LAYER VI3 ;
  RECT 56.880 5.940 57.080 6.140 ;
  LAYER VI3 ;
  RECT 56.480 6.340 56.680 6.540 ;
  LAYER VI3 ;
  RECT 56.480 5.940 56.680 6.140 ;
  LAYER VI3 ;
  RECT 56.080 6.340 56.280 6.540 ;
  LAYER VI3 ;
  RECT 56.080 5.940 56.280 6.140 ;
  LAYER VI3 ;
  RECT 55.680 6.340 55.880 6.540 ;
  LAYER VI3 ;
  RECT 55.680 5.940 55.880 6.140 ;
  LAYER VI3 ;
  RECT 55.280 6.340 55.480 6.540 ;
  LAYER VI3 ;
  RECT 55.280 5.940 55.480 6.140 ;
  LAYER VI3 ;
  RECT 54.880 6.340 55.080 6.540 ;
  LAYER VI3 ;
  RECT 54.880 5.940 55.080 6.140 ;
  LAYER VI3 ;
  RECT 54.480 6.340 54.680 6.540 ;
  LAYER VI3 ;
  RECT 54.480 5.940 54.680 6.140 ;
  LAYER VI3 ;
  RECT 54.080 6.340 54.280 6.540 ;
  LAYER VI3 ;
  RECT 54.080 5.940 54.280 6.140 ;
  LAYER VI3 ;
  RECT 53.680 6.340 53.880 6.540 ;
  LAYER VI3 ;
  RECT 53.680 5.940 53.880 6.140 ;
  LAYER VI3 ;
  RECT 53.280 6.340 53.480 6.540 ;
  LAYER VI3 ;
  RECT 53.280 5.940 53.480 6.140 ;
  LAYER VI3 ;
  RECT 52.880 6.340 53.080 6.540 ;
  LAYER VI3 ;
  RECT 52.880 5.940 53.080 6.140 ;
  LAYER VI3 ;
  RECT 52.480 6.340 52.680 6.540 ;
  LAYER VI3 ;
  RECT 52.480 5.940 52.680 6.140 ;
  LAYER VI3 ;
  RECT 52.080 6.340 52.280 6.540 ;
  LAYER VI3 ;
  RECT 52.080 5.940 52.280 6.140 ;
  LAYER VI3 ;
  RECT 51.680 6.340 51.880 6.540 ;
  LAYER VI3 ;
  RECT 51.680 5.940 51.880 6.140 ;
  LAYER VI3 ;
  RECT 51.280 6.340 51.480 6.540 ;
  LAYER VI3 ;
  RECT 51.280 5.940 51.480 6.140 ;
  LAYER VI3 ;
  RECT 50.880 6.340 51.080 6.540 ;
  LAYER VI3 ;
  RECT 50.880 5.940 51.080 6.140 ;
  LAYER VI3 ;
  RECT 50.480 6.340 50.680 6.540 ;
  LAYER VI3 ;
  RECT 50.480 5.940 50.680 6.140 ;
  LAYER VI3 ;
  RECT 50.080 6.340 50.280 6.540 ;
  LAYER VI3 ;
  RECT 50.080 5.940 50.280 6.140 ;
  LAYER VI3 ;
  RECT 49.680 6.340 49.880 6.540 ;
  LAYER VI3 ;
  RECT 49.680 5.940 49.880 6.140 ;
  LAYER VI3 ;
  RECT 49.280 6.340 49.480 6.540 ;
  LAYER VI3 ;
  RECT 49.280 5.940 49.480 6.140 ;
  LAYER VI3 ;
  RECT 69.120 5.880 77.120 6.740 ;
  LAYER VI3 ;
  RECT 76.720 6.340 76.920 6.540 ;
  LAYER VI3 ;
  RECT 76.720 5.940 76.920 6.140 ;
  LAYER VI3 ;
  RECT 76.320 6.340 76.520 6.540 ;
  LAYER VI3 ;
  RECT 76.320 5.940 76.520 6.140 ;
  LAYER VI3 ;
  RECT 75.920 6.340 76.120 6.540 ;
  LAYER VI3 ;
  RECT 75.920 5.940 76.120 6.140 ;
  LAYER VI3 ;
  RECT 75.520 6.340 75.720 6.540 ;
  LAYER VI3 ;
  RECT 75.520 5.940 75.720 6.140 ;
  LAYER VI3 ;
  RECT 75.120 6.340 75.320 6.540 ;
  LAYER VI3 ;
  RECT 75.120 5.940 75.320 6.140 ;
  LAYER VI3 ;
  RECT 74.720 6.340 74.920 6.540 ;
  LAYER VI3 ;
  RECT 74.720 5.940 74.920 6.140 ;
  LAYER VI3 ;
  RECT 74.320 6.340 74.520 6.540 ;
  LAYER VI3 ;
  RECT 74.320 5.940 74.520 6.140 ;
  LAYER VI3 ;
  RECT 73.920 6.340 74.120 6.540 ;
  LAYER VI3 ;
  RECT 73.920 5.940 74.120 6.140 ;
  LAYER VI3 ;
  RECT 73.520 6.340 73.720 6.540 ;
  LAYER VI3 ;
  RECT 73.520 5.940 73.720 6.140 ;
  LAYER VI3 ;
  RECT 73.120 6.340 73.320 6.540 ;
  LAYER VI3 ;
  RECT 73.120 5.940 73.320 6.140 ;
  LAYER VI3 ;
  RECT 72.720 6.340 72.920 6.540 ;
  LAYER VI3 ;
  RECT 72.720 5.940 72.920 6.140 ;
  LAYER VI3 ;
  RECT 72.320 6.340 72.520 6.540 ;
  LAYER VI3 ;
  RECT 72.320 5.940 72.520 6.140 ;
  LAYER VI3 ;
  RECT 71.920 6.340 72.120 6.540 ;
  LAYER VI3 ;
  RECT 71.920 5.940 72.120 6.140 ;
  LAYER VI3 ;
  RECT 71.520 6.340 71.720 6.540 ;
  LAYER VI3 ;
  RECT 71.520 5.940 71.720 6.140 ;
  LAYER VI3 ;
  RECT 71.120 6.340 71.320 6.540 ;
  LAYER VI3 ;
  RECT 71.120 5.940 71.320 6.140 ;
  LAYER VI3 ;
  RECT 70.720 6.340 70.920 6.540 ;
  LAYER VI3 ;
  RECT 70.720 5.940 70.920 6.140 ;
  LAYER VI3 ;
  RECT 70.320 6.340 70.520 6.540 ;
  LAYER VI3 ;
  RECT 70.320 5.940 70.520 6.140 ;
  LAYER VI3 ;
  RECT 69.920 6.340 70.120 6.540 ;
  LAYER VI3 ;
  RECT 69.920 5.940 70.120 6.140 ;
  LAYER VI3 ;
  RECT 69.520 6.340 69.720 6.540 ;
  LAYER VI3 ;
  RECT 69.520 5.940 69.720 6.140 ;
  LAYER VI3 ;
  RECT 69.120 6.340 69.320 6.540 ;
  LAYER VI3 ;
  RECT 69.120 5.940 69.320 6.140 ;
  LAYER VI3 ;
  RECT 90.200 5.880 98.200 6.740 ;
  LAYER VI3 ;
  RECT 97.800 6.340 98.000 6.540 ;
  LAYER VI3 ;
  RECT 97.800 5.940 98.000 6.140 ;
  LAYER VI3 ;
  RECT 97.400 6.340 97.600 6.540 ;
  LAYER VI3 ;
  RECT 97.400 5.940 97.600 6.140 ;
  LAYER VI3 ;
  RECT 97.000 6.340 97.200 6.540 ;
  LAYER VI3 ;
  RECT 97.000 5.940 97.200 6.140 ;
  LAYER VI3 ;
  RECT 96.600 6.340 96.800 6.540 ;
  LAYER VI3 ;
  RECT 96.600 5.940 96.800 6.140 ;
  LAYER VI3 ;
  RECT 96.200 6.340 96.400 6.540 ;
  LAYER VI3 ;
  RECT 96.200 5.940 96.400 6.140 ;
  LAYER VI3 ;
  RECT 95.800 6.340 96.000 6.540 ;
  LAYER VI3 ;
  RECT 95.800 5.940 96.000 6.140 ;
  LAYER VI3 ;
  RECT 95.400 6.340 95.600 6.540 ;
  LAYER VI3 ;
  RECT 95.400 5.940 95.600 6.140 ;
  LAYER VI3 ;
  RECT 95.000 6.340 95.200 6.540 ;
  LAYER VI3 ;
  RECT 95.000 5.940 95.200 6.140 ;
  LAYER VI3 ;
  RECT 94.600 6.340 94.800 6.540 ;
  LAYER VI3 ;
  RECT 94.600 5.940 94.800 6.140 ;
  LAYER VI3 ;
  RECT 94.200 6.340 94.400 6.540 ;
  LAYER VI3 ;
  RECT 94.200 5.940 94.400 6.140 ;
  LAYER VI3 ;
  RECT 93.800 6.340 94.000 6.540 ;
  LAYER VI3 ;
  RECT 93.800 5.940 94.000 6.140 ;
  LAYER VI3 ;
  RECT 93.400 6.340 93.600 6.540 ;
  LAYER VI3 ;
  RECT 93.400 5.940 93.600 6.140 ;
  LAYER VI3 ;
  RECT 93.000 6.340 93.200 6.540 ;
  LAYER VI3 ;
  RECT 93.000 5.940 93.200 6.140 ;
  LAYER VI3 ;
  RECT 92.600 6.340 92.800 6.540 ;
  LAYER VI3 ;
  RECT 92.600 5.940 92.800 6.140 ;
  LAYER VI3 ;
  RECT 92.200 6.340 92.400 6.540 ;
  LAYER VI3 ;
  RECT 92.200 5.940 92.400 6.140 ;
  LAYER VI3 ;
  RECT 91.800 6.340 92.000 6.540 ;
  LAYER VI3 ;
  RECT 91.800 5.940 92.000 6.140 ;
  LAYER VI3 ;
  RECT 91.400 6.340 91.600 6.540 ;
  LAYER VI3 ;
  RECT 91.400 5.940 91.600 6.140 ;
  LAYER VI3 ;
  RECT 91.000 6.340 91.200 6.540 ;
  LAYER VI3 ;
  RECT 91.000 5.940 91.200 6.140 ;
  LAYER VI3 ;
  RECT 90.600 6.340 90.800 6.540 ;
  LAYER VI3 ;
  RECT 90.600 5.940 90.800 6.140 ;
  LAYER VI3 ;
  RECT 90.200 6.340 90.400 6.540 ;
  LAYER VI3 ;
  RECT 90.200 5.940 90.400 6.140 ;
  LAYER VI3 ;
  RECT 110.040 5.880 118.040 6.740 ;
  LAYER VI3 ;
  RECT 117.640 6.340 117.840 6.540 ;
  LAYER VI3 ;
  RECT 117.640 5.940 117.840 6.140 ;
  LAYER VI3 ;
  RECT 117.240 6.340 117.440 6.540 ;
  LAYER VI3 ;
  RECT 117.240 5.940 117.440 6.140 ;
  LAYER VI3 ;
  RECT 116.840 6.340 117.040 6.540 ;
  LAYER VI3 ;
  RECT 116.840 5.940 117.040 6.140 ;
  LAYER VI3 ;
  RECT 116.440 6.340 116.640 6.540 ;
  LAYER VI3 ;
  RECT 116.440 5.940 116.640 6.140 ;
  LAYER VI3 ;
  RECT 116.040 6.340 116.240 6.540 ;
  LAYER VI3 ;
  RECT 116.040 5.940 116.240 6.140 ;
  LAYER VI3 ;
  RECT 115.640 6.340 115.840 6.540 ;
  LAYER VI3 ;
  RECT 115.640 5.940 115.840 6.140 ;
  LAYER VI3 ;
  RECT 115.240 6.340 115.440 6.540 ;
  LAYER VI3 ;
  RECT 115.240 5.940 115.440 6.140 ;
  LAYER VI3 ;
  RECT 114.840 6.340 115.040 6.540 ;
  LAYER VI3 ;
  RECT 114.840 5.940 115.040 6.140 ;
  LAYER VI3 ;
  RECT 114.440 6.340 114.640 6.540 ;
  LAYER VI3 ;
  RECT 114.440 5.940 114.640 6.140 ;
  LAYER VI3 ;
  RECT 114.040 6.340 114.240 6.540 ;
  LAYER VI3 ;
  RECT 114.040 5.940 114.240 6.140 ;
  LAYER VI3 ;
  RECT 113.640 6.340 113.840 6.540 ;
  LAYER VI3 ;
  RECT 113.640 5.940 113.840 6.140 ;
  LAYER VI3 ;
  RECT 113.240 6.340 113.440 6.540 ;
  LAYER VI3 ;
  RECT 113.240 5.940 113.440 6.140 ;
  LAYER VI3 ;
  RECT 112.840 6.340 113.040 6.540 ;
  LAYER VI3 ;
  RECT 112.840 5.940 113.040 6.140 ;
  LAYER VI3 ;
  RECT 112.440 6.340 112.640 6.540 ;
  LAYER VI3 ;
  RECT 112.440 5.940 112.640 6.140 ;
  LAYER VI3 ;
  RECT 112.040 6.340 112.240 6.540 ;
  LAYER VI3 ;
  RECT 112.040 5.940 112.240 6.140 ;
  LAYER VI3 ;
  RECT 111.640 6.340 111.840 6.540 ;
  LAYER VI3 ;
  RECT 111.640 5.940 111.840 6.140 ;
  LAYER VI3 ;
  RECT 111.240 6.340 111.440 6.540 ;
  LAYER VI3 ;
  RECT 111.240 5.940 111.440 6.140 ;
  LAYER VI3 ;
  RECT 110.840 6.340 111.040 6.540 ;
  LAYER VI3 ;
  RECT 110.840 5.940 111.040 6.140 ;
  LAYER VI3 ;
  RECT 110.440 6.340 110.640 6.540 ;
  LAYER VI3 ;
  RECT 110.440 5.940 110.640 6.140 ;
  LAYER VI3 ;
  RECT 110.040 6.340 110.240 6.540 ;
  LAYER VI3 ;
  RECT 110.040 5.940 110.240 6.140 ;
  LAYER VI3 ;
  RECT 131.120 5.880 139.120 6.740 ;
  LAYER VI3 ;
  RECT 138.720 6.340 138.920 6.540 ;
  LAYER VI3 ;
  RECT 138.720 5.940 138.920 6.140 ;
  LAYER VI3 ;
  RECT 138.320 6.340 138.520 6.540 ;
  LAYER VI3 ;
  RECT 138.320 5.940 138.520 6.140 ;
  LAYER VI3 ;
  RECT 137.920 6.340 138.120 6.540 ;
  LAYER VI3 ;
  RECT 137.920 5.940 138.120 6.140 ;
  LAYER VI3 ;
  RECT 137.520 6.340 137.720 6.540 ;
  LAYER VI3 ;
  RECT 137.520 5.940 137.720 6.140 ;
  LAYER VI3 ;
  RECT 137.120 6.340 137.320 6.540 ;
  LAYER VI3 ;
  RECT 137.120 5.940 137.320 6.140 ;
  LAYER VI3 ;
  RECT 136.720 6.340 136.920 6.540 ;
  LAYER VI3 ;
  RECT 136.720 5.940 136.920 6.140 ;
  LAYER VI3 ;
  RECT 136.320 6.340 136.520 6.540 ;
  LAYER VI3 ;
  RECT 136.320 5.940 136.520 6.140 ;
  LAYER VI3 ;
  RECT 135.920 6.340 136.120 6.540 ;
  LAYER VI3 ;
  RECT 135.920 5.940 136.120 6.140 ;
  LAYER VI3 ;
  RECT 135.520 6.340 135.720 6.540 ;
  LAYER VI3 ;
  RECT 135.520 5.940 135.720 6.140 ;
  LAYER VI3 ;
  RECT 135.120 6.340 135.320 6.540 ;
  LAYER VI3 ;
  RECT 135.120 5.940 135.320 6.140 ;
  LAYER VI3 ;
  RECT 134.720 6.340 134.920 6.540 ;
  LAYER VI3 ;
  RECT 134.720 5.940 134.920 6.140 ;
  LAYER VI3 ;
  RECT 134.320 6.340 134.520 6.540 ;
  LAYER VI3 ;
  RECT 134.320 5.940 134.520 6.140 ;
  LAYER VI3 ;
  RECT 133.920 6.340 134.120 6.540 ;
  LAYER VI3 ;
  RECT 133.920 5.940 134.120 6.140 ;
  LAYER VI3 ;
  RECT 133.520 6.340 133.720 6.540 ;
  LAYER VI3 ;
  RECT 133.520 5.940 133.720 6.140 ;
  LAYER VI3 ;
  RECT 133.120 6.340 133.320 6.540 ;
  LAYER VI3 ;
  RECT 133.120 5.940 133.320 6.140 ;
  LAYER VI3 ;
  RECT 132.720 6.340 132.920 6.540 ;
  LAYER VI3 ;
  RECT 132.720 5.940 132.920 6.140 ;
  LAYER VI3 ;
  RECT 132.320 6.340 132.520 6.540 ;
  LAYER VI3 ;
  RECT 132.320 5.940 132.520 6.140 ;
  LAYER VI3 ;
  RECT 131.920 6.340 132.120 6.540 ;
  LAYER VI3 ;
  RECT 131.920 5.940 132.120 6.140 ;
  LAYER VI3 ;
  RECT 131.520 6.340 131.720 6.540 ;
  LAYER VI3 ;
  RECT 131.520 5.940 131.720 6.140 ;
  LAYER VI3 ;
  RECT 131.120 6.340 131.320 6.540 ;
  LAYER VI3 ;
  RECT 131.120 5.940 131.320 6.140 ;
  LAYER VI3 ;
  RECT 150.960 5.880 158.960 6.740 ;
  LAYER VI3 ;
  RECT 158.560 6.340 158.760 6.540 ;
  LAYER VI3 ;
  RECT 158.560 5.940 158.760 6.140 ;
  LAYER VI3 ;
  RECT 158.160 6.340 158.360 6.540 ;
  LAYER VI3 ;
  RECT 158.160 5.940 158.360 6.140 ;
  LAYER VI3 ;
  RECT 157.760 6.340 157.960 6.540 ;
  LAYER VI3 ;
  RECT 157.760 5.940 157.960 6.140 ;
  LAYER VI3 ;
  RECT 157.360 6.340 157.560 6.540 ;
  LAYER VI3 ;
  RECT 157.360 5.940 157.560 6.140 ;
  LAYER VI3 ;
  RECT 156.960 6.340 157.160 6.540 ;
  LAYER VI3 ;
  RECT 156.960 5.940 157.160 6.140 ;
  LAYER VI3 ;
  RECT 156.560 6.340 156.760 6.540 ;
  LAYER VI3 ;
  RECT 156.560 5.940 156.760 6.140 ;
  LAYER VI3 ;
  RECT 156.160 6.340 156.360 6.540 ;
  LAYER VI3 ;
  RECT 156.160 5.940 156.360 6.140 ;
  LAYER VI3 ;
  RECT 155.760 6.340 155.960 6.540 ;
  LAYER VI3 ;
  RECT 155.760 5.940 155.960 6.140 ;
  LAYER VI3 ;
  RECT 155.360 6.340 155.560 6.540 ;
  LAYER VI3 ;
  RECT 155.360 5.940 155.560 6.140 ;
  LAYER VI3 ;
  RECT 154.960 6.340 155.160 6.540 ;
  LAYER VI3 ;
  RECT 154.960 5.940 155.160 6.140 ;
  LAYER VI3 ;
  RECT 154.560 6.340 154.760 6.540 ;
  LAYER VI3 ;
  RECT 154.560 5.940 154.760 6.140 ;
  LAYER VI3 ;
  RECT 154.160 6.340 154.360 6.540 ;
  LAYER VI3 ;
  RECT 154.160 5.940 154.360 6.140 ;
  LAYER VI3 ;
  RECT 153.760 6.340 153.960 6.540 ;
  LAYER VI3 ;
  RECT 153.760 5.940 153.960 6.140 ;
  LAYER VI3 ;
  RECT 153.360 6.340 153.560 6.540 ;
  LAYER VI3 ;
  RECT 153.360 5.940 153.560 6.140 ;
  LAYER VI3 ;
  RECT 152.960 6.340 153.160 6.540 ;
  LAYER VI3 ;
  RECT 152.960 5.940 153.160 6.140 ;
  LAYER VI3 ;
  RECT 152.560 6.340 152.760 6.540 ;
  LAYER VI3 ;
  RECT 152.560 5.940 152.760 6.140 ;
  LAYER VI3 ;
  RECT 152.160 6.340 152.360 6.540 ;
  LAYER VI3 ;
  RECT 152.160 5.940 152.360 6.140 ;
  LAYER VI3 ;
  RECT 151.760 6.340 151.960 6.540 ;
  LAYER VI3 ;
  RECT 151.760 5.940 151.960 6.140 ;
  LAYER VI3 ;
  RECT 151.360 6.340 151.560 6.540 ;
  LAYER VI3 ;
  RECT 151.360 5.940 151.560 6.140 ;
  LAYER VI3 ;
  RECT 150.960 6.340 151.160 6.540 ;
  LAYER VI3 ;
  RECT 150.960 5.940 151.160 6.140 ;
  LAYER VI3 ;
  RECT 172.040 5.880 180.040 6.740 ;
  LAYER VI3 ;
  RECT 179.640 6.340 179.840 6.540 ;
  LAYER VI3 ;
  RECT 179.640 5.940 179.840 6.140 ;
  LAYER VI3 ;
  RECT 179.240 6.340 179.440 6.540 ;
  LAYER VI3 ;
  RECT 179.240 5.940 179.440 6.140 ;
  LAYER VI3 ;
  RECT 178.840 6.340 179.040 6.540 ;
  LAYER VI3 ;
  RECT 178.840 5.940 179.040 6.140 ;
  LAYER VI3 ;
  RECT 178.440 6.340 178.640 6.540 ;
  LAYER VI3 ;
  RECT 178.440 5.940 178.640 6.140 ;
  LAYER VI3 ;
  RECT 178.040 6.340 178.240 6.540 ;
  LAYER VI3 ;
  RECT 178.040 5.940 178.240 6.140 ;
  LAYER VI3 ;
  RECT 177.640 6.340 177.840 6.540 ;
  LAYER VI3 ;
  RECT 177.640 5.940 177.840 6.140 ;
  LAYER VI3 ;
  RECT 177.240 6.340 177.440 6.540 ;
  LAYER VI3 ;
  RECT 177.240 5.940 177.440 6.140 ;
  LAYER VI3 ;
  RECT 176.840 6.340 177.040 6.540 ;
  LAYER VI3 ;
  RECT 176.840 5.940 177.040 6.140 ;
  LAYER VI3 ;
  RECT 176.440 6.340 176.640 6.540 ;
  LAYER VI3 ;
  RECT 176.440 5.940 176.640 6.140 ;
  LAYER VI3 ;
  RECT 176.040 6.340 176.240 6.540 ;
  LAYER VI3 ;
  RECT 176.040 5.940 176.240 6.140 ;
  LAYER VI3 ;
  RECT 175.640 6.340 175.840 6.540 ;
  LAYER VI3 ;
  RECT 175.640 5.940 175.840 6.140 ;
  LAYER VI3 ;
  RECT 175.240 6.340 175.440 6.540 ;
  LAYER VI3 ;
  RECT 175.240 5.940 175.440 6.140 ;
  LAYER VI3 ;
  RECT 174.840 6.340 175.040 6.540 ;
  LAYER VI3 ;
  RECT 174.840 5.940 175.040 6.140 ;
  LAYER VI3 ;
  RECT 174.440 6.340 174.640 6.540 ;
  LAYER VI3 ;
  RECT 174.440 5.940 174.640 6.140 ;
  LAYER VI3 ;
  RECT 174.040 6.340 174.240 6.540 ;
  LAYER VI3 ;
  RECT 174.040 5.940 174.240 6.140 ;
  LAYER VI3 ;
  RECT 173.640 6.340 173.840 6.540 ;
  LAYER VI3 ;
  RECT 173.640 5.940 173.840 6.140 ;
  LAYER VI3 ;
  RECT 173.240 6.340 173.440 6.540 ;
  LAYER VI3 ;
  RECT 173.240 5.940 173.440 6.140 ;
  LAYER VI3 ;
  RECT 172.840 6.340 173.040 6.540 ;
  LAYER VI3 ;
  RECT 172.840 5.940 173.040 6.140 ;
  LAYER VI3 ;
  RECT 172.440 6.340 172.640 6.540 ;
  LAYER VI3 ;
  RECT 172.440 5.940 172.640 6.140 ;
  LAYER VI3 ;
  RECT 172.040 6.340 172.240 6.540 ;
  LAYER VI3 ;
  RECT 172.040 5.940 172.240 6.140 ;
  LAYER VI3 ;
  RECT 191.880 5.880 199.880 6.740 ;
  LAYER VI3 ;
  RECT 199.480 6.340 199.680 6.540 ;
  LAYER VI3 ;
  RECT 199.480 5.940 199.680 6.140 ;
  LAYER VI3 ;
  RECT 199.080 6.340 199.280 6.540 ;
  LAYER VI3 ;
  RECT 199.080 5.940 199.280 6.140 ;
  LAYER VI3 ;
  RECT 198.680 6.340 198.880 6.540 ;
  LAYER VI3 ;
  RECT 198.680 5.940 198.880 6.140 ;
  LAYER VI3 ;
  RECT 198.280 6.340 198.480 6.540 ;
  LAYER VI3 ;
  RECT 198.280 5.940 198.480 6.140 ;
  LAYER VI3 ;
  RECT 197.880 6.340 198.080 6.540 ;
  LAYER VI3 ;
  RECT 197.880 5.940 198.080 6.140 ;
  LAYER VI3 ;
  RECT 197.480 6.340 197.680 6.540 ;
  LAYER VI3 ;
  RECT 197.480 5.940 197.680 6.140 ;
  LAYER VI3 ;
  RECT 197.080 6.340 197.280 6.540 ;
  LAYER VI3 ;
  RECT 197.080 5.940 197.280 6.140 ;
  LAYER VI3 ;
  RECT 196.680 6.340 196.880 6.540 ;
  LAYER VI3 ;
  RECT 196.680 5.940 196.880 6.140 ;
  LAYER VI3 ;
  RECT 196.280 6.340 196.480 6.540 ;
  LAYER VI3 ;
  RECT 196.280 5.940 196.480 6.140 ;
  LAYER VI3 ;
  RECT 195.880 6.340 196.080 6.540 ;
  LAYER VI3 ;
  RECT 195.880 5.940 196.080 6.140 ;
  LAYER VI3 ;
  RECT 195.480 6.340 195.680 6.540 ;
  LAYER VI3 ;
  RECT 195.480 5.940 195.680 6.140 ;
  LAYER VI3 ;
  RECT 195.080 6.340 195.280 6.540 ;
  LAYER VI3 ;
  RECT 195.080 5.940 195.280 6.140 ;
  LAYER VI3 ;
  RECT 194.680 6.340 194.880 6.540 ;
  LAYER VI3 ;
  RECT 194.680 5.940 194.880 6.140 ;
  LAYER VI3 ;
  RECT 194.280 6.340 194.480 6.540 ;
  LAYER VI3 ;
  RECT 194.280 5.940 194.480 6.140 ;
  LAYER VI3 ;
  RECT 193.880 6.340 194.080 6.540 ;
  LAYER VI3 ;
  RECT 193.880 5.940 194.080 6.140 ;
  LAYER VI3 ;
  RECT 193.480 6.340 193.680 6.540 ;
  LAYER VI3 ;
  RECT 193.480 5.940 193.680 6.140 ;
  LAYER VI3 ;
  RECT 193.080 6.340 193.280 6.540 ;
  LAYER VI3 ;
  RECT 193.080 5.940 193.280 6.140 ;
  LAYER VI3 ;
  RECT 192.680 6.340 192.880 6.540 ;
  LAYER VI3 ;
  RECT 192.680 5.940 192.880 6.140 ;
  LAYER VI3 ;
  RECT 192.280 6.340 192.480 6.540 ;
  LAYER VI3 ;
  RECT 192.280 5.940 192.480 6.140 ;
  LAYER VI3 ;
  RECT 191.880 6.340 192.080 6.540 ;
  LAYER VI3 ;
  RECT 191.880 5.940 192.080 6.140 ;
  LAYER VI3 ;
  RECT 212.960 5.880 220.960 6.740 ;
  LAYER VI3 ;
  RECT 220.560 6.340 220.760 6.540 ;
  LAYER VI3 ;
  RECT 220.560 5.940 220.760 6.140 ;
  LAYER VI3 ;
  RECT 220.160 6.340 220.360 6.540 ;
  LAYER VI3 ;
  RECT 220.160 5.940 220.360 6.140 ;
  LAYER VI3 ;
  RECT 219.760 6.340 219.960 6.540 ;
  LAYER VI3 ;
  RECT 219.760 5.940 219.960 6.140 ;
  LAYER VI3 ;
  RECT 219.360 6.340 219.560 6.540 ;
  LAYER VI3 ;
  RECT 219.360 5.940 219.560 6.140 ;
  LAYER VI3 ;
  RECT 218.960 6.340 219.160 6.540 ;
  LAYER VI3 ;
  RECT 218.960 5.940 219.160 6.140 ;
  LAYER VI3 ;
  RECT 218.560 6.340 218.760 6.540 ;
  LAYER VI3 ;
  RECT 218.560 5.940 218.760 6.140 ;
  LAYER VI3 ;
  RECT 218.160 6.340 218.360 6.540 ;
  LAYER VI3 ;
  RECT 218.160 5.940 218.360 6.140 ;
  LAYER VI3 ;
  RECT 217.760 6.340 217.960 6.540 ;
  LAYER VI3 ;
  RECT 217.760 5.940 217.960 6.140 ;
  LAYER VI3 ;
  RECT 217.360 6.340 217.560 6.540 ;
  LAYER VI3 ;
  RECT 217.360 5.940 217.560 6.140 ;
  LAYER VI3 ;
  RECT 216.960 6.340 217.160 6.540 ;
  LAYER VI3 ;
  RECT 216.960 5.940 217.160 6.140 ;
  LAYER VI3 ;
  RECT 216.560 6.340 216.760 6.540 ;
  LAYER VI3 ;
  RECT 216.560 5.940 216.760 6.140 ;
  LAYER VI3 ;
  RECT 216.160 6.340 216.360 6.540 ;
  LAYER VI3 ;
  RECT 216.160 5.940 216.360 6.140 ;
  LAYER VI3 ;
  RECT 215.760 6.340 215.960 6.540 ;
  LAYER VI3 ;
  RECT 215.760 5.940 215.960 6.140 ;
  LAYER VI3 ;
  RECT 215.360 6.340 215.560 6.540 ;
  LAYER VI3 ;
  RECT 215.360 5.940 215.560 6.140 ;
  LAYER VI3 ;
  RECT 214.960 6.340 215.160 6.540 ;
  LAYER VI3 ;
  RECT 214.960 5.940 215.160 6.140 ;
  LAYER VI3 ;
  RECT 214.560 6.340 214.760 6.540 ;
  LAYER VI3 ;
  RECT 214.560 5.940 214.760 6.140 ;
  LAYER VI3 ;
  RECT 214.160 6.340 214.360 6.540 ;
  LAYER VI3 ;
  RECT 214.160 5.940 214.360 6.140 ;
  LAYER VI3 ;
  RECT 213.760 6.340 213.960 6.540 ;
  LAYER VI3 ;
  RECT 213.760 5.940 213.960 6.140 ;
  LAYER VI3 ;
  RECT 213.360 6.340 213.560 6.540 ;
  LAYER VI3 ;
  RECT 213.360 5.940 213.560 6.140 ;
  LAYER VI3 ;
  RECT 212.960 6.340 213.160 6.540 ;
  LAYER VI3 ;
  RECT 212.960 5.940 213.160 6.140 ;
  LAYER VI3 ;
  RECT 232.800 5.880 240.800 6.740 ;
  LAYER VI3 ;
  RECT 240.400 6.340 240.600 6.540 ;
  LAYER VI3 ;
  RECT 240.400 5.940 240.600 6.140 ;
  LAYER VI3 ;
  RECT 240.000 6.340 240.200 6.540 ;
  LAYER VI3 ;
  RECT 240.000 5.940 240.200 6.140 ;
  LAYER VI3 ;
  RECT 239.600 6.340 239.800 6.540 ;
  LAYER VI3 ;
  RECT 239.600 5.940 239.800 6.140 ;
  LAYER VI3 ;
  RECT 239.200 6.340 239.400 6.540 ;
  LAYER VI3 ;
  RECT 239.200 5.940 239.400 6.140 ;
  LAYER VI3 ;
  RECT 238.800 6.340 239.000 6.540 ;
  LAYER VI3 ;
  RECT 238.800 5.940 239.000 6.140 ;
  LAYER VI3 ;
  RECT 238.400 6.340 238.600 6.540 ;
  LAYER VI3 ;
  RECT 238.400 5.940 238.600 6.140 ;
  LAYER VI3 ;
  RECT 238.000 6.340 238.200 6.540 ;
  LAYER VI3 ;
  RECT 238.000 5.940 238.200 6.140 ;
  LAYER VI3 ;
  RECT 237.600 6.340 237.800 6.540 ;
  LAYER VI3 ;
  RECT 237.600 5.940 237.800 6.140 ;
  LAYER VI3 ;
  RECT 237.200 6.340 237.400 6.540 ;
  LAYER VI3 ;
  RECT 237.200 5.940 237.400 6.140 ;
  LAYER VI3 ;
  RECT 236.800 6.340 237.000 6.540 ;
  LAYER VI3 ;
  RECT 236.800 5.940 237.000 6.140 ;
  LAYER VI3 ;
  RECT 236.400 6.340 236.600 6.540 ;
  LAYER VI3 ;
  RECT 236.400 5.940 236.600 6.140 ;
  LAYER VI3 ;
  RECT 236.000 6.340 236.200 6.540 ;
  LAYER VI3 ;
  RECT 236.000 5.940 236.200 6.140 ;
  LAYER VI3 ;
  RECT 235.600 6.340 235.800 6.540 ;
  LAYER VI3 ;
  RECT 235.600 5.940 235.800 6.140 ;
  LAYER VI3 ;
  RECT 235.200 6.340 235.400 6.540 ;
  LAYER VI3 ;
  RECT 235.200 5.940 235.400 6.140 ;
  LAYER VI3 ;
  RECT 234.800 6.340 235.000 6.540 ;
  LAYER VI3 ;
  RECT 234.800 5.940 235.000 6.140 ;
  LAYER VI3 ;
  RECT 234.400 6.340 234.600 6.540 ;
  LAYER VI3 ;
  RECT 234.400 5.940 234.600 6.140 ;
  LAYER VI3 ;
  RECT 234.000 6.340 234.200 6.540 ;
  LAYER VI3 ;
  RECT 234.000 5.940 234.200 6.140 ;
  LAYER VI3 ;
  RECT 233.600 6.340 233.800 6.540 ;
  LAYER VI3 ;
  RECT 233.600 5.940 233.800 6.140 ;
  LAYER VI3 ;
  RECT 233.200 6.340 233.400 6.540 ;
  LAYER VI3 ;
  RECT 233.200 5.940 233.400 6.140 ;
  LAYER VI3 ;
  RECT 232.800 6.340 233.000 6.540 ;
  LAYER VI3 ;
  RECT 232.800 5.940 233.000 6.140 ;
  LAYER VI3 ;
  RECT 253.880 5.880 261.880 6.740 ;
  LAYER VI3 ;
  RECT 261.480 6.340 261.680 6.540 ;
  LAYER VI3 ;
  RECT 261.480 5.940 261.680 6.140 ;
  LAYER VI3 ;
  RECT 261.080 6.340 261.280 6.540 ;
  LAYER VI3 ;
  RECT 261.080 5.940 261.280 6.140 ;
  LAYER VI3 ;
  RECT 260.680 6.340 260.880 6.540 ;
  LAYER VI3 ;
  RECT 260.680 5.940 260.880 6.140 ;
  LAYER VI3 ;
  RECT 260.280 6.340 260.480 6.540 ;
  LAYER VI3 ;
  RECT 260.280 5.940 260.480 6.140 ;
  LAYER VI3 ;
  RECT 259.880 6.340 260.080 6.540 ;
  LAYER VI3 ;
  RECT 259.880 5.940 260.080 6.140 ;
  LAYER VI3 ;
  RECT 259.480 6.340 259.680 6.540 ;
  LAYER VI3 ;
  RECT 259.480 5.940 259.680 6.140 ;
  LAYER VI3 ;
  RECT 259.080 6.340 259.280 6.540 ;
  LAYER VI3 ;
  RECT 259.080 5.940 259.280 6.140 ;
  LAYER VI3 ;
  RECT 258.680 6.340 258.880 6.540 ;
  LAYER VI3 ;
  RECT 258.680 5.940 258.880 6.140 ;
  LAYER VI3 ;
  RECT 258.280 6.340 258.480 6.540 ;
  LAYER VI3 ;
  RECT 258.280 5.940 258.480 6.140 ;
  LAYER VI3 ;
  RECT 257.880 6.340 258.080 6.540 ;
  LAYER VI3 ;
  RECT 257.880 5.940 258.080 6.140 ;
  LAYER VI3 ;
  RECT 257.480 6.340 257.680 6.540 ;
  LAYER VI3 ;
  RECT 257.480 5.940 257.680 6.140 ;
  LAYER VI3 ;
  RECT 257.080 6.340 257.280 6.540 ;
  LAYER VI3 ;
  RECT 257.080 5.940 257.280 6.140 ;
  LAYER VI3 ;
  RECT 256.680 6.340 256.880 6.540 ;
  LAYER VI3 ;
  RECT 256.680 5.940 256.880 6.140 ;
  LAYER VI3 ;
  RECT 256.280 6.340 256.480 6.540 ;
  LAYER VI3 ;
  RECT 256.280 5.940 256.480 6.140 ;
  LAYER VI3 ;
  RECT 255.880 6.340 256.080 6.540 ;
  LAYER VI3 ;
  RECT 255.880 5.940 256.080 6.140 ;
  LAYER VI3 ;
  RECT 255.480 6.340 255.680 6.540 ;
  LAYER VI3 ;
  RECT 255.480 5.940 255.680 6.140 ;
  LAYER VI3 ;
  RECT 255.080 6.340 255.280 6.540 ;
  LAYER VI3 ;
  RECT 255.080 5.940 255.280 6.140 ;
  LAYER VI3 ;
  RECT 254.680 6.340 254.880 6.540 ;
  LAYER VI3 ;
  RECT 254.680 5.940 254.880 6.140 ;
  LAYER VI3 ;
  RECT 254.280 6.340 254.480 6.540 ;
  LAYER VI3 ;
  RECT 254.280 5.940 254.480 6.140 ;
  LAYER VI3 ;
  RECT 253.880 6.340 254.080 6.540 ;
  LAYER VI3 ;
  RECT 253.880 5.940 254.080 6.140 ;
  LAYER VI3 ;
  RECT 273.720 5.880 281.720 6.740 ;
  LAYER VI3 ;
  RECT 281.320 6.340 281.520 6.540 ;
  LAYER VI3 ;
  RECT 281.320 5.940 281.520 6.140 ;
  LAYER VI3 ;
  RECT 280.920 6.340 281.120 6.540 ;
  LAYER VI3 ;
  RECT 280.920 5.940 281.120 6.140 ;
  LAYER VI3 ;
  RECT 280.520 6.340 280.720 6.540 ;
  LAYER VI3 ;
  RECT 280.520 5.940 280.720 6.140 ;
  LAYER VI3 ;
  RECT 280.120 6.340 280.320 6.540 ;
  LAYER VI3 ;
  RECT 280.120 5.940 280.320 6.140 ;
  LAYER VI3 ;
  RECT 279.720 6.340 279.920 6.540 ;
  LAYER VI3 ;
  RECT 279.720 5.940 279.920 6.140 ;
  LAYER VI3 ;
  RECT 279.320 6.340 279.520 6.540 ;
  LAYER VI3 ;
  RECT 279.320 5.940 279.520 6.140 ;
  LAYER VI3 ;
  RECT 278.920 6.340 279.120 6.540 ;
  LAYER VI3 ;
  RECT 278.920 5.940 279.120 6.140 ;
  LAYER VI3 ;
  RECT 278.520 6.340 278.720 6.540 ;
  LAYER VI3 ;
  RECT 278.520 5.940 278.720 6.140 ;
  LAYER VI3 ;
  RECT 278.120 6.340 278.320 6.540 ;
  LAYER VI3 ;
  RECT 278.120 5.940 278.320 6.140 ;
  LAYER VI3 ;
  RECT 277.720 6.340 277.920 6.540 ;
  LAYER VI3 ;
  RECT 277.720 5.940 277.920 6.140 ;
  LAYER VI3 ;
  RECT 277.320 6.340 277.520 6.540 ;
  LAYER VI3 ;
  RECT 277.320 5.940 277.520 6.140 ;
  LAYER VI3 ;
  RECT 276.920 6.340 277.120 6.540 ;
  LAYER VI3 ;
  RECT 276.920 5.940 277.120 6.140 ;
  LAYER VI3 ;
  RECT 276.520 6.340 276.720 6.540 ;
  LAYER VI3 ;
  RECT 276.520 5.940 276.720 6.140 ;
  LAYER VI3 ;
  RECT 276.120 6.340 276.320 6.540 ;
  LAYER VI3 ;
  RECT 276.120 5.940 276.320 6.140 ;
  LAYER VI3 ;
  RECT 275.720 6.340 275.920 6.540 ;
  LAYER VI3 ;
  RECT 275.720 5.940 275.920 6.140 ;
  LAYER VI3 ;
  RECT 275.320 6.340 275.520 6.540 ;
  LAYER VI3 ;
  RECT 275.320 5.940 275.520 6.140 ;
  LAYER VI3 ;
  RECT 274.920 6.340 275.120 6.540 ;
  LAYER VI3 ;
  RECT 274.920 5.940 275.120 6.140 ;
  LAYER VI3 ;
  RECT 274.520 6.340 274.720 6.540 ;
  LAYER VI3 ;
  RECT 274.520 5.940 274.720 6.140 ;
  LAYER VI3 ;
  RECT 274.120 6.340 274.320 6.540 ;
  LAYER VI3 ;
  RECT 274.120 5.940 274.320 6.140 ;
  LAYER VI3 ;
  RECT 273.720 6.340 273.920 6.540 ;
  LAYER VI3 ;
  RECT 273.720 5.940 273.920 6.140 ;
  LAYER VI3 ;
  RECT 294.800 5.880 302.800 6.740 ;
  LAYER VI3 ;
  RECT 302.400 6.340 302.600 6.540 ;
  LAYER VI3 ;
  RECT 302.400 5.940 302.600 6.140 ;
  LAYER VI3 ;
  RECT 302.000 6.340 302.200 6.540 ;
  LAYER VI3 ;
  RECT 302.000 5.940 302.200 6.140 ;
  LAYER VI3 ;
  RECT 301.600 6.340 301.800 6.540 ;
  LAYER VI3 ;
  RECT 301.600 5.940 301.800 6.140 ;
  LAYER VI3 ;
  RECT 301.200 6.340 301.400 6.540 ;
  LAYER VI3 ;
  RECT 301.200 5.940 301.400 6.140 ;
  LAYER VI3 ;
  RECT 300.800 6.340 301.000 6.540 ;
  LAYER VI3 ;
  RECT 300.800 5.940 301.000 6.140 ;
  LAYER VI3 ;
  RECT 300.400 6.340 300.600 6.540 ;
  LAYER VI3 ;
  RECT 300.400 5.940 300.600 6.140 ;
  LAYER VI3 ;
  RECT 300.000 6.340 300.200 6.540 ;
  LAYER VI3 ;
  RECT 300.000 5.940 300.200 6.140 ;
  LAYER VI3 ;
  RECT 299.600 6.340 299.800 6.540 ;
  LAYER VI3 ;
  RECT 299.600 5.940 299.800 6.140 ;
  LAYER VI3 ;
  RECT 299.200 6.340 299.400 6.540 ;
  LAYER VI3 ;
  RECT 299.200 5.940 299.400 6.140 ;
  LAYER VI3 ;
  RECT 298.800 6.340 299.000 6.540 ;
  LAYER VI3 ;
  RECT 298.800 5.940 299.000 6.140 ;
  LAYER VI3 ;
  RECT 298.400 6.340 298.600 6.540 ;
  LAYER VI3 ;
  RECT 298.400 5.940 298.600 6.140 ;
  LAYER VI3 ;
  RECT 298.000 6.340 298.200 6.540 ;
  LAYER VI3 ;
  RECT 298.000 5.940 298.200 6.140 ;
  LAYER VI3 ;
  RECT 297.600 6.340 297.800 6.540 ;
  LAYER VI3 ;
  RECT 297.600 5.940 297.800 6.140 ;
  LAYER VI3 ;
  RECT 297.200 6.340 297.400 6.540 ;
  LAYER VI3 ;
  RECT 297.200 5.940 297.400 6.140 ;
  LAYER VI3 ;
  RECT 296.800 6.340 297.000 6.540 ;
  LAYER VI3 ;
  RECT 296.800 5.940 297.000 6.140 ;
  LAYER VI3 ;
  RECT 296.400 6.340 296.600 6.540 ;
  LAYER VI3 ;
  RECT 296.400 5.940 296.600 6.140 ;
  LAYER VI3 ;
  RECT 296.000 6.340 296.200 6.540 ;
  LAYER VI3 ;
  RECT 296.000 5.940 296.200 6.140 ;
  LAYER VI3 ;
  RECT 295.600 6.340 295.800 6.540 ;
  LAYER VI3 ;
  RECT 295.600 5.940 295.800 6.140 ;
  LAYER VI3 ;
  RECT 295.200 6.340 295.400 6.540 ;
  LAYER VI3 ;
  RECT 295.200 5.940 295.400 6.140 ;
  LAYER VI3 ;
  RECT 294.800 6.340 295.000 6.540 ;
  LAYER VI3 ;
  RECT 294.800 5.940 295.000 6.140 ;
  LAYER VI3 ;
  RECT 314.640 5.880 322.640 6.740 ;
  LAYER VI3 ;
  RECT 322.240 6.340 322.440 6.540 ;
  LAYER VI3 ;
  RECT 322.240 5.940 322.440 6.140 ;
  LAYER VI3 ;
  RECT 321.840 6.340 322.040 6.540 ;
  LAYER VI3 ;
  RECT 321.840 5.940 322.040 6.140 ;
  LAYER VI3 ;
  RECT 321.440 6.340 321.640 6.540 ;
  LAYER VI3 ;
  RECT 321.440 5.940 321.640 6.140 ;
  LAYER VI3 ;
  RECT 321.040 6.340 321.240 6.540 ;
  LAYER VI3 ;
  RECT 321.040 5.940 321.240 6.140 ;
  LAYER VI3 ;
  RECT 320.640 6.340 320.840 6.540 ;
  LAYER VI3 ;
  RECT 320.640 5.940 320.840 6.140 ;
  LAYER VI3 ;
  RECT 320.240 6.340 320.440 6.540 ;
  LAYER VI3 ;
  RECT 320.240 5.940 320.440 6.140 ;
  LAYER VI3 ;
  RECT 319.840 6.340 320.040 6.540 ;
  LAYER VI3 ;
  RECT 319.840 5.940 320.040 6.140 ;
  LAYER VI3 ;
  RECT 319.440 6.340 319.640 6.540 ;
  LAYER VI3 ;
  RECT 319.440 5.940 319.640 6.140 ;
  LAYER VI3 ;
  RECT 319.040 6.340 319.240 6.540 ;
  LAYER VI3 ;
  RECT 319.040 5.940 319.240 6.140 ;
  LAYER VI3 ;
  RECT 318.640 6.340 318.840 6.540 ;
  LAYER VI3 ;
  RECT 318.640 5.940 318.840 6.140 ;
  LAYER VI3 ;
  RECT 318.240 6.340 318.440 6.540 ;
  LAYER VI3 ;
  RECT 318.240 5.940 318.440 6.140 ;
  LAYER VI3 ;
  RECT 317.840 6.340 318.040 6.540 ;
  LAYER VI3 ;
  RECT 317.840 5.940 318.040 6.140 ;
  LAYER VI3 ;
  RECT 317.440 6.340 317.640 6.540 ;
  LAYER VI3 ;
  RECT 317.440 5.940 317.640 6.140 ;
  LAYER VI3 ;
  RECT 317.040 6.340 317.240 6.540 ;
  LAYER VI3 ;
  RECT 317.040 5.940 317.240 6.140 ;
  LAYER VI3 ;
  RECT 316.640 6.340 316.840 6.540 ;
  LAYER VI3 ;
  RECT 316.640 5.940 316.840 6.140 ;
  LAYER VI3 ;
  RECT 316.240 6.340 316.440 6.540 ;
  LAYER VI3 ;
  RECT 316.240 5.940 316.440 6.140 ;
  LAYER VI3 ;
  RECT 315.840 6.340 316.040 6.540 ;
  LAYER VI3 ;
  RECT 315.840 5.940 316.040 6.140 ;
  LAYER VI3 ;
  RECT 315.440 6.340 315.640 6.540 ;
  LAYER VI3 ;
  RECT 315.440 5.940 315.640 6.140 ;
  LAYER VI3 ;
  RECT 315.040 6.340 315.240 6.540 ;
  LAYER VI3 ;
  RECT 315.040 5.940 315.240 6.140 ;
  LAYER VI3 ;
  RECT 314.640 6.340 314.840 6.540 ;
  LAYER VI3 ;
  RECT 314.640 5.940 314.840 6.140 ;
  LAYER VI3 ;
  RECT 335.720 5.880 343.720 6.740 ;
  LAYER VI3 ;
  RECT 343.320 6.340 343.520 6.540 ;
  LAYER VI3 ;
  RECT 343.320 5.940 343.520 6.140 ;
  LAYER VI3 ;
  RECT 342.920 6.340 343.120 6.540 ;
  LAYER VI3 ;
  RECT 342.920 5.940 343.120 6.140 ;
  LAYER VI3 ;
  RECT 342.520 6.340 342.720 6.540 ;
  LAYER VI3 ;
  RECT 342.520 5.940 342.720 6.140 ;
  LAYER VI3 ;
  RECT 342.120 6.340 342.320 6.540 ;
  LAYER VI3 ;
  RECT 342.120 5.940 342.320 6.140 ;
  LAYER VI3 ;
  RECT 341.720 6.340 341.920 6.540 ;
  LAYER VI3 ;
  RECT 341.720 5.940 341.920 6.140 ;
  LAYER VI3 ;
  RECT 341.320 6.340 341.520 6.540 ;
  LAYER VI3 ;
  RECT 341.320 5.940 341.520 6.140 ;
  LAYER VI3 ;
  RECT 340.920 6.340 341.120 6.540 ;
  LAYER VI3 ;
  RECT 340.920 5.940 341.120 6.140 ;
  LAYER VI3 ;
  RECT 340.520 6.340 340.720 6.540 ;
  LAYER VI3 ;
  RECT 340.520 5.940 340.720 6.140 ;
  LAYER VI3 ;
  RECT 340.120 6.340 340.320 6.540 ;
  LAYER VI3 ;
  RECT 340.120 5.940 340.320 6.140 ;
  LAYER VI3 ;
  RECT 339.720 6.340 339.920 6.540 ;
  LAYER VI3 ;
  RECT 339.720 5.940 339.920 6.140 ;
  LAYER VI3 ;
  RECT 339.320 6.340 339.520 6.540 ;
  LAYER VI3 ;
  RECT 339.320 5.940 339.520 6.140 ;
  LAYER VI3 ;
  RECT 338.920 6.340 339.120 6.540 ;
  LAYER VI3 ;
  RECT 338.920 5.940 339.120 6.140 ;
  LAYER VI3 ;
  RECT 338.520 6.340 338.720 6.540 ;
  LAYER VI3 ;
  RECT 338.520 5.940 338.720 6.140 ;
  LAYER VI3 ;
  RECT 338.120 6.340 338.320 6.540 ;
  LAYER VI3 ;
  RECT 338.120 5.940 338.320 6.140 ;
  LAYER VI3 ;
  RECT 337.720 6.340 337.920 6.540 ;
  LAYER VI3 ;
  RECT 337.720 5.940 337.920 6.140 ;
  LAYER VI3 ;
  RECT 337.320 6.340 337.520 6.540 ;
  LAYER VI3 ;
  RECT 337.320 5.940 337.520 6.140 ;
  LAYER VI3 ;
  RECT 336.920 6.340 337.120 6.540 ;
  LAYER VI3 ;
  RECT 336.920 5.940 337.120 6.140 ;
  LAYER VI3 ;
  RECT 336.520 6.340 336.720 6.540 ;
  LAYER VI3 ;
  RECT 336.520 5.940 336.720 6.140 ;
  LAYER VI3 ;
  RECT 336.120 6.340 336.320 6.540 ;
  LAYER VI3 ;
  RECT 336.120 5.940 336.320 6.140 ;
  LAYER VI3 ;
  RECT 335.720 6.340 335.920 6.540 ;
  LAYER VI3 ;
  RECT 335.720 5.940 335.920 6.140 ;
  LAYER VI3 ;
  RECT 355.560 5.880 363.560 6.740 ;
  LAYER VI3 ;
  RECT 363.160 6.340 363.360 6.540 ;
  LAYER VI3 ;
  RECT 363.160 5.940 363.360 6.140 ;
  LAYER VI3 ;
  RECT 362.760 6.340 362.960 6.540 ;
  LAYER VI3 ;
  RECT 362.760 5.940 362.960 6.140 ;
  LAYER VI3 ;
  RECT 362.360 6.340 362.560 6.540 ;
  LAYER VI3 ;
  RECT 362.360 5.940 362.560 6.140 ;
  LAYER VI3 ;
  RECT 361.960 6.340 362.160 6.540 ;
  LAYER VI3 ;
  RECT 361.960 5.940 362.160 6.140 ;
  LAYER VI3 ;
  RECT 361.560 6.340 361.760 6.540 ;
  LAYER VI3 ;
  RECT 361.560 5.940 361.760 6.140 ;
  LAYER VI3 ;
  RECT 361.160 6.340 361.360 6.540 ;
  LAYER VI3 ;
  RECT 361.160 5.940 361.360 6.140 ;
  LAYER VI3 ;
  RECT 360.760 6.340 360.960 6.540 ;
  LAYER VI3 ;
  RECT 360.760 5.940 360.960 6.140 ;
  LAYER VI3 ;
  RECT 360.360 6.340 360.560 6.540 ;
  LAYER VI3 ;
  RECT 360.360 5.940 360.560 6.140 ;
  LAYER VI3 ;
  RECT 359.960 6.340 360.160 6.540 ;
  LAYER VI3 ;
  RECT 359.960 5.940 360.160 6.140 ;
  LAYER VI3 ;
  RECT 359.560 6.340 359.760 6.540 ;
  LAYER VI3 ;
  RECT 359.560 5.940 359.760 6.140 ;
  LAYER VI3 ;
  RECT 359.160 6.340 359.360 6.540 ;
  LAYER VI3 ;
  RECT 359.160 5.940 359.360 6.140 ;
  LAYER VI3 ;
  RECT 358.760 6.340 358.960 6.540 ;
  LAYER VI3 ;
  RECT 358.760 5.940 358.960 6.140 ;
  LAYER VI3 ;
  RECT 358.360 6.340 358.560 6.540 ;
  LAYER VI3 ;
  RECT 358.360 5.940 358.560 6.140 ;
  LAYER VI3 ;
  RECT 357.960 6.340 358.160 6.540 ;
  LAYER VI3 ;
  RECT 357.960 5.940 358.160 6.140 ;
  LAYER VI3 ;
  RECT 357.560 6.340 357.760 6.540 ;
  LAYER VI3 ;
  RECT 357.560 5.940 357.760 6.140 ;
  LAYER VI3 ;
  RECT 357.160 6.340 357.360 6.540 ;
  LAYER VI3 ;
  RECT 357.160 5.940 357.360 6.140 ;
  LAYER VI3 ;
  RECT 356.760 6.340 356.960 6.540 ;
  LAYER VI3 ;
  RECT 356.760 5.940 356.960 6.140 ;
  LAYER VI3 ;
  RECT 356.360 6.340 356.560 6.540 ;
  LAYER VI3 ;
  RECT 356.360 5.940 356.560 6.140 ;
  LAYER VI3 ;
  RECT 355.960 6.340 356.160 6.540 ;
  LAYER VI3 ;
  RECT 355.960 5.940 356.160 6.140 ;
  LAYER VI3 ;
  RECT 355.560 6.340 355.760 6.540 ;
  LAYER VI3 ;
  RECT 355.560 5.940 355.760 6.140 ;
  LAYER VI3 ;
  RECT 376.640 5.880 384.640 6.740 ;
  LAYER VI3 ;
  RECT 384.240 6.340 384.440 6.540 ;
  LAYER VI3 ;
  RECT 384.240 5.940 384.440 6.140 ;
  LAYER VI3 ;
  RECT 383.840 6.340 384.040 6.540 ;
  LAYER VI3 ;
  RECT 383.840 5.940 384.040 6.140 ;
  LAYER VI3 ;
  RECT 383.440 6.340 383.640 6.540 ;
  LAYER VI3 ;
  RECT 383.440 5.940 383.640 6.140 ;
  LAYER VI3 ;
  RECT 383.040 6.340 383.240 6.540 ;
  LAYER VI3 ;
  RECT 383.040 5.940 383.240 6.140 ;
  LAYER VI3 ;
  RECT 382.640 6.340 382.840 6.540 ;
  LAYER VI3 ;
  RECT 382.640 5.940 382.840 6.140 ;
  LAYER VI3 ;
  RECT 382.240 6.340 382.440 6.540 ;
  LAYER VI3 ;
  RECT 382.240 5.940 382.440 6.140 ;
  LAYER VI3 ;
  RECT 381.840 6.340 382.040 6.540 ;
  LAYER VI3 ;
  RECT 381.840 5.940 382.040 6.140 ;
  LAYER VI3 ;
  RECT 381.440 6.340 381.640 6.540 ;
  LAYER VI3 ;
  RECT 381.440 5.940 381.640 6.140 ;
  LAYER VI3 ;
  RECT 381.040 6.340 381.240 6.540 ;
  LAYER VI3 ;
  RECT 381.040 5.940 381.240 6.140 ;
  LAYER VI3 ;
  RECT 380.640 6.340 380.840 6.540 ;
  LAYER VI3 ;
  RECT 380.640 5.940 380.840 6.140 ;
  LAYER VI3 ;
  RECT 380.240 6.340 380.440 6.540 ;
  LAYER VI3 ;
  RECT 380.240 5.940 380.440 6.140 ;
  LAYER VI3 ;
  RECT 379.840 6.340 380.040 6.540 ;
  LAYER VI3 ;
  RECT 379.840 5.940 380.040 6.140 ;
  LAYER VI3 ;
  RECT 379.440 6.340 379.640 6.540 ;
  LAYER VI3 ;
  RECT 379.440 5.940 379.640 6.140 ;
  LAYER VI3 ;
  RECT 379.040 6.340 379.240 6.540 ;
  LAYER VI3 ;
  RECT 379.040 5.940 379.240 6.140 ;
  LAYER VI3 ;
  RECT 378.640 6.340 378.840 6.540 ;
  LAYER VI3 ;
  RECT 378.640 5.940 378.840 6.140 ;
  LAYER VI3 ;
  RECT 378.240 6.340 378.440 6.540 ;
  LAYER VI3 ;
  RECT 378.240 5.940 378.440 6.140 ;
  LAYER VI3 ;
  RECT 377.840 6.340 378.040 6.540 ;
  LAYER VI3 ;
  RECT 377.840 5.940 378.040 6.140 ;
  LAYER VI3 ;
  RECT 377.440 6.340 377.640 6.540 ;
  LAYER VI3 ;
  RECT 377.440 5.940 377.640 6.140 ;
  LAYER VI3 ;
  RECT 377.040 6.340 377.240 6.540 ;
  LAYER VI3 ;
  RECT 377.040 5.940 377.240 6.140 ;
  LAYER VI3 ;
  RECT 376.640 6.340 376.840 6.540 ;
  LAYER VI3 ;
  RECT 376.640 5.940 376.840 6.140 ;
  LAYER VI3 ;
  RECT 396.480 5.880 404.480 6.740 ;
  LAYER VI3 ;
  RECT 404.080 6.340 404.280 6.540 ;
  LAYER VI3 ;
  RECT 404.080 5.940 404.280 6.140 ;
  LAYER VI3 ;
  RECT 403.680 6.340 403.880 6.540 ;
  LAYER VI3 ;
  RECT 403.680 5.940 403.880 6.140 ;
  LAYER VI3 ;
  RECT 403.280 6.340 403.480 6.540 ;
  LAYER VI3 ;
  RECT 403.280 5.940 403.480 6.140 ;
  LAYER VI3 ;
  RECT 402.880 6.340 403.080 6.540 ;
  LAYER VI3 ;
  RECT 402.880 5.940 403.080 6.140 ;
  LAYER VI3 ;
  RECT 402.480 6.340 402.680 6.540 ;
  LAYER VI3 ;
  RECT 402.480 5.940 402.680 6.140 ;
  LAYER VI3 ;
  RECT 402.080 6.340 402.280 6.540 ;
  LAYER VI3 ;
  RECT 402.080 5.940 402.280 6.140 ;
  LAYER VI3 ;
  RECT 401.680 6.340 401.880 6.540 ;
  LAYER VI3 ;
  RECT 401.680 5.940 401.880 6.140 ;
  LAYER VI3 ;
  RECT 401.280 6.340 401.480 6.540 ;
  LAYER VI3 ;
  RECT 401.280 5.940 401.480 6.140 ;
  LAYER VI3 ;
  RECT 400.880 6.340 401.080 6.540 ;
  LAYER VI3 ;
  RECT 400.880 5.940 401.080 6.140 ;
  LAYER VI3 ;
  RECT 400.480 6.340 400.680 6.540 ;
  LAYER VI3 ;
  RECT 400.480 5.940 400.680 6.140 ;
  LAYER VI3 ;
  RECT 400.080 6.340 400.280 6.540 ;
  LAYER VI3 ;
  RECT 400.080 5.940 400.280 6.140 ;
  LAYER VI3 ;
  RECT 399.680 6.340 399.880 6.540 ;
  LAYER VI3 ;
  RECT 399.680 5.940 399.880 6.140 ;
  LAYER VI3 ;
  RECT 399.280 6.340 399.480 6.540 ;
  LAYER VI3 ;
  RECT 399.280 5.940 399.480 6.140 ;
  LAYER VI3 ;
  RECT 398.880 6.340 399.080 6.540 ;
  LAYER VI3 ;
  RECT 398.880 5.940 399.080 6.140 ;
  LAYER VI3 ;
  RECT 398.480 6.340 398.680 6.540 ;
  LAYER VI3 ;
  RECT 398.480 5.940 398.680 6.140 ;
  LAYER VI3 ;
  RECT 398.080 6.340 398.280 6.540 ;
  LAYER VI3 ;
  RECT 398.080 5.940 398.280 6.140 ;
  LAYER VI3 ;
  RECT 397.680 6.340 397.880 6.540 ;
  LAYER VI3 ;
  RECT 397.680 5.940 397.880 6.140 ;
  LAYER VI3 ;
  RECT 397.280 6.340 397.480 6.540 ;
  LAYER VI3 ;
  RECT 397.280 5.940 397.480 6.140 ;
  LAYER VI3 ;
  RECT 396.880 6.340 397.080 6.540 ;
  LAYER VI3 ;
  RECT 396.880 5.940 397.080 6.140 ;
  LAYER VI3 ;
  RECT 396.480 6.340 396.680 6.540 ;
  LAYER VI3 ;
  RECT 396.480 5.940 396.680 6.140 ;
  LAYER VI3 ;
  RECT 417.560 5.880 425.560 6.740 ;
  LAYER VI3 ;
  RECT 425.160 6.340 425.360 6.540 ;
  LAYER VI3 ;
  RECT 425.160 5.940 425.360 6.140 ;
  LAYER VI3 ;
  RECT 424.760 6.340 424.960 6.540 ;
  LAYER VI3 ;
  RECT 424.760 5.940 424.960 6.140 ;
  LAYER VI3 ;
  RECT 424.360 6.340 424.560 6.540 ;
  LAYER VI3 ;
  RECT 424.360 5.940 424.560 6.140 ;
  LAYER VI3 ;
  RECT 423.960 6.340 424.160 6.540 ;
  LAYER VI3 ;
  RECT 423.960 5.940 424.160 6.140 ;
  LAYER VI3 ;
  RECT 423.560 6.340 423.760 6.540 ;
  LAYER VI3 ;
  RECT 423.560 5.940 423.760 6.140 ;
  LAYER VI3 ;
  RECT 423.160 6.340 423.360 6.540 ;
  LAYER VI3 ;
  RECT 423.160 5.940 423.360 6.140 ;
  LAYER VI3 ;
  RECT 422.760 6.340 422.960 6.540 ;
  LAYER VI3 ;
  RECT 422.760 5.940 422.960 6.140 ;
  LAYER VI3 ;
  RECT 422.360 6.340 422.560 6.540 ;
  LAYER VI3 ;
  RECT 422.360 5.940 422.560 6.140 ;
  LAYER VI3 ;
  RECT 421.960 6.340 422.160 6.540 ;
  LAYER VI3 ;
  RECT 421.960 5.940 422.160 6.140 ;
  LAYER VI3 ;
  RECT 421.560 6.340 421.760 6.540 ;
  LAYER VI3 ;
  RECT 421.560 5.940 421.760 6.140 ;
  LAYER VI3 ;
  RECT 421.160 6.340 421.360 6.540 ;
  LAYER VI3 ;
  RECT 421.160 5.940 421.360 6.140 ;
  LAYER VI3 ;
  RECT 420.760 6.340 420.960 6.540 ;
  LAYER VI3 ;
  RECT 420.760 5.940 420.960 6.140 ;
  LAYER VI3 ;
  RECT 420.360 6.340 420.560 6.540 ;
  LAYER VI3 ;
  RECT 420.360 5.940 420.560 6.140 ;
  LAYER VI3 ;
  RECT 419.960 6.340 420.160 6.540 ;
  LAYER VI3 ;
  RECT 419.960 5.940 420.160 6.140 ;
  LAYER VI3 ;
  RECT 419.560 6.340 419.760 6.540 ;
  LAYER VI3 ;
  RECT 419.560 5.940 419.760 6.140 ;
  LAYER VI3 ;
  RECT 419.160 6.340 419.360 6.540 ;
  LAYER VI3 ;
  RECT 419.160 5.940 419.360 6.140 ;
  LAYER VI3 ;
  RECT 418.760 6.340 418.960 6.540 ;
  LAYER VI3 ;
  RECT 418.760 5.940 418.960 6.140 ;
  LAYER VI3 ;
  RECT 418.360 6.340 418.560 6.540 ;
  LAYER VI3 ;
  RECT 418.360 5.940 418.560 6.140 ;
  LAYER VI3 ;
  RECT 417.960 6.340 418.160 6.540 ;
  LAYER VI3 ;
  RECT 417.960 5.940 418.160 6.140 ;
  LAYER VI3 ;
  RECT 417.560 6.340 417.760 6.540 ;
  LAYER VI3 ;
  RECT 417.560 5.940 417.760 6.140 ;
  LAYER VI3 ;
  RECT 437.400 5.880 445.400 6.740 ;
  LAYER VI3 ;
  RECT 445.000 6.340 445.200 6.540 ;
  LAYER VI3 ;
  RECT 445.000 5.940 445.200 6.140 ;
  LAYER VI3 ;
  RECT 444.600 6.340 444.800 6.540 ;
  LAYER VI3 ;
  RECT 444.600 5.940 444.800 6.140 ;
  LAYER VI3 ;
  RECT 444.200 6.340 444.400 6.540 ;
  LAYER VI3 ;
  RECT 444.200 5.940 444.400 6.140 ;
  LAYER VI3 ;
  RECT 443.800 6.340 444.000 6.540 ;
  LAYER VI3 ;
  RECT 443.800 5.940 444.000 6.140 ;
  LAYER VI3 ;
  RECT 443.400 6.340 443.600 6.540 ;
  LAYER VI3 ;
  RECT 443.400 5.940 443.600 6.140 ;
  LAYER VI3 ;
  RECT 443.000 6.340 443.200 6.540 ;
  LAYER VI3 ;
  RECT 443.000 5.940 443.200 6.140 ;
  LAYER VI3 ;
  RECT 442.600 6.340 442.800 6.540 ;
  LAYER VI3 ;
  RECT 442.600 5.940 442.800 6.140 ;
  LAYER VI3 ;
  RECT 442.200 6.340 442.400 6.540 ;
  LAYER VI3 ;
  RECT 442.200 5.940 442.400 6.140 ;
  LAYER VI3 ;
  RECT 441.800 6.340 442.000 6.540 ;
  LAYER VI3 ;
  RECT 441.800 5.940 442.000 6.140 ;
  LAYER VI3 ;
  RECT 441.400 6.340 441.600 6.540 ;
  LAYER VI3 ;
  RECT 441.400 5.940 441.600 6.140 ;
  LAYER VI3 ;
  RECT 441.000 6.340 441.200 6.540 ;
  LAYER VI3 ;
  RECT 441.000 5.940 441.200 6.140 ;
  LAYER VI3 ;
  RECT 440.600 6.340 440.800 6.540 ;
  LAYER VI3 ;
  RECT 440.600 5.940 440.800 6.140 ;
  LAYER VI3 ;
  RECT 440.200 6.340 440.400 6.540 ;
  LAYER VI3 ;
  RECT 440.200 5.940 440.400 6.140 ;
  LAYER VI3 ;
  RECT 439.800 6.340 440.000 6.540 ;
  LAYER VI3 ;
  RECT 439.800 5.940 440.000 6.140 ;
  LAYER VI3 ;
  RECT 439.400 6.340 439.600 6.540 ;
  LAYER VI3 ;
  RECT 439.400 5.940 439.600 6.140 ;
  LAYER VI3 ;
  RECT 439.000 6.340 439.200 6.540 ;
  LAYER VI3 ;
  RECT 439.000 5.940 439.200 6.140 ;
  LAYER VI3 ;
  RECT 438.600 6.340 438.800 6.540 ;
  LAYER VI3 ;
  RECT 438.600 5.940 438.800 6.140 ;
  LAYER VI3 ;
  RECT 438.200 6.340 438.400 6.540 ;
  LAYER VI3 ;
  RECT 438.200 5.940 438.400 6.140 ;
  LAYER VI3 ;
  RECT 437.800 6.340 438.000 6.540 ;
  LAYER VI3 ;
  RECT 437.800 5.940 438.000 6.140 ;
  LAYER VI3 ;
  RECT 437.400 6.340 437.600 6.540 ;
  LAYER VI3 ;
  RECT 437.400 5.940 437.600 6.140 ;
  LAYER VI3 ;
  RECT 458.480 5.880 466.480 6.740 ;
  LAYER VI3 ;
  RECT 466.080 6.340 466.280 6.540 ;
  LAYER VI3 ;
  RECT 466.080 5.940 466.280 6.140 ;
  LAYER VI3 ;
  RECT 465.680 6.340 465.880 6.540 ;
  LAYER VI3 ;
  RECT 465.680 5.940 465.880 6.140 ;
  LAYER VI3 ;
  RECT 465.280 6.340 465.480 6.540 ;
  LAYER VI3 ;
  RECT 465.280 5.940 465.480 6.140 ;
  LAYER VI3 ;
  RECT 464.880 6.340 465.080 6.540 ;
  LAYER VI3 ;
  RECT 464.880 5.940 465.080 6.140 ;
  LAYER VI3 ;
  RECT 464.480 6.340 464.680 6.540 ;
  LAYER VI3 ;
  RECT 464.480 5.940 464.680 6.140 ;
  LAYER VI3 ;
  RECT 464.080 6.340 464.280 6.540 ;
  LAYER VI3 ;
  RECT 464.080 5.940 464.280 6.140 ;
  LAYER VI3 ;
  RECT 463.680 6.340 463.880 6.540 ;
  LAYER VI3 ;
  RECT 463.680 5.940 463.880 6.140 ;
  LAYER VI3 ;
  RECT 463.280 6.340 463.480 6.540 ;
  LAYER VI3 ;
  RECT 463.280 5.940 463.480 6.140 ;
  LAYER VI3 ;
  RECT 462.880 6.340 463.080 6.540 ;
  LAYER VI3 ;
  RECT 462.880 5.940 463.080 6.140 ;
  LAYER VI3 ;
  RECT 462.480 6.340 462.680 6.540 ;
  LAYER VI3 ;
  RECT 462.480 5.940 462.680 6.140 ;
  LAYER VI3 ;
  RECT 462.080 6.340 462.280 6.540 ;
  LAYER VI3 ;
  RECT 462.080 5.940 462.280 6.140 ;
  LAYER VI3 ;
  RECT 461.680 6.340 461.880 6.540 ;
  LAYER VI3 ;
  RECT 461.680 5.940 461.880 6.140 ;
  LAYER VI3 ;
  RECT 461.280 6.340 461.480 6.540 ;
  LAYER VI3 ;
  RECT 461.280 5.940 461.480 6.140 ;
  LAYER VI3 ;
  RECT 460.880 6.340 461.080 6.540 ;
  LAYER VI3 ;
  RECT 460.880 5.940 461.080 6.140 ;
  LAYER VI3 ;
  RECT 460.480 6.340 460.680 6.540 ;
  LAYER VI3 ;
  RECT 460.480 5.940 460.680 6.140 ;
  LAYER VI3 ;
  RECT 460.080 6.340 460.280 6.540 ;
  LAYER VI3 ;
  RECT 460.080 5.940 460.280 6.140 ;
  LAYER VI3 ;
  RECT 459.680 6.340 459.880 6.540 ;
  LAYER VI3 ;
  RECT 459.680 5.940 459.880 6.140 ;
  LAYER VI3 ;
  RECT 459.280 6.340 459.480 6.540 ;
  LAYER VI3 ;
  RECT 459.280 5.940 459.480 6.140 ;
  LAYER VI3 ;
  RECT 458.880 6.340 459.080 6.540 ;
  LAYER VI3 ;
  RECT 458.880 5.940 459.080 6.140 ;
  LAYER VI3 ;
  RECT 458.480 6.340 458.680 6.540 ;
  LAYER VI3 ;
  RECT 458.480 5.940 458.680 6.140 ;
  LAYER VI3 ;
  RECT 478.320 5.880 486.320 6.740 ;
  LAYER VI3 ;
  RECT 485.920 6.340 486.120 6.540 ;
  LAYER VI3 ;
  RECT 485.920 5.940 486.120 6.140 ;
  LAYER VI3 ;
  RECT 485.520 6.340 485.720 6.540 ;
  LAYER VI3 ;
  RECT 485.520 5.940 485.720 6.140 ;
  LAYER VI3 ;
  RECT 485.120 6.340 485.320 6.540 ;
  LAYER VI3 ;
  RECT 485.120 5.940 485.320 6.140 ;
  LAYER VI3 ;
  RECT 484.720 6.340 484.920 6.540 ;
  LAYER VI3 ;
  RECT 484.720 5.940 484.920 6.140 ;
  LAYER VI3 ;
  RECT 484.320 6.340 484.520 6.540 ;
  LAYER VI3 ;
  RECT 484.320 5.940 484.520 6.140 ;
  LAYER VI3 ;
  RECT 483.920 6.340 484.120 6.540 ;
  LAYER VI3 ;
  RECT 483.920 5.940 484.120 6.140 ;
  LAYER VI3 ;
  RECT 483.520 6.340 483.720 6.540 ;
  LAYER VI3 ;
  RECT 483.520 5.940 483.720 6.140 ;
  LAYER VI3 ;
  RECT 483.120 6.340 483.320 6.540 ;
  LAYER VI3 ;
  RECT 483.120 5.940 483.320 6.140 ;
  LAYER VI3 ;
  RECT 482.720 6.340 482.920 6.540 ;
  LAYER VI3 ;
  RECT 482.720 5.940 482.920 6.140 ;
  LAYER VI3 ;
  RECT 482.320 6.340 482.520 6.540 ;
  LAYER VI3 ;
  RECT 482.320 5.940 482.520 6.140 ;
  LAYER VI3 ;
  RECT 481.920 6.340 482.120 6.540 ;
  LAYER VI3 ;
  RECT 481.920 5.940 482.120 6.140 ;
  LAYER VI3 ;
  RECT 481.520 6.340 481.720 6.540 ;
  LAYER VI3 ;
  RECT 481.520 5.940 481.720 6.140 ;
  LAYER VI3 ;
  RECT 481.120 6.340 481.320 6.540 ;
  LAYER VI3 ;
  RECT 481.120 5.940 481.320 6.140 ;
  LAYER VI3 ;
  RECT 480.720 6.340 480.920 6.540 ;
  LAYER VI3 ;
  RECT 480.720 5.940 480.920 6.140 ;
  LAYER VI3 ;
  RECT 480.320 6.340 480.520 6.540 ;
  LAYER VI3 ;
  RECT 480.320 5.940 480.520 6.140 ;
  LAYER VI3 ;
  RECT 479.920 6.340 480.120 6.540 ;
  LAYER VI3 ;
  RECT 479.920 5.940 480.120 6.140 ;
  LAYER VI3 ;
  RECT 479.520 6.340 479.720 6.540 ;
  LAYER VI3 ;
  RECT 479.520 5.940 479.720 6.140 ;
  LAYER VI3 ;
  RECT 479.120 6.340 479.320 6.540 ;
  LAYER VI3 ;
  RECT 479.120 5.940 479.320 6.140 ;
  LAYER VI3 ;
  RECT 478.720 6.340 478.920 6.540 ;
  LAYER VI3 ;
  RECT 478.720 5.940 478.920 6.140 ;
  LAYER VI3 ;
  RECT 478.320 6.340 478.520 6.540 ;
  LAYER VI3 ;
  RECT 478.320 5.940 478.520 6.140 ;
  LAYER VI3 ;
  RECT 499.400 5.880 507.400 6.740 ;
  LAYER VI3 ;
  RECT 507.000 6.340 507.200 6.540 ;
  LAYER VI3 ;
  RECT 507.000 5.940 507.200 6.140 ;
  LAYER VI3 ;
  RECT 506.600 6.340 506.800 6.540 ;
  LAYER VI3 ;
  RECT 506.600 5.940 506.800 6.140 ;
  LAYER VI3 ;
  RECT 506.200 6.340 506.400 6.540 ;
  LAYER VI3 ;
  RECT 506.200 5.940 506.400 6.140 ;
  LAYER VI3 ;
  RECT 505.800 6.340 506.000 6.540 ;
  LAYER VI3 ;
  RECT 505.800 5.940 506.000 6.140 ;
  LAYER VI3 ;
  RECT 505.400 6.340 505.600 6.540 ;
  LAYER VI3 ;
  RECT 505.400 5.940 505.600 6.140 ;
  LAYER VI3 ;
  RECT 505.000 6.340 505.200 6.540 ;
  LAYER VI3 ;
  RECT 505.000 5.940 505.200 6.140 ;
  LAYER VI3 ;
  RECT 504.600 6.340 504.800 6.540 ;
  LAYER VI3 ;
  RECT 504.600 5.940 504.800 6.140 ;
  LAYER VI3 ;
  RECT 504.200 6.340 504.400 6.540 ;
  LAYER VI3 ;
  RECT 504.200 5.940 504.400 6.140 ;
  LAYER VI3 ;
  RECT 503.800 6.340 504.000 6.540 ;
  LAYER VI3 ;
  RECT 503.800 5.940 504.000 6.140 ;
  LAYER VI3 ;
  RECT 503.400 6.340 503.600 6.540 ;
  LAYER VI3 ;
  RECT 503.400 5.940 503.600 6.140 ;
  LAYER VI3 ;
  RECT 503.000 6.340 503.200 6.540 ;
  LAYER VI3 ;
  RECT 503.000 5.940 503.200 6.140 ;
  LAYER VI3 ;
  RECT 502.600 6.340 502.800 6.540 ;
  LAYER VI3 ;
  RECT 502.600 5.940 502.800 6.140 ;
  LAYER VI3 ;
  RECT 502.200 6.340 502.400 6.540 ;
  LAYER VI3 ;
  RECT 502.200 5.940 502.400 6.140 ;
  LAYER VI3 ;
  RECT 501.800 6.340 502.000 6.540 ;
  LAYER VI3 ;
  RECT 501.800 5.940 502.000 6.140 ;
  LAYER VI3 ;
  RECT 501.400 6.340 501.600 6.540 ;
  LAYER VI3 ;
  RECT 501.400 5.940 501.600 6.140 ;
  LAYER VI3 ;
  RECT 501.000 6.340 501.200 6.540 ;
  LAYER VI3 ;
  RECT 501.000 5.940 501.200 6.140 ;
  LAYER VI3 ;
  RECT 500.600 6.340 500.800 6.540 ;
  LAYER VI3 ;
  RECT 500.600 5.940 500.800 6.140 ;
  LAYER VI3 ;
  RECT 500.200 6.340 500.400 6.540 ;
  LAYER VI3 ;
  RECT 500.200 5.940 500.400 6.140 ;
  LAYER VI3 ;
  RECT 499.800 6.340 500.000 6.540 ;
  LAYER VI3 ;
  RECT 499.800 5.940 500.000 6.140 ;
  LAYER VI3 ;
  RECT 499.400 6.340 499.600 6.540 ;
  LAYER VI3 ;
  RECT 499.400 5.940 499.600 6.140 ;
  LAYER VI3 ;
  RECT 519.240 5.880 527.240 6.740 ;
  LAYER VI3 ;
  RECT 526.840 6.340 527.040 6.540 ;
  LAYER VI3 ;
  RECT 526.840 5.940 527.040 6.140 ;
  LAYER VI3 ;
  RECT 526.440 6.340 526.640 6.540 ;
  LAYER VI3 ;
  RECT 526.440 5.940 526.640 6.140 ;
  LAYER VI3 ;
  RECT 526.040 6.340 526.240 6.540 ;
  LAYER VI3 ;
  RECT 526.040 5.940 526.240 6.140 ;
  LAYER VI3 ;
  RECT 525.640 6.340 525.840 6.540 ;
  LAYER VI3 ;
  RECT 525.640 5.940 525.840 6.140 ;
  LAYER VI3 ;
  RECT 525.240 6.340 525.440 6.540 ;
  LAYER VI3 ;
  RECT 525.240 5.940 525.440 6.140 ;
  LAYER VI3 ;
  RECT 524.840 6.340 525.040 6.540 ;
  LAYER VI3 ;
  RECT 524.840 5.940 525.040 6.140 ;
  LAYER VI3 ;
  RECT 524.440 6.340 524.640 6.540 ;
  LAYER VI3 ;
  RECT 524.440 5.940 524.640 6.140 ;
  LAYER VI3 ;
  RECT 524.040 6.340 524.240 6.540 ;
  LAYER VI3 ;
  RECT 524.040 5.940 524.240 6.140 ;
  LAYER VI3 ;
  RECT 523.640 6.340 523.840 6.540 ;
  LAYER VI3 ;
  RECT 523.640 5.940 523.840 6.140 ;
  LAYER VI3 ;
  RECT 523.240 6.340 523.440 6.540 ;
  LAYER VI3 ;
  RECT 523.240 5.940 523.440 6.140 ;
  LAYER VI3 ;
  RECT 522.840 6.340 523.040 6.540 ;
  LAYER VI3 ;
  RECT 522.840 5.940 523.040 6.140 ;
  LAYER VI3 ;
  RECT 522.440 6.340 522.640 6.540 ;
  LAYER VI3 ;
  RECT 522.440 5.940 522.640 6.140 ;
  LAYER VI3 ;
  RECT 522.040 6.340 522.240 6.540 ;
  LAYER VI3 ;
  RECT 522.040 5.940 522.240 6.140 ;
  LAYER VI3 ;
  RECT 521.640 6.340 521.840 6.540 ;
  LAYER VI3 ;
  RECT 521.640 5.940 521.840 6.140 ;
  LAYER VI3 ;
  RECT 521.240 6.340 521.440 6.540 ;
  LAYER VI3 ;
  RECT 521.240 5.940 521.440 6.140 ;
  LAYER VI3 ;
  RECT 520.840 6.340 521.040 6.540 ;
  LAYER VI3 ;
  RECT 520.840 5.940 521.040 6.140 ;
  LAYER VI3 ;
  RECT 520.440 6.340 520.640 6.540 ;
  LAYER VI3 ;
  RECT 520.440 5.940 520.640 6.140 ;
  LAYER VI3 ;
  RECT 520.040 6.340 520.240 6.540 ;
  LAYER VI3 ;
  RECT 520.040 5.940 520.240 6.140 ;
  LAYER VI3 ;
  RECT 519.640 6.340 519.840 6.540 ;
  LAYER VI3 ;
  RECT 519.640 5.940 519.840 6.140 ;
  LAYER VI3 ;
  RECT 519.240 6.340 519.440 6.540 ;
  LAYER VI3 ;
  RECT 519.240 5.940 519.440 6.140 ;
  LAYER VI3 ;
  RECT 540.320 5.880 548.320 6.740 ;
  LAYER VI3 ;
  RECT 547.920 6.340 548.120 6.540 ;
  LAYER VI3 ;
  RECT 547.920 5.940 548.120 6.140 ;
  LAYER VI3 ;
  RECT 547.520 6.340 547.720 6.540 ;
  LAYER VI3 ;
  RECT 547.520 5.940 547.720 6.140 ;
  LAYER VI3 ;
  RECT 547.120 6.340 547.320 6.540 ;
  LAYER VI3 ;
  RECT 547.120 5.940 547.320 6.140 ;
  LAYER VI3 ;
  RECT 546.720 6.340 546.920 6.540 ;
  LAYER VI3 ;
  RECT 546.720 5.940 546.920 6.140 ;
  LAYER VI3 ;
  RECT 546.320 6.340 546.520 6.540 ;
  LAYER VI3 ;
  RECT 546.320 5.940 546.520 6.140 ;
  LAYER VI3 ;
  RECT 545.920 6.340 546.120 6.540 ;
  LAYER VI3 ;
  RECT 545.920 5.940 546.120 6.140 ;
  LAYER VI3 ;
  RECT 545.520 6.340 545.720 6.540 ;
  LAYER VI3 ;
  RECT 545.520 5.940 545.720 6.140 ;
  LAYER VI3 ;
  RECT 545.120 6.340 545.320 6.540 ;
  LAYER VI3 ;
  RECT 545.120 5.940 545.320 6.140 ;
  LAYER VI3 ;
  RECT 544.720 6.340 544.920 6.540 ;
  LAYER VI3 ;
  RECT 544.720 5.940 544.920 6.140 ;
  LAYER VI3 ;
  RECT 544.320 6.340 544.520 6.540 ;
  LAYER VI3 ;
  RECT 544.320 5.940 544.520 6.140 ;
  LAYER VI3 ;
  RECT 543.920 6.340 544.120 6.540 ;
  LAYER VI3 ;
  RECT 543.920 5.940 544.120 6.140 ;
  LAYER VI3 ;
  RECT 543.520 6.340 543.720 6.540 ;
  LAYER VI3 ;
  RECT 543.520 5.940 543.720 6.140 ;
  LAYER VI3 ;
  RECT 543.120 6.340 543.320 6.540 ;
  LAYER VI3 ;
  RECT 543.120 5.940 543.320 6.140 ;
  LAYER VI3 ;
  RECT 542.720 6.340 542.920 6.540 ;
  LAYER VI3 ;
  RECT 542.720 5.940 542.920 6.140 ;
  LAYER VI3 ;
  RECT 542.320 6.340 542.520 6.540 ;
  LAYER VI3 ;
  RECT 542.320 5.940 542.520 6.140 ;
  LAYER VI3 ;
  RECT 541.920 6.340 542.120 6.540 ;
  LAYER VI3 ;
  RECT 541.920 5.940 542.120 6.140 ;
  LAYER VI3 ;
  RECT 541.520 6.340 541.720 6.540 ;
  LAYER VI3 ;
  RECT 541.520 5.940 541.720 6.140 ;
  LAYER VI3 ;
  RECT 541.120 6.340 541.320 6.540 ;
  LAYER VI3 ;
  RECT 541.120 5.940 541.320 6.140 ;
  LAYER VI3 ;
  RECT 540.720 6.340 540.920 6.540 ;
  LAYER VI3 ;
  RECT 540.720 5.940 540.920 6.140 ;
  LAYER VI3 ;
  RECT 540.320 6.340 540.520 6.540 ;
  LAYER VI3 ;
  RECT 540.320 5.940 540.520 6.140 ;
  LAYER VI3 ;
  RECT 560.160 5.880 568.160 6.740 ;
  LAYER VI3 ;
  RECT 567.760 6.340 567.960 6.540 ;
  LAYER VI3 ;
  RECT 567.760 5.940 567.960 6.140 ;
  LAYER VI3 ;
  RECT 567.360 6.340 567.560 6.540 ;
  LAYER VI3 ;
  RECT 567.360 5.940 567.560 6.140 ;
  LAYER VI3 ;
  RECT 566.960 6.340 567.160 6.540 ;
  LAYER VI3 ;
  RECT 566.960 5.940 567.160 6.140 ;
  LAYER VI3 ;
  RECT 566.560 6.340 566.760 6.540 ;
  LAYER VI3 ;
  RECT 566.560 5.940 566.760 6.140 ;
  LAYER VI3 ;
  RECT 566.160 6.340 566.360 6.540 ;
  LAYER VI3 ;
  RECT 566.160 5.940 566.360 6.140 ;
  LAYER VI3 ;
  RECT 565.760 6.340 565.960 6.540 ;
  LAYER VI3 ;
  RECT 565.760 5.940 565.960 6.140 ;
  LAYER VI3 ;
  RECT 565.360 6.340 565.560 6.540 ;
  LAYER VI3 ;
  RECT 565.360 5.940 565.560 6.140 ;
  LAYER VI3 ;
  RECT 564.960 6.340 565.160 6.540 ;
  LAYER VI3 ;
  RECT 564.960 5.940 565.160 6.140 ;
  LAYER VI3 ;
  RECT 564.560 6.340 564.760 6.540 ;
  LAYER VI3 ;
  RECT 564.560 5.940 564.760 6.140 ;
  LAYER VI3 ;
  RECT 564.160 6.340 564.360 6.540 ;
  LAYER VI3 ;
  RECT 564.160 5.940 564.360 6.140 ;
  LAYER VI3 ;
  RECT 563.760 6.340 563.960 6.540 ;
  LAYER VI3 ;
  RECT 563.760 5.940 563.960 6.140 ;
  LAYER VI3 ;
  RECT 563.360 6.340 563.560 6.540 ;
  LAYER VI3 ;
  RECT 563.360 5.940 563.560 6.140 ;
  LAYER VI3 ;
  RECT 562.960 6.340 563.160 6.540 ;
  LAYER VI3 ;
  RECT 562.960 5.940 563.160 6.140 ;
  LAYER VI3 ;
  RECT 562.560 6.340 562.760 6.540 ;
  LAYER VI3 ;
  RECT 562.560 5.940 562.760 6.140 ;
  LAYER VI3 ;
  RECT 562.160 6.340 562.360 6.540 ;
  LAYER VI3 ;
  RECT 562.160 5.940 562.360 6.140 ;
  LAYER VI3 ;
  RECT 561.760 6.340 561.960 6.540 ;
  LAYER VI3 ;
  RECT 561.760 5.940 561.960 6.140 ;
  LAYER VI3 ;
  RECT 561.360 6.340 561.560 6.540 ;
  LAYER VI3 ;
  RECT 561.360 5.940 561.560 6.140 ;
  LAYER VI3 ;
  RECT 560.960 6.340 561.160 6.540 ;
  LAYER VI3 ;
  RECT 560.960 5.940 561.160 6.140 ;
  LAYER VI3 ;
  RECT 560.560 6.340 560.760 6.540 ;
  LAYER VI3 ;
  RECT 560.560 5.940 560.760 6.140 ;
  LAYER VI3 ;
  RECT 560.160 6.340 560.360 6.540 ;
  LAYER VI3 ;
  RECT 560.160 5.940 560.360 6.140 ;
  LAYER VI3 ;
  RECT 581.240 5.880 589.240 6.740 ;
  LAYER VI3 ;
  RECT 588.840 6.340 589.040 6.540 ;
  LAYER VI3 ;
  RECT 588.840 5.940 589.040 6.140 ;
  LAYER VI3 ;
  RECT 588.440 6.340 588.640 6.540 ;
  LAYER VI3 ;
  RECT 588.440 5.940 588.640 6.140 ;
  LAYER VI3 ;
  RECT 588.040 6.340 588.240 6.540 ;
  LAYER VI3 ;
  RECT 588.040 5.940 588.240 6.140 ;
  LAYER VI3 ;
  RECT 587.640 6.340 587.840 6.540 ;
  LAYER VI3 ;
  RECT 587.640 5.940 587.840 6.140 ;
  LAYER VI3 ;
  RECT 587.240 6.340 587.440 6.540 ;
  LAYER VI3 ;
  RECT 587.240 5.940 587.440 6.140 ;
  LAYER VI3 ;
  RECT 586.840 6.340 587.040 6.540 ;
  LAYER VI3 ;
  RECT 586.840 5.940 587.040 6.140 ;
  LAYER VI3 ;
  RECT 586.440 6.340 586.640 6.540 ;
  LAYER VI3 ;
  RECT 586.440 5.940 586.640 6.140 ;
  LAYER VI3 ;
  RECT 586.040 6.340 586.240 6.540 ;
  LAYER VI3 ;
  RECT 586.040 5.940 586.240 6.140 ;
  LAYER VI3 ;
  RECT 585.640 6.340 585.840 6.540 ;
  LAYER VI3 ;
  RECT 585.640 5.940 585.840 6.140 ;
  LAYER VI3 ;
  RECT 585.240 6.340 585.440 6.540 ;
  LAYER VI3 ;
  RECT 585.240 5.940 585.440 6.140 ;
  LAYER VI3 ;
  RECT 584.840 6.340 585.040 6.540 ;
  LAYER VI3 ;
  RECT 584.840 5.940 585.040 6.140 ;
  LAYER VI3 ;
  RECT 584.440 6.340 584.640 6.540 ;
  LAYER VI3 ;
  RECT 584.440 5.940 584.640 6.140 ;
  LAYER VI3 ;
  RECT 584.040 6.340 584.240 6.540 ;
  LAYER VI3 ;
  RECT 584.040 5.940 584.240 6.140 ;
  LAYER VI3 ;
  RECT 583.640 6.340 583.840 6.540 ;
  LAYER VI3 ;
  RECT 583.640 5.940 583.840 6.140 ;
  LAYER VI3 ;
  RECT 583.240 6.340 583.440 6.540 ;
  LAYER VI3 ;
  RECT 583.240 5.940 583.440 6.140 ;
  LAYER VI3 ;
  RECT 582.840 6.340 583.040 6.540 ;
  LAYER VI3 ;
  RECT 582.840 5.940 583.040 6.140 ;
  LAYER VI3 ;
  RECT 582.440 6.340 582.640 6.540 ;
  LAYER VI3 ;
  RECT 582.440 5.940 582.640 6.140 ;
  LAYER VI3 ;
  RECT 582.040 6.340 582.240 6.540 ;
  LAYER VI3 ;
  RECT 582.040 5.940 582.240 6.140 ;
  LAYER VI3 ;
  RECT 581.640 6.340 581.840 6.540 ;
  LAYER VI3 ;
  RECT 581.640 5.940 581.840 6.140 ;
  LAYER VI3 ;
  RECT 581.240 6.340 581.440 6.540 ;
  LAYER VI3 ;
  RECT 581.240 5.940 581.440 6.140 ;
  LAYER VI3 ;
  RECT 601.080 5.880 609.080 6.740 ;
  LAYER VI3 ;
  RECT 608.680 6.340 608.880 6.540 ;
  LAYER VI3 ;
  RECT 608.680 5.940 608.880 6.140 ;
  LAYER VI3 ;
  RECT 608.280 6.340 608.480 6.540 ;
  LAYER VI3 ;
  RECT 608.280 5.940 608.480 6.140 ;
  LAYER VI3 ;
  RECT 607.880 6.340 608.080 6.540 ;
  LAYER VI3 ;
  RECT 607.880 5.940 608.080 6.140 ;
  LAYER VI3 ;
  RECT 607.480 6.340 607.680 6.540 ;
  LAYER VI3 ;
  RECT 607.480 5.940 607.680 6.140 ;
  LAYER VI3 ;
  RECT 607.080 6.340 607.280 6.540 ;
  LAYER VI3 ;
  RECT 607.080 5.940 607.280 6.140 ;
  LAYER VI3 ;
  RECT 606.680 6.340 606.880 6.540 ;
  LAYER VI3 ;
  RECT 606.680 5.940 606.880 6.140 ;
  LAYER VI3 ;
  RECT 606.280 6.340 606.480 6.540 ;
  LAYER VI3 ;
  RECT 606.280 5.940 606.480 6.140 ;
  LAYER VI3 ;
  RECT 605.880 6.340 606.080 6.540 ;
  LAYER VI3 ;
  RECT 605.880 5.940 606.080 6.140 ;
  LAYER VI3 ;
  RECT 605.480 6.340 605.680 6.540 ;
  LAYER VI3 ;
  RECT 605.480 5.940 605.680 6.140 ;
  LAYER VI3 ;
  RECT 605.080 6.340 605.280 6.540 ;
  LAYER VI3 ;
  RECT 605.080 5.940 605.280 6.140 ;
  LAYER VI3 ;
  RECT 604.680 6.340 604.880 6.540 ;
  LAYER VI3 ;
  RECT 604.680 5.940 604.880 6.140 ;
  LAYER VI3 ;
  RECT 604.280 6.340 604.480 6.540 ;
  LAYER VI3 ;
  RECT 604.280 5.940 604.480 6.140 ;
  LAYER VI3 ;
  RECT 603.880 6.340 604.080 6.540 ;
  LAYER VI3 ;
  RECT 603.880 5.940 604.080 6.140 ;
  LAYER VI3 ;
  RECT 603.480 6.340 603.680 6.540 ;
  LAYER VI3 ;
  RECT 603.480 5.940 603.680 6.140 ;
  LAYER VI3 ;
  RECT 603.080 6.340 603.280 6.540 ;
  LAYER VI3 ;
  RECT 603.080 5.940 603.280 6.140 ;
  LAYER VI3 ;
  RECT 602.680 6.340 602.880 6.540 ;
  LAYER VI3 ;
  RECT 602.680 5.940 602.880 6.140 ;
  LAYER VI3 ;
  RECT 602.280 6.340 602.480 6.540 ;
  LAYER VI3 ;
  RECT 602.280 5.940 602.480 6.140 ;
  LAYER VI3 ;
  RECT 601.880 6.340 602.080 6.540 ;
  LAYER VI3 ;
  RECT 601.880 5.940 602.080 6.140 ;
  LAYER VI3 ;
  RECT 601.480 6.340 601.680 6.540 ;
  LAYER VI3 ;
  RECT 601.480 5.940 601.680 6.140 ;
  LAYER VI3 ;
  RECT 601.080 6.340 601.280 6.540 ;
  LAYER VI3 ;
  RECT 601.080 5.940 601.280 6.140 ;
  LAYER VI3 ;
  RECT 622.160 5.880 630.160 6.740 ;
  LAYER VI3 ;
  RECT 629.760 6.340 629.960 6.540 ;
  LAYER VI3 ;
  RECT 629.760 5.940 629.960 6.140 ;
  LAYER VI3 ;
  RECT 629.360 6.340 629.560 6.540 ;
  LAYER VI3 ;
  RECT 629.360 5.940 629.560 6.140 ;
  LAYER VI3 ;
  RECT 628.960 6.340 629.160 6.540 ;
  LAYER VI3 ;
  RECT 628.960 5.940 629.160 6.140 ;
  LAYER VI3 ;
  RECT 628.560 6.340 628.760 6.540 ;
  LAYER VI3 ;
  RECT 628.560 5.940 628.760 6.140 ;
  LAYER VI3 ;
  RECT 628.160 6.340 628.360 6.540 ;
  LAYER VI3 ;
  RECT 628.160 5.940 628.360 6.140 ;
  LAYER VI3 ;
  RECT 627.760 6.340 627.960 6.540 ;
  LAYER VI3 ;
  RECT 627.760 5.940 627.960 6.140 ;
  LAYER VI3 ;
  RECT 627.360 6.340 627.560 6.540 ;
  LAYER VI3 ;
  RECT 627.360 5.940 627.560 6.140 ;
  LAYER VI3 ;
  RECT 626.960 6.340 627.160 6.540 ;
  LAYER VI3 ;
  RECT 626.960 5.940 627.160 6.140 ;
  LAYER VI3 ;
  RECT 626.560 6.340 626.760 6.540 ;
  LAYER VI3 ;
  RECT 626.560 5.940 626.760 6.140 ;
  LAYER VI3 ;
  RECT 626.160 6.340 626.360 6.540 ;
  LAYER VI3 ;
  RECT 626.160 5.940 626.360 6.140 ;
  LAYER VI3 ;
  RECT 625.760 6.340 625.960 6.540 ;
  LAYER VI3 ;
  RECT 625.760 5.940 625.960 6.140 ;
  LAYER VI3 ;
  RECT 625.360 6.340 625.560 6.540 ;
  LAYER VI3 ;
  RECT 625.360 5.940 625.560 6.140 ;
  LAYER VI3 ;
  RECT 624.960 6.340 625.160 6.540 ;
  LAYER VI3 ;
  RECT 624.960 5.940 625.160 6.140 ;
  LAYER VI3 ;
  RECT 624.560 6.340 624.760 6.540 ;
  LAYER VI3 ;
  RECT 624.560 5.940 624.760 6.140 ;
  LAYER VI3 ;
  RECT 624.160 6.340 624.360 6.540 ;
  LAYER VI3 ;
  RECT 624.160 5.940 624.360 6.140 ;
  LAYER VI3 ;
  RECT 623.760 6.340 623.960 6.540 ;
  LAYER VI3 ;
  RECT 623.760 5.940 623.960 6.140 ;
  LAYER VI3 ;
  RECT 623.360 6.340 623.560 6.540 ;
  LAYER VI3 ;
  RECT 623.360 5.940 623.560 6.140 ;
  LAYER VI3 ;
  RECT 622.960 6.340 623.160 6.540 ;
  LAYER VI3 ;
  RECT 622.960 5.940 623.160 6.140 ;
  LAYER VI3 ;
  RECT 622.560 6.340 622.760 6.540 ;
  LAYER VI3 ;
  RECT 622.560 5.940 622.760 6.140 ;
  LAYER VI3 ;
  RECT 622.160 6.340 622.360 6.540 ;
  LAYER VI3 ;
  RECT 622.160 5.940 622.360 6.140 ;
  LAYER VI3 ;
  RECT 642.000 5.880 650.000 6.740 ;
  LAYER VI3 ;
  RECT 649.600 6.340 649.800 6.540 ;
  LAYER VI3 ;
  RECT 649.600 5.940 649.800 6.140 ;
  LAYER VI3 ;
  RECT 649.200 6.340 649.400 6.540 ;
  LAYER VI3 ;
  RECT 649.200 5.940 649.400 6.140 ;
  LAYER VI3 ;
  RECT 648.800 6.340 649.000 6.540 ;
  LAYER VI3 ;
  RECT 648.800 5.940 649.000 6.140 ;
  LAYER VI3 ;
  RECT 648.400 6.340 648.600 6.540 ;
  LAYER VI3 ;
  RECT 648.400 5.940 648.600 6.140 ;
  LAYER VI3 ;
  RECT 648.000 6.340 648.200 6.540 ;
  LAYER VI3 ;
  RECT 648.000 5.940 648.200 6.140 ;
  LAYER VI3 ;
  RECT 647.600 6.340 647.800 6.540 ;
  LAYER VI3 ;
  RECT 647.600 5.940 647.800 6.140 ;
  LAYER VI3 ;
  RECT 647.200 6.340 647.400 6.540 ;
  LAYER VI3 ;
  RECT 647.200 5.940 647.400 6.140 ;
  LAYER VI3 ;
  RECT 646.800 6.340 647.000 6.540 ;
  LAYER VI3 ;
  RECT 646.800 5.940 647.000 6.140 ;
  LAYER VI3 ;
  RECT 646.400 6.340 646.600 6.540 ;
  LAYER VI3 ;
  RECT 646.400 5.940 646.600 6.140 ;
  LAYER VI3 ;
  RECT 646.000 6.340 646.200 6.540 ;
  LAYER VI3 ;
  RECT 646.000 5.940 646.200 6.140 ;
  LAYER VI3 ;
  RECT 645.600 6.340 645.800 6.540 ;
  LAYER VI3 ;
  RECT 645.600 5.940 645.800 6.140 ;
  LAYER VI3 ;
  RECT 645.200 6.340 645.400 6.540 ;
  LAYER VI3 ;
  RECT 645.200 5.940 645.400 6.140 ;
  LAYER VI3 ;
  RECT 644.800 6.340 645.000 6.540 ;
  LAYER VI3 ;
  RECT 644.800 5.940 645.000 6.140 ;
  LAYER VI3 ;
  RECT 644.400 6.340 644.600 6.540 ;
  LAYER VI3 ;
  RECT 644.400 5.940 644.600 6.140 ;
  LAYER VI3 ;
  RECT 644.000 6.340 644.200 6.540 ;
  LAYER VI3 ;
  RECT 644.000 5.940 644.200 6.140 ;
  LAYER VI3 ;
  RECT 643.600 6.340 643.800 6.540 ;
  LAYER VI3 ;
  RECT 643.600 5.940 643.800 6.140 ;
  LAYER VI3 ;
  RECT 643.200 6.340 643.400 6.540 ;
  LAYER VI3 ;
  RECT 643.200 5.940 643.400 6.140 ;
  LAYER VI3 ;
  RECT 642.800 6.340 643.000 6.540 ;
  LAYER VI3 ;
  RECT 642.800 5.940 643.000 6.140 ;
  LAYER VI3 ;
  RECT 642.400 6.340 642.600 6.540 ;
  LAYER VI3 ;
  RECT 642.400 5.940 642.600 6.140 ;
  LAYER VI3 ;
  RECT 642.000 6.340 642.200 6.540 ;
  LAYER VI3 ;
  RECT 642.000 5.940 642.200 6.140 ;
  LAYER VI3 ;
  RECT 1374.360 545.220 1375.220 545.600 ;
  LAYER VI3 ;
  RECT 1374.760 545.280 1374.960 545.480 ;
  LAYER VI3 ;
  RECT 1374.360 545.280 1374.560 545.480 ;
  LAYER VI2 ;
  RECT 1374.360 545.220 1375.220 545.600 ;
  LAYER VI2 ;
  RECT 1374.760 545.280 1374.960 545.480 ;
  LAYER VI2 ;
  RECT 1374.360 545.280 1374.560 545.480 ;
  LAYER VI3 ;
  RECT 1374.360 537.300 1375.220 537.580 ;
  LAYER VI3 ;
  RECT 1374.820 537.300 1375.020 537.500 ;
  LAYER VI3 ;
  RECT 1374.420 537.300 1374.620 537.500 ;
  LAYER VI2 ;
  RECT 1374.360 537.300 1375.220 537.580 ;
  LAYER VI2 ;
  RECT 1374.820 537.300 1375.020 537.500 ;
  LAYER VI2 ;
  RECT 1374.420 537.300 1374.620 537.500 ;
  LAYER VI3 ;
  RECT 1374.360 533.620 1375.220 533.900 ;
  LAYER VI3 ;
  RECT 1374.820 533.620 1375.020 533.820 ;
  LAYER VI3 ;
  RECT 1374.420 533.620 1374.620 533.820 ;
  LAYER VI2 ;
  RECT 1374.360 533.620 1375.220 533.900 ;
  LAYER VI2 ;
  RECT 1374.820 533.620 1375.020 533.820 ;
  LAYER VI2 ;
  RECT 1374.420 533.620 1374.620 533.820 ;
  LAYER VI3 ;
  RECT 1374.360 529.940 1375.220 530.220 ;
  LAYER VI3 ;
  RECT 1374.820 529.940 1375.020 530.140 ;
  LAYER VI3 ;
  RECT 1374.420 529.940 1374.620 530.140 ;
  LAYER VI2 ;
  RECT 1374.360 529.940 1375.220 530.220 ;
  LAYER VI2 ;
  RECT 1374.820 529.940 1375.020 530.140 ;
  LAYER VI2 ;
  RECT 1374.420 529.940 1374.620 530.140 ;
  LAYER VI3 ;
  RECT 1374.360 526.260 1375.220 526.540 ;
  LAYER VI3 ;
  RECT 1374.820 526.260 1375.020 526.460 ;
  LAYER VI3 ;
  RECT 1374.420 526.260 1374.620 526.460 ;
  LAYER VI2 ;
  RECT 1374.360 526.260 1375.220 526.540 ;
  LAYER VI2 ;
  RECT 1374.820 526.260 1375.020 526.460 ;
  LAYER VI2 ;
  RECT 1374.420 526.260 1374.620 526.460 ;
  LAYER VI3 ;
  RECT 1374.360 522.580 1375.220 522.860 ;
  LAYER VI3 ;
  RECT 1374.820 522.580 1375.020 522.780 ;
  LAYER VI3 ;
  RECT 1374.420 522.580 1374.620 522.780 ;
  LAYER VI2 ;
  RECT 1374.360 522.580 1375.220 522.860 ;
  LAYER VI2 ;
  RECT 1374.820 522.580 1375.020 522.780 ;
  LAYER VI2 ;
  RECT 1374.420 522.580 1374.620 522.780 ;
  LAYER VI3 ;
  RECT 1374.360 518.900 1375.220 519.180 ;
  LAYER VI3 ;
  RECT 1374.820 518.900 1375.020 519.100 ;
  LAYER VI3 ;
  RECT 1374.420 518.900 1374.620 519.100 ;
  LAYER VI2 ;
  RECT 1374.360 518.900 1375.220 519.180 ;
  LAYER VI2 ;
  RECT 1374.820 518.900 1375.020 519.100 ;
  LAYER VI2 ;
  RECT 1374.420 518.900 1374.620 519.100 ;
  LAYER VI3 ;
  RECT 1374.360 515.220 1375.220 515.500 ;
  LAYER VI3 ;
  RECT 1374.820 515.220 1375.020 515.420 ;
  LAYER VI3 ;
  RECT 1374.420 515.220 1374.620 515.420 ;
  LAYER VI2 ;
  RECT 1374.360 515.220 1375.220 515.500 ;
  LAYER VI2 ;
  RECT 1374.820 515.220 1375.020 515.420 ;
  LAYER VI2 ;
  RECT 1374.420 515.220 1374.620 515.420 ;
  LAYER VI3 ;
  RECT 1374.360 511.540 1375.220 511.820 ;
  LAYER VI3 ;
  RECT 1374.820 511.540 1375.020 511.740 ;
  LAYER VI3 ;
  RECT 1374.420 511.540 1374.620 511.740 ;
  LAYER VI2 ;
  RECT 1374.360 511.540 1375.220 511.820 ;
  LAYER VI2 ;
  RECT 1374.820 511.540 1375.020 511.740 ;
  LAYER VI2 ;
  RECT 1374.420 511.540 1374.620 511.740 ;
  LAYER VI3 ;
  RECT 1374.360 507.860 1375.220 508.140 ;
  LAYER VI3 ;
  RECT 1374.820 507.860 1375.020 508.060 ;
  LAYER VI3 ;
  RECT 1374.420 507.860 1374.620 508.060 ;
  LAYER VI2 ;
  RECT 1374.360 507.860 1375.220 508.140 ;
  LAYER VI2 ;
  RECT 1374.820 507.860 1375.020 508.060 ;
  LAYER VI2 ;
  RECT 1374.420 507.860 1374.620 508.060 ;
  LAYER VI3 ;
  RECT 1374.360 504.180 1375.220 504.460 ;
  LAYER VI3 ;
  RECT 1374.820 504.180 1375.020 504.380 ;
  LAYER VI3 ;
  RECT 1374.420 504.180 1374.620 504.380 ;
  LAYER VI2 ;
  RECT 1374.360 504.180 1375.220 504.460 ;
  LAYER VI2 ;
  RECT 1374.820 504.180 1375.020 504.380 ;
  LAYER VI2 ;
  RECT 1374.420 504.180 1374.620 504.380 ;
  LAYER VI3 ;
  RECT 1374.360 500.500 1375.220 500.780 ;
  LAYER VI3 ;
  RECT 1374.820 500.500 1375.020 500.700 ;
  LAYER VI3 ;
  RECT 1374.420 500.500 1374.620 500.700 ;
  LAYER VI2 ;
  RECT 1374.360 500.500 1375.220 500.780 ;
  LAYER VI2 ;
  RECT 1374.820 500.500 1375.020 500.700 ;
  LAYER VI2 ;
  RECT 1374.420 500.500 1374.620 500.700 ;
  LAYER VI3 ;
  RECT 1374.360 496.820 1375.220 497.100 ;
  LAYER VI3 ;
  RECT 1374.820 496.820 1375.020 497.020 ;
  LAYER VI3 ;
  RECT 1374.420 496.820 1374.620 497.020 ;
  LAYER VI2 ;
  RECT 1374.360 496.820 1375.220 497.100 ;
  LAYER VI2 ;
  RECT 1374.820 496.820 1375.020 497.020 ;
  LAYER VI2 ;
  RECT 1374.420 496.820 1374.620 497.020 ;
  LAYER VI3 ;
  RECT 1374.360 493.140 1375.220 493.420 ;
  LAYER VI3 ;
  RECT 1374.820 493.140 1375.020 493.340 ;
  LAYER VI3 ;
  RECT 1374.420 493.140 1374.620 493.340 ;
  LAYER VI2 ;
  RECT 1374.360 493.140 1375.220 493.420 ;
  LAYER VI2 ;
  RECT 1374.820 493.140 1375.020 493.340 ;
  LAYER VI2 ;
  RECT 1374.420 493.140 1374.620 493.340 ;
  LAYER VI3 ;
  RECT 1374.360 489.460 1375.220 489.740 ;
  LAYER VI3 ;
  RECT 1374.820 489.460 1375.020 489.660 ;
  LAYER VI3 ;
  RECT 1374.420 489.460 1374.620 489.660 ;
  LAYER VI2 ;
  RECT 1374.360 489.460 1375.220 489.740 ;
  LAYER VI2 ;
  RECT 1374.820 489.460 1375.020 489.660 ;
  LAYER VI2 ;
  RECT 1374.420 489.460 1374.620 489.660 ;
  LAYER VI3 ;
  RECT 1374.360 485.780 1375.220 486.060 ;
  LAYER VI3 ;
  RECT 1374.820 485.780 1375.020 485.980 ;
  LAYER VI3 ;
  RECT 1374.420 485.780 1374.620 485.980 ;
  LAYER VI2 ;
  RECT 1374.360 485.780 1375.220 486.060 ;
  LAYER VI2 ;
  RECT 1374.820 485.780 1375.020 485.980 ;
  LAYER VI2 ;
  RECT 1374.420 485.780 1374.620 485.980 ;
  LAYER VI3 ;
  RECT 1374.360 482.100 1375.220 482.380 ;
  LAYER VI3 ;
  RECT 1374.820 482.100 1375.020 482.300 ;
  LAYER VI3 ;
  RECT 1374.420 482.100 1374.620 482.300 ;
  LAYER VI2 ;
  RECT 1374.360 482.100 1375.220 482.380 ;
  LAYER VI2 ;
  RECT 1374.820 482.100 1375.020 482.300 ;
  LAYER VI2 ;
  RECT 1374.420 482.100 1374.620 482.300 ;
  LAYER VI3 ;
  RECT 1374.360 478.420 1375.220 478.700 ;
  LAYER VI3 ;
  RECT 1374.820 478.420 1375.020 478.620 ;
  LAYER VI3 ;
  RECT 1374.420 478.420 1374.620 478.620 ;
  LAYER VI2 ;
  RECT 1374.360 478.420 1375.220 478.700 ;
  LAYER VI2 ;
  RECT 1374.820 478.420 1375.020 478.620 ;
  LAYER VI2 ;
  RECT 1374.420 478.420 1374.620 478.620 ;
  LAYER VI3 ;
  RECT 1374.360 474.740 1375.220 475.020 ;
  LAYER VI3 ;
  RECT 1374.820 474.740 1375.020 474.940 ;
  LAYER VI3 ;
  RECT 1374.420 474.740 1374.620 474.940 ;
  LAYER VI2 ;
  RECT 1374.360 474.740 1375.220 475.020 ;
  LAYER VI2 ;
  RECT 1374.820 474.740 1375.020 474.940 ;
  LAYER VI2 ;
  RECT 1374.420 474.740 1374.620 474.940 ;
  LAYER VI3 ;
  RECT 1374.360 471.060 1375.220 471.340 ;
  LAYER VI3 ;
  RECT 1374.820 471.060 1375.020 471.260 ;
  LAYER VI3 ;
  RECT 1374.420 471.060 1374.620 471.260 ;
  LAYER VI2 ;
  RECT 1374.360 471.060 1375.220 471.340 ;
  LAYER VI2 ;
  RECT 1374.820 471.060 1375.020 471.260 ;
  LAYER VI2 ;
  RECT 1374.420 471.060 1374.620 471.260 ;
  LAYER VI3 ;
  RECT 1374.360 467.380 1375.220 467.660 ;
  LAYER VI3 ;
  RECT 1374.820 467.380 1375.020 467.580 ;
  LAYER VI3 ;
  RECT 1374.420 467.380 1374.620 467.580 ;
  LAYER VI2 ;
  RECT 1374.360 467.380 1375.220 467.660 ;
  LAYER VI2 ;
  RECT 1374.820 467.380 1375.020 467.580 ;
  LAYER VI2 ;
  RECT 1374.420 467.380 1374.620 467.580 ;
  LAYER VI3 ;
  RECT 1374.360 463.700 1375.220 463.980 ;
  LAYER VI3 ;
  RECT 1374.820 463.700 1375.020 463.900 ;
  LAYER VI3 ;
  RECT 1374.420 463.700 1374.620 463.900 ;
  LAYER VI2 ;
  RECT 1374.360 463.700 1375.220 463.980 ;
  LAYER VI2 ;
  RECT 1374.820 463.700 1375.020 463.900 ;
  LAYER VI2 ;
  RECT 1374.420 463.700 1374.620 463.900 ;
  LAYER VI3 ;
  RECT 1374.360 460.020 1375.220 460.300 ;
  LAYER VI3 ;
  RECT 1374.820 460.020 1375.020 460.220 ;
  LAYER VI3 ;
  RECT 1374.420 460.020 1374.620 460.220 ;
  LAYER VI2 ;
  RECT 1374.360 460.020 1375.220 460.300 ;
  LAYER VI2 ;
  RECT 1374.820 460.020 1375.020 460.220 ;
  LAYER VI2 ;
  RECT 1374.420 460.020 1374.620 460.220 ;
  LAYER VI3 ;
  RECT 1374.360 456.340 1375.220 456.620 ;
  LAYER VI3 ;
  RECT 1374.820 456.340 1375.020 456.540 ;
  LAYER VI3 ;
  RECT 1374.420 456.340 1374.620 456.540 ;
  LAYER VI2 ;
  RECT 1374.360 456.340 1375.220 456.620 ;
  LAYER VI2 ;
  RECT 1374.820 456.340 1375.020 456.540 ;
  LAYER VI2 ;
  RECT 1374.420 456.340 1374.620 456.540 ;
  LAYER VI3 ;
  RECT 1374.360 452.660 1375.220 452.940 ;
  LAYER VI3 ;
  RECT 1374.820 452.660 1375.020 452.860 ;
  LAYER VI3 ;
  RECT 1374.420 452.660 1374.620 452.860 ;
  LAYER VI2 ;
  RECT 1374.360 452.660 1375.220 452.940 ;
  LAYER VI2 ;
  RECT 1374.820 452.660 1375.020 452.860 ;
  LAYER VI2 ;
  RECT 1374.420 452.660 1374.620 452.860 ;
  LAYER VI3 ;
  RECT 1374.360 448.980 1375.220 449.260 ;
  LAYER VI3 ;
  RECT 1374.820 448.980 1375.020 449.180 ;
  LAYER VI3 ;
  RECT 1374.420 448.980 1374.620 449.180 ;
  LAYER VI2 ;
  RECT 1374.360 448.980 1375.220 449.260 ;
  LAYER VI2 ;
  RECT 1374.820 448.980 1375.020 449.180 ;
  LAYER VI2 ;
  RECT 1374.420 448.980 1374.620 449.180 ;
  LAYER VI3 ;
  RECT 1374.360 445.300 1375.220 445.580 ;
  LAYER VI3 ;
  RECT 1374.820 445.300 1375.020 445.500 ;
  LAYER VI3 ;
  RECT 1374.420 445.300 1374.620 445.500 ;
  LAYER VI2 ;
  RECT 1374.360 445.300 1375.220 445.580 ;
  LAYER VI2 ;
  RECT 1374.820 445.300 1375.020 445.500 ;
  LAYER VI2 ;
  RECT 1374.420 445.300 1374.620 445.500 ;
  LAYER VI3 ;
  RECT 1374.360 441.620 1375.220 441.900 ;
  LAYER VI3 ;
  RECT 1374.820 441.620 1375.020 441.820 ;
  LAYER VI3 ;
  RECT 1374.420 441.620 1374.620 441.820 ;
  LAYER VI2 ;
  RECT 1374.360 441.620 1375.220 441.900 ;
  LAYER VI2 ;
  RECT 1374.820 441.620 1375.020 441.820 ;
  LAYER VI2 ;
  RECT 1374.420 441.620 1374.620 441.820 ;
  LAYER VI3 ;
  RECT 1374.360 437.940 1375.220 438.220 ;
  LAYER VI3 ;
  RECT 1374.820 437.940 1375.020 438.140 ;
  LAYER VI3 ;
  RECT 1374.420 437.940 1374.620 438.140 ;
  LAYER VI2 ;
  RECT 1374.360 437.940 1375.220 438.220 ;
  LAYER VI2 ;
  RECT 1374.820 437.940 1375.020 438.140 ;
  LAYER VI2 ;
  RECT 1374.420 437.940 1374.620 438.140 ;
  LAYER VI3 ;
  RECT 1374.360 434.260 1375.220 434.540 ;
  LAYER VI3 ;
  RECT 1374.820 434.260 1375.020 434.460 ;
  LAYER VI3 ;
  RECT 1374.420 434.260 1374.620 434.460 ;
  LAYER VI2 ;
  RECT 1374.360 434.260 1375.220 434.540 ;
  LAYER VI2 ;
  RECT 1374.820 434.260 1375.020 434.460 ;
  LAYER VI2 ;
  RECT 1374.420 434.260 1374.620 434.460 ;
  LAYER VI3 ;
  RECT 1374.360 430.580 1375.220 430.860 ;
  LAYER VI3 ;
  RECT 1374.820 430.580 1375.020 430.780 ;
  LAYER VI3 ;
  RECT 1374.420 430.580 1374.620 430.780 ;
  LAYER VI2 ;
  RECT 1374.360 430.580 1375.220 430.860 ;
  LAYER VI2 ;
  RECT 1374.820 430.580 1375.020 430.780 ;
  LAYER VI2 ;
  RECT 1374.420 430.580 1374.620 430.780 ;
  LAYER VI3 ;
  RECT 1374.360 426.900 1375.220 427.180 ;
  LAYER VI3 ;
  RECT 1374.820 426.900 1375.020 427.100 ;
  LAYER VI3 ;
  RECT 1374.420 426.900 1374.620 427.100 ;
  LAYER VI2 ;
  RECT 1374.360 426.900 1375.220 427.180 ;
  LAYER VI2 ;
  RECT 1374.820 426.900 1375.020 427.100 ;
  LAYER VI2 ;
  RECT 1374.420 426.900 1374.620 427.100 ;
  LAYER VI3 ;
  RECT 1374.360 423.220 1375.220 423.500 ;
  LAYER VI3 ;
  RECT 1374.820 423.220 1375.020 423.420 ;
  LAYER VI3 ;
  RECT 1374.420 423.220 1374.620 423.420 ;
  LAYER VI2 ;
  RECT 1374.360 423.220 1375.220 423.500 ;
  LAYER VI2 ;
  RECT 1374.820 423.220 1375.020 423.420 ;
  LAYER VI2 ;
  RECT 1374.420 423.220 1374.620 423.420 ;
  LAYER VI3 ;
  RECT 1374.360 419.540 1375.220 419.820 ;
  LAYER VI3 ;
  RECT 1374.820 419.540 1375.020 419.740 ;
  LAYER VI3 ;
  RECT 1374.420 419.540 1374.620 419.740 ;
  LAYER VI2 ;
  RECT 1374.360 419.540 1375.220 419.820 ;
  LAYER VI2 ;
  RECT 1374.820 419.540 1375.020 419.740 ;
  LAYER VI2 ;
  RECT 1374.420 419.540 1374.620 419.740 ;
  LAYER VI3 ;
  RECT 1374.360 415.860 1375.220 416.140 ;
  LAYER VI3 ;
  RECT 1374.820 415.860 1375.020 416.060 ;
  LAYER VI3 ;
  RECT 1374.420 415.860 1374.620 416.060 ;
  LAYER VI2 ;
  RECT 1374.360 415.860 1375.220 416.140 ;
  LAYER VI2 ;
  RECT 1374.820 415.860 1375.020 416.060 ;
  LAYER VI2 ;
  RECT 1374.420 415.860 1374.620 416.060 ;
  LAYER VI3 ;
  RECT 1374.360 412.180 1375.220 412.460 ;
  LAYER VI3 ;
  RECT 1374.820 412.180 1375.020 412.380 ;
  LAYER VI3 ;
  RECT 1374.420 412.180 1374.620 412.380 ;
  LAYER VI2 ;
  RECT 1374.360 412.180 1375.220 412.460 ;
  LAYER VI2 ;
  RECT 1374.820 412.180 1375.020 412.380 ;
  LAYER VI2 ;
  RECT 1374.420 412.180 1374.620 412.380 ;
  LAYER VI3 ;
  RECT 1374.360 408.500 1375.220 408.780 ;
  LAYER VI3 ;
  RECT 1374.820 408.500 1375.020 408.700 ;
  LAYER VI3 ;
  RECT 1374.420 408.500 1374.620 408.700 ;
  LAYER VI2 ;
  RECT 1374.360 408.500 1375.220 408.780 ;
  LAYER VI2 ;
  RECT 1374.820 408.500 1375.020 408.700 ;
  LAYER VI2 ;
  RECT 1374.420 408.500 1374.620 408.700 ;
  LAYER VI3 ;
  RECT 1374.360 404.820 1375.220 405.100 ;
  LAYER VI3 ;
  RECT 1374.820 404.820 1375.020 405.020 ;
  LAYER VI3 ;
  RECT 1374.420 404.820 1374.620 405.020 ;
  LAYER VI2 ;
  RECT 1374.360 404.820 1375.220 405.100 ;
  LAYER VI2 ;
  RECT 1374.820 404.820 1375.020 405.020 ;
  LAYER VI2 ;
  RECT 1374.420 404.820 1374.620 405.020 ;
  LAYER VI3 ;
  RECT 1374.360 401.140 1375.220 401.420 ;
  LAYER VI3 ;
  RECT 1374.820 401.140 1375.020 401.340 ;
  LAYER VI3 ;
  RECT 1374.420 401.140 1374.620 401.340 ;
  LAYER VI2 ;
  RECT 1374.360 401.140 1375.220 401.420 ;
  LAYER VI2 ;
  RECT 1374.820 401.140 1375.020 401.340 ;
  LAYER VI2 ;
  RECT 1374.420 401.140 1374.620 401.340 ;
  LAYER VI3 ;
  RECT 1374.360 397.460 1375.220 397.740 ;
  LAYER VI3 ;
  RECT 1374.820 397.460 1375.020 397.660 ;
  LAYER VI3 ;
  RECT 1374.420 397.460 1374.620 397.660 ;
  LAYER VI2 ;
  RECT 1374.360 397.460 1375.220 397.740 ;
  LAYER VI2 ;
  RECT 1374.820 397.460 1375.020 397.660 ;
  LAYER VI2 ;
  RECT 1374.420 397.460 1374.620 397.660 ;
  LAYER VI3 ;
  RECT 1374.360 393.780 1375.220 394.060 ;
  LAYER VI3 ;
  RECT 1374.820 393.780 1375.020 393.980 ;
  LAYER VI3 ;
  RECT 1374.420 393.780 1374.620 393.980 ;
  LAYER VI2 ;
  RECT 1374.360 393.780 1375.220 394.060 ;
  LAYER VI2 ;
  RECT 1374.820 393.780 1375.020 393.980 ;
  LAYER VI2 ;
  RECT 1374.420 393.780 1374.620 393.980 ;
  LAYER VI3 ;
  RECT 1374.360 390.100 1375.220 390.380 ;
  LAYER VI3 ;
  RECT 1374.820 390.100 1375.020 390.300 ;
  LAYER VI3 ;
  RECT 1374.420 390.100 1374.620 390.300 ;
  LAYER VI2 ;
  RECT 1374.360 390.100 1375.220 390.380 ;
  LAYER VI2 ;
  RECT 1374.820 390.100 1375.020 390.300 ;
  LAYER VI2 ;
  RECT 1374.420 390.100 1374.620 390.300 ;
  LAYER VI3 ;
  RECT 1374.360 386.420 1375.220 386.700 ;
  LAYER VI3 ;
  RECT 1374.820 386.420 1375.020 386.620 ;
  LAYER VI3 ;
  RECT 1374.420 386.420 1374.620 386.620 ;
  LAYER VI2 ;
  RECT 1374.360 386.420 1375.220 386.700 ;
  LAYER VI2 ;
  RECT 1374.820 386.420 1375.020 386.620 ;
  LAYER VI2 ;
  RECT 1374.420 386.420 1374.620 386.620 ;
  LAYER VI3 ;
  RECT 1374.360 382.740 1375.220 383.020 ;
  LAYER VI3 ;
  RECT 1374.820 382.740 1375.020 382.940 ;
  LAYER VI3 ;
  RECT 1374.420 382.740 1374.620 382.940 ;
  LAYER VI2 ;
  RECT 1374.360 382.740 1375.220 383.020 ;
  LAYER VI2 ;
  RECT 1374.820 382.740 1375.020 382.940 ;
  LAYER VI2 ;
  RECT 1374.420 382.740 1374.620 382.940 ;
  LAYER VI3 ;
  RECT 1374.360 379.060 1375.220 379.340 ;
  LAYER VI3 ;
  RECT 1374.820 379.060 1375.020 379.260 ;
  LAYER VI3 ;
  RECT 1374.420 379.060 1374.620 379.260 ;
  LAYER VI2 ;
  RECT 1374.360 379.060 1375.220 379.340 ;
  LAYER VI2 ;
  RECT 1374.820 379.060 1375.020 379.260 ;
  LAYER VI2 ;
  RECT 1374.420 379.060 1374.620 379.260 ;
  LAYER VI3 ;
  RECT 1374.360 375.380 1375.220 375.660 ;
  LAYER VI3 ;
  RECT 1374.820 375.380 1375.020 375.580 ;
  LAYER VI3 ;
  RECT 1374.420 375.380 1374.620 375.580 ;
  LAYER VI2 ;
  RECT 1374.360 375.380 1375.220 375.660 ;
  LAYER VI2 ;
  RECT 1374.820 375.380 1375.020 375.580 ;
  LAYER VI2 ;
  RECT 1374.420 375.380 1374.620 375.580 ;
  LAYER VI3 ;
  RECT 1374.360 371.700 1375.220 371.980 ;
  LAYER VI3 ;
  RECT 1374.820 371.700 1375.020 371.900 ;
  LAYER VI3 ;
  RECT 1374.420 371.700 1374.620 371.900 ;
  LAYER VI2 ;
  RECT 1374.360 371.700 1375.220 371.980 ;
  LAYER VI2 ;
  RECT 1374.820 371.700 1375.020 371.900 ;
  LAYER VI2 ;
  RECT 1374.420 371.700 1374.620 371.900 ;
  LAYER VI3 ;
  RECT 1374.360 368.020 1375.220 368.300 ;
  LAYER VI3 ;
  RECT 1374.820 368.020 1375.020 368.220 ;
  LAYER VI3 ;
  RECT 1374.420 368.020 1374.620 368.220 ;
  LAYER VI2 ;
  RECT 1374.360 368.020 1375.220 368.300 ;
  LAYER VI2 ;
  RECT 1374.820 368.020 1375.020 368.220 ;
  LAYER VI2 ;
  RECT 1374.420 368.020 1374.620 368.220 ;
  LAYER VI3 ;
  RECT 1374.360 364.340 1375.220 364.620 ;
  LAYER VI3 ;
  RECT 1374.820 364.340 1375.020 364.540 ;
  LAYER VI3 ;
  RECT 1374.420 364.340 1374.620 364.540 ;
  LAYER VI2 ;
  RECT 1374.360 364.340 1375.220 364.620 ;
  LAYER VI2 ;
  RECT 1374.820 364.340 1375.020 364.540 ;
  LAYER VI2 ;
  RECT 1374.420 364.340 1374.620 364.540 ;
  LAYER VI3 ;
  RECT 1374.360 360.660 1375.220 360.940 ;
  LAYER VI3 ;
  RECT 1374.820 360.660 1375.020 360.860 ;
  LAYER VI3 ;
  RECT 1374.420 360.660 1374.620 360.860 ;
  LAYER VI2 ;
  RECT 1374.360 360.660 1375.220 360.940 ;
  LAYER VI2 ;
  RECT 1374.820 360.660 1375.020 360.860 ;
  LAYER VI2 ;
  RECT 1374.420 360.660 1374.620 360.860 ;
  LAYER VI3 ;
  RECT 1374.360 356.980 1375.220 357.260 ;
  LAYER VI3 ;
  RECT 1374.820 356.980 1375.020 357.180 ;
  LAYER VI3 ;
  RECT 1374.420 356.980 1374.620 357.180 ;
  LAYER VI2 ;
  RECT 1374.360 356.980 1375.220 357.260 ;
  LAYER VI2 ;
  RECT 1374.820 356.980 1375.020 357.180 ;
  LAYER VI2 ;
  RECT 1374.420 356.980 1374.620 357.180 ;
  LAYER VI3 ;
  RECT 1374.360 353.300 1375.220 353.580 ;
  LAYER VI3 ;
  RECT 1374.820 353.300 1375.020 353.500 ;
  LAYER VI3 ;
  RECT 1374.420 353.300 1374.620 353.500 ;
  LAYER VI2 ;
  RECT 1374.360 353.300 1375.220 353.580 ;
  LAYER VI2 ;
  RECT 1374.820 353.300 1375.020 353.500 ;
  LAYER VI2 ;
  RECT 1374.420 353.300 1374.620 353.500 ;
  LAYER VI3 ;
  RECT 1374.360 349.620 1375.220 349.900 ;
  LAYER VI3 ;
  RECT 1374.820 349.620 1375.020 349.820 ;
  LAYER VI3 ;
  RECT 1374.420 349.620 1374.620 349.820 ;
  LAYER VI2 ;
  RECT 1374.360 349.620 1375.220 349.900 ;
  LAYER VI2 ;
  RECT 1374.820 349.620 1375.020 349.820 ;
  LAYER VI2 ;
  RECT 1374.420 349.620 1374.620 349.820 ;
  LAYER VI3 ;
  RECT 1374.360 345.940 1375.220 346.220 ;
  LAYER VI3 ;
  RECT 1374.820 345.940 1375.020 346.140 ;
  LAYER VI3 ;
  RECT 1374.420 345.940 1374.620 346.140 ;
  LAYER VI2 ;
  RECT 1374.360 345.940 1375.220 346.220 ;
  LAYER VI2 ;
  RECT 1374.820 345.940 1375.020 346.140 ;
  LAYER VI2 ;
  RECT 1374.420 345.940 1374.620 346.140 ;
  LAYER VI3 ;
  RECT 1374.360 342.260 1375.220 342.540 ;
  LAYER VI3 ;
  RECT 1374.820 342.260 1375.020 342.460 ;
  LAYER VI3 ;
  RECT 1374.420 342.260 1374.620 342.460 ;
  LAYER VI2 ;
  RECT 1374.360 342.260 1375.220 342.540 ;
  LAYER VI2 ;
  RECT 1374.820 342.260 1375.020 342.460 ;
  LAYER VI2 ;
  RECT 1374.420 342.260 1374.620 342.460 ;
  LAYER VI3 ;
  RECT 1374.360 338.580 1375.220 338.860 ;
  LAYER VI3 ;
  RECT 1374.820 338.580 1375.020 338.780 ;
  LAYER VI3 ;
  RECT 1374.420 338.580 1374.620 338.780 ;
  LAYER VI2 ;
  RECT 1374.360 338.580 1375.220 338.860 ;
  LAYER VI2 ;
  RECT 1374.820 338.580 1375.020 338.780 ;
  LAYER VI2 ;
  RECT 1374.420 338.580 1374.620 338.780 ;
  LAYER VI3 ;
  RECT 1374.360 334.900 1375.220 335.180 ;
  LAYER VI3 ;
  RECT 1374.820 334.900 1375.020 335.100 ;
  LAYER VI3 ;
  RECT 1374.420 334.900 1374.620 335.100 ;
  LAYER VI2 ;
  RECT 1374.360 334.900 1375.220 335.180 ;
  LAYER VI2 ;
  RECT 1374.820 334.900 1375.020 335.100 ;
  LAYER VI2 ;
  RECT 1374.420 334.900 1374.620 335.100 ;
  LAYER VI3 ;
  RECT 1374.360 331.220 1375.220 331.500 ;
  LAYER VI3 ;
  RECT 1374.820 331.220 1375.020 331.420 ;
  LAYER VI3 ;
  RECT 1374.420 331.220 1374.620 331.420 ;
  LAYER VI2 ;
  RECT 1374.360 331.220 1375.220 331.500 ;
  LAYER VI2 ;
  RECT 1374.820 331.220 1375.020 331.420 ;
  LAYER VI2 ;
  RECT 1374.420 331.220 1374.620 331.420 ;
  LAYER VI3 ;
  RECT 1374.360 327.540 1375.220 327.820 ;
  LAYER VI3 ;
  RECT 1374.820 327.540 1375.020 327.740 ;
  LAYER VI3 ;
  RECT 1374.420 327.540 1374.620 327.740 ;
  LAYER VI2 ;
  RECT 1374.360 327.540 1375.220 327.820 ;
  LAYER VI2 ;
  RECT 1374.820 327.540 1375.020 327.740 ;
  LAYER VI2 ;
  RECT 1374.420 327.540 1374.620 327.740 ;
  LAYER VI3 ;
  RECT 1374.360 323.860 1375.220 324.140 ;
  LAYER VI3 ;
  RECT 1374.820 323.860 1375.020 324.060 ;
  LAYER VI3 ;
  RECT 1374.420 323.860 1374.620 324.060 ;
  LAYER VI2 ;
  RECT 1374.360 323.860 1375.220 324.140 ;
  LAYER VI2 ;
  RECT 1374.820 323.860 1375.020 324.060 ;
  LAYER VI2 ;
  RECT 1374.420 323.860 1374.620 324.060 ;
  LAYER VI3 ;
  RECT 1374.360 320.180 1375.220 320.460 ;
  LAYER VI3 ;
  RECT 1374.820 320.180 1375.020 320.380 ;
  LAYER VI3 ;
  RECT 1374.420 320.180 1374.620 320.380 ;
  LAYER VI2 ;
  RECT 1374.360 320.180 1375.220 320.460 ;
  LAYER VI2 ;
  RECT 1374.820 320.180 1375.020 320.380 ;
  LAYER VI2 ;
  RECT 1374.420 320.180 1374.620 320.380 ;
  LAYER VI3 ;
  RECT 1374.360 316.500 1375.220 316.780 ;
  LAYER VI3 ;
  RECT 1374.820 316.500 1375.020 316.700 ;
  LAYER VI3 ;
  RECT 1374.420 316.500 1374.620 316.700 ;
  LAYER VI2 ;
  RECT 1374.360 316.500 1375.220 316.780 ;
  LAYER VI2 ;
  RECT 1374.820 316.500 1375.020 316.700 ;
  LAYER VI2 ;
  RECT 1374.420 316.500 1374.620 316.700 ;
  LAYER VI3 ;
  RECT 1374.360 312.820 1375.220 313.100 ;
  LAYER VI3 ;
  RECT 1374.820 312.820 1375.020 313.020 ;
  LAYER VI3 ;
  RECT 1374.420 312.820 1374.620 313.020 ;
  LAYER VI2 ;
  RECT 1374.360 312.820 1375.220 313.100 ;
  LAYER VI2 ;
  RECT 1374.820 312.820 1375.020 313.020 ;
  LAYER VI2 ;
  RECT 1374.420 312.820 1374.620 313.020 ;
  LAYER VI3 ;
  RECT 1374.360 309.140 1375.220 309.420 ;
  LAYER VI3 ;
  RECT 1374.820 309.140 1375.020 309.340 ;
  LAYER VI3 ;
  RECT 1374.420 309.140 1374.620 309.340 ;
  LAYER VI2 ;
  RECT 1374.360 309.140 1375.220 309.420 ;
  LAYER VI2 ;
  RECT 1374.820 309.140 1375.020 309.340 ;
  LAYER VI2 ;
  RECT 1374.420 309.140 1374.620 309.340 ;
  LAYER VI3 ;
  RECT 1374.360 305.460 1375.220 305.740 ;
  LAYER VI3 ;
  RECT 1374.820 305.460 1375.020 305.660 ;
  LAYER VI3 ;
  RECT 1374.420 305.460 1374.620 305.660 ;
  LAYER VI2 ;
  RECT 1374.360 305.460 1375.220 305.740 ;
  LAYER VI2 ;
  RECT 1374.820 305.460 1375.020 305.660 ;
  LAYER VI2 ;
  RECT 1374.420 305.460 1374.620 305.660 ;
  LAYER VI3 ;
  RECT 1374.360 301.780 1375.220 302.060 ;
  LAYER VI3 ;
  RECT 1374.820 301.780 1375.020 301.980 ;
  LAYER VI3 ;
  RECT 1374.420 301.780 1374.620 301.980 ;
  LAYER VI2 ;
  RECT 1374.360 301.780 1375.220 302.060 ;
  LAYER VI2 ;
  RECT 1374.820 301.780 1375.020 301.980 ;
  LAYER VI2 ;
  RECT 1374.420 301.780 1374.620 301.980 ;
  LAYER VI3 ;
  RECT 1374.360 298.100 1375.220 298.380 ;
  LAYER VI3 ;
  RECT 1374.820 298.100 1375.020 298.300 ;
  LAYER VI3 ;
  RECT 1374.420 298.100 1374.620 298.300 ;
  LAYER VI2 ;
  RECT 1374.360 298.100 1375.220 298.380 ;
  LAYER VI2 ;
  RECT 1374.820 298.100 1375.020 298.300 ;
  LAYER VI2 ;
  RECT 1374.420 298.100 1374.620 298.300 ;
  LAYER VI3 ;
  RECT 1374.360 294.420 1375.220 294.700 ;
  LAYER VI3 ;
  RECT 1374.820 294.420 1375.020 294.620 ;
  LAYER VI3 ;
  RECT 1374.420 294.420 1374.620 294.620 ;
  LAYER VI2 ;
  RECT 1374.360 294.420 1375.220 294.700 ;
  LAYER VI2 ;
  RECT 1374.820 294.420 1375.020 294.620 ;
  LAYER VI2 ;
  RECT 1374.420 294.420 1374.620 294.620 ;
  LAYER VI3 ;
  RECT 1374.360 290.740 1375.220 291.020 ;
  LAYER VI3 ;
  RECT 1374.820 290.740 1375.020 290.940 ;
  LAYER VI3 ;
  RECT 1374.420 290.740 1374.620 290.940 ;
  LAYER VI2 ;
  RECT 1374.360 290.740 1375.220 291.020 ;
  LAYER VI2 ;
  RECT 1374.820 290.740 1375.020 290.940 ;
  LAYER VI2 ;
  RECT 1374.420 290.740 1374.620 290.940 ;
  LAYER VI3 ;
  RECT 1374.360 287.060 1375.220 287.340 ;
  LAYER VI3 ;
  RECT 1374.820 287.060 1375.020 287.260 ;
  LAYER VI3 ;
  RECT 1374.420 287.060 1374.620 287.260 ;
  LAYER VI2 ;
  RECT 1374.360 287.060 1375.220 287.340 ;
  LAYER VI2 ;
  RECT 1374.820 287.060 1375.020 287.260 ;
  LAYER VI2 ;
  RECT 1374.420 287.060 1374.620 287.260 ;
  LAYER VI3 ;
  RECT 1374.360 283.380 1375.220 283.660 ;
  LAYER VI3 ;
  RECT 1374.820 283.380 1375.020 283.580 ;
  LAYER VI3 ;
  RECT 1374.420 283.380 1374.620 283.580 ;
  LAYER VI2 ;
  RECT 1374.360 283.380 1375.220 283.660 ;
  LAYER VI2 ;
  RECT 1374.820 283.380 1375.020 283.580 ;
  LAYER VI2 ;
  RECT 1374.420 283.380 1374.620 283.580 ;
  LAYER VI3 ;
  RECT 1374.360 279.700 1375.220 279.980 ;
  LAYER VI3 ;
  RECT 1374.820 279.700 1375.020 279.900 ;
  LAYER VI3 ;
  RECT 1374.420 279.700 1374.620 279.900 ;
  LAYER VI2 ;
  RECT 1374.360 279.700 1375.220 279.980 ;
  LAYER VI2 ;
  RECT 1374.820 279.700 1375.020 279.900 ;
  LAYER VI2 ;
  RECT 1374.420 279.700 1374.620 279.900 ;
  LAYER VI3 ;
  RECT 1374.360 276.020 1375.220 276.300 ;
  LAYER VI3 ;
  RECT 1374.820 276.020 1375.020 276.220 ;
  LAYER VI3 ;
  RECT 1374.420 276.020 1374.620 276.220 ;
  LAYER VI2 ;
  RECT 1374.360 276.020 1375.220 276.300 ;
  LAYER VI2 ;
  RECT 1374.820 276.020 1375.020 276.220 ;
  LAYER VI2 ;
  RECT 1374.420 276.020 1374.620 276.220 ;
  LAYER VI3 ;
  RECT 1374.360 272.340 1375.220 272.620 ;
  LAYER VI3 ;
  RECT 1374.820 272.340 1375.020 272.540 ;
  LAYER VI3 ;
  RECT 1374.420 272.340 1374.620 272.540 ;
  LAYER VI2 ;
  RECT 1374.360 272.340 1375.220 272.620 ;
  LAYER VI2 ;
  RECT 1374.820 272.340 1375.020 272.540 ;
  LAYER VI2 ;
  RECT 1374.420 272.340 1374.620 272.540 ;
  LAYER VI3 ;
  RECT 1374.360 268.660 1375.220 268.940 ;
  LAYER VI3 ;
  RECT 1374.820 268.660 1375.020 268.860 ;
  LAYER VI3 ;
  RECT 1374.420 268.660 1374.620 268.860 ;
  LAYER VI2 ;
  RECT 1374.360 268.660 1375.220 268.940 ;
  LAYER VI2 ;
  RECT 1374.820 268.660 1375.020 268.860 ;
  LAYER VI2 ;
  RECT 1374.420 268.660 1374.620 268.860 ;
  LAYER VI3 ;
  RECT 1374.360 264.980 1375.220 265.260 ;
  LAYER VI3 ;
  RECT 1374.820 264.980 1375.020 265.180 ;
  LAYER VI3 ;
  RECT 1374.420 264.980 1374.620 265.180 ;
  LAYER VI2 ;
  RECT 1374.360 264.980 1375.220 265.260 ;
  LAYER VI2 ;
  RECT 1374.820 264.980 1375.020 265.180 ;
  LAYER VI2 ;
  RECT 1374.420 264.980 1374.620 265.180 ;
  LAYER VI3 ;
  RECT 1374.360 261.300 1375.220 261.580 ;
  LAYER VI3 ;
  RECT 1374.820 261.300 1375.020 261.500 ;
  LAYER VI3 ;
  RECT 1374.420 261.300 1374.620 261.500 ;
  LAYER VI2 ;
  RECT 1374.360 261.300 1375.220 261.580 ;
  LAYER VI2 ;
  RECT 1374.820 261.300 1375.020 261.500 ;
  LAYER VI2 ;
  RECT 1374.420 261.300 1374.620 261.500 ;
  LAYER VI3 ;
  RECT 1374.360 257.620 1375.220 257.900 ;
  LAYER VI3 ;
  RECT 1374.820 257.620 1375.020 257.820 ;
  LAYER VI3 ;
  RECT 1374.420 257.620 1374.620 257.820 ;
  LAYER VI2 ;
  RECT 1374.360 257.620 1375.220 257.900 ;
  LAYER VI2 ;
  RECT 1374.820 257.620 1375.020 257.820 ;
  LAYER VI2 ;
  RECT 1374.420 257.620 1374.620 257.820 ;
  LAYER VI3 ;
  RECT 1374.360 253.940 1375.220 254.220 ;
  LAYER VI3 ;
  RECT 1374.820 253.940 1375.020 254.140 ;
  LAYER VI3 ;
  RECT 1374.420 253.940 1374.620 254.140 ;
  LAYER VI2 ;
  RECT 1374.360 253.940 1375.220 254.220 ;
  LAYER VI2 ;
  RECT 1374.820 253.940 1375.020 254.140 ;
  LAYER VI2 ;
  RECT 1374.420 253.940 1374.620 254.140 ;
  LAYER VI3 ;
  RECT 1374.360 250.260 1375.220 250.540 ;
  LAYER VI3 ;
  RECT 1374.820 250.260 1375.020 250.460 ;
  LAYER VI3 ;
  RECT 1374.420 250.260 1374.620 250.460 ;
  LAYER VI2 ;
  RECT 1374.360 250.260 1375.220 250.540 ;
  LAYER VI2 ;
  RECT 1374.820 250.260 1375.020 250.460 ;
  LAYER VI2 ;
  RECT 1374.420 250.260 1374.620 250.460 ;
  LAYER VI3 ;
  RECT 1374.360 246.580 1375.220 246.860 ;
  LAYER VI3 ;
  RECT 1374.820 246.580 1375.020 246.780 ;
  LAYER VI3 ;
  RECT 1374.420 246.580 1374.620 246.780 ;
  LAYER VI2 ;
  RECT 1374.360 246.580 1375.220 246.860 ;
  LAYER VI2 ;
  RECT 1374.820 246.580 1375.020 246.780 ;
  LAYER VI2 ;
  RECT 1374.420 246.580 1374.620 246.780 ;
  LAYER VI3 ;
  RECT 1374.360 242.900 1375.220 243.180 ;
  LAYER VI3 ;
  RECT 1374.820 242.900 1375.020 243.100 ;
  LAYER VI3 ;
  RECT 1374.420 242.900 1374.620 243.100 ;
  LAYER VI2 ;
  RECT 1374.360 242.900 1375.220 243.180 ;
  LAYER VI2 ;
  RECT 1374.820 242.900 1375.020 243.100 ;
  LAYER VI2 ;
  RECT 1374.420 242.900 1374.620 243.100 ;
  LAYER VI3 ;
  RECT 1374.360 239.220 1375.220 239.500 ;
  LAYER VI3 ;
  RECT 1374.820 239.220 1375.020 239.420 ;
  LAYER VI3 ;
  RECT 1374.420 239.220 1374.620 239.420 ;
  LAYER VI2 ;
  RECT 1374.360 239.220 1375.220 239.500 ;
  LAYER VI2 ;
  RECT 1374.820 239.220 1375.020 239.420 ;
  LAYER VI2 ;
  RECT 1374.420 239.220 1374.620 239.420 ;
  LAYER VI3 ;
  RECT 1374.360 235.540 1375.220 235.820 ;
  LAYER VI3 ;
  RECT 1374.820 235.540 1375.020 235.740 ;
  LAYER VI3 ;
  RECT 1374.420 235.540 1374.620 235.740 ;
  LAYER VI2 ;
  RECT 1374.360 235.540 1375.220 235.820 ;
  LAYER VI2 ;
  RECT 1374.820 235.540 1375.020 235.740 ;
  LAYER VI2 ;
  RECT 1374.420 235.540 1374.620 235.740 ;
  LAYER VI3 ;
  RECT 1374.360 231.860 1375.220 232.140 ;
  LAYER VI3 ;
  RECT 1374.820 231.860 1375.020 232.060 ;
  LAYER VI3 ;
  RECT 1374.420 231.860 1374.620 232.060 ;
  LAYER VI2 ;
  RECT 1374.360 231.860 1375.220 232.140 ;
  LAYER VI2 ;
  RECT 1374.820 231.860 1375.020 232.060 ;
  LAYER VI2 ;
  RECT 1374.420 231.860 1374.620 232.060 ;
  LAYER VI3 ;
  RECT 1374.360 228.180 1375.220 228.460 ;
  LAYER VI3 ;
  RECT 1374.820 228.180 1375.020 228.380 ;
  LAYER VI3 ;
  RECT 1374.420 228.180 1374.620 228.380 ;
  LAYER VI2 ;
  RECT 1374.360 228.180 1375.220 228.460 ;
  LAYER VI2 ;
  RECT 1374.820 228.180 1375.020 228.380 ;
  LAYER VI2 ;
  RECT 1374.420 228.180 1374.620 228.380 ;
  LAYER VI3 ;
  RECT 1374.360 224.500 1375.220 224.780 ;
  LAYER VI3 ;
  RECT 1374.820 224.500 1375.020 224.700 ;
  LAYER VI3 ;
  RECT 1374.420 224.500 1374.620 224.700 ;
  LAYER VI2 ;
  RECT 1374.360 224.500 1375.220 224.780 ;
  LAYER VI2 ;
  RECT 1374.820 224.500 1375.020 224.700 ;
  LAYER VI2 ;
  RECT 1374.420 224.500 1374.620 224.700 ;
  LAYER VI3 ;
  RECT 1374.360 220.820 1375.220 221.100 ;
  LAYER VI3 ;
  RECT 1374.820 220.820 1375.020 221.020 ;
  LAYER VI3 ;
  RECT 1374.420 220.820 1374.620 221.020 ;
  LAYER VI2 ;
  RECT 1374.360 220.820 1375.220 221.100 ;
  LAYER VI2 ;
  RECT 1374.820 220.820 1375.020 221.020 ;
  LAYER VI2 ;
  RECT 1374.420 220.820 1374.620 221.020 ;
  LAYER VI3 ;
  RECT 1374.360 217.140 1375.220 217.420 ;
  LAYER VI3 ;
  RECT 1374.820 217.140 1375.020 217.340 ;
  LAYER VI3 ;
  RECT 1374.420 217.140 1374.620 217.340 ;
  LAYER VI2 ;
  RECT 1374.360 217.140 1375.220 217.420 ;
  LAYER VI2 ;
  RECT 1374.820 217.140 1375.020 217.340 ;
  LAYER VI2 ;
  RECT 1374.420 217.140 1374.620 217.340 ;
  LAYER VI3 ;
  RECT 1374.360 213.460 1375.220 213.740 ;
  LAYER VI3 ;
  RECT 1374.820 213.460 1375.020 213.660 ;
  LAYER VI3 ;
  RECT 1374.420 213.460 1374.620 213.660 ;
  LAYER VI2 ;
  RECT 1374.360 213.460 1375.220 213.740 ;
  LAYER VI2 ;
  RECT 1374.820 213.460 1375.020 213.660 ;
  LAYER VI2 ;
  RECT 1374.420 213.460 1374.620 213.660 ;
  LAYER VI3 ;
  RECT 1374.360 209.780 1375.220 210.060 ;
  LAYER VI3 ;
  RECT 1374.820 209.780 1375.020 209.980 ;
  LAYER VI3 ;
  RECT 1374.420 209.780 1374.620 209.980 ;
  LAYER VI2 ;
  RECT 1374.360 209.780 1375.220 210.060 ;
  LAYER VI2 ;
  RECT 1374.820 209.780 1375.020 209.980 ;
  LAYER VI2 ;
  RECT 1374.420 209.780 1374.620 209.980 ;
  LAYER VI3 ;
  RECT 1374.360 206.100 1375.220 206.380 ;
  LAYER VI3 ;
  RECT 1374.820 206.100 1375.020 206.300 ;
  LAYER VI3 ;
  RECT 1374.420 206.100 1374.620 206.300 ;
  LAYER VI2 ;
  RECT 1374.360 206.100 1375.220 206.380 ;
  LAYER VI2 ;
  RECT 1374.820 206.100 1375.020 206.300 ;
  LAYER VI2 ;
  RECT 1374.420 206.100 1374.620 206.300 ;
  LAYER VI3 ;
  RECT 1374.360 202.420 1375.220 202.700 ;
  LAYER VI3 ;
  RECT 1374.820 202.420 1375.020 202.620 ;
  LAYER VI3 ;
  RECT 1374.420 202.420 1374.620 202.620 ;
  LAYER VI2 ;
  RECT 1374.360 202.420 1375.220 202.700 ;
  LAYER VI2 ;
  RECT 1374.820 202.420 1375.020 202.620 ;
  LAYER VI2 ;
  RECT 1374.420 202.420 1374.620 202.620 ;
  LAYER VI3 ;
  RECT 1374.360 198.740 1375.220 199.020 ;
  LAYER VI3 ;
  RECT 1374.820 198.740 1375.020 198.940 ;
  LAYER VI3 ;
  RECT 1374.420 198.740 1374.620 198.940 ;
  LAYER VI2 ;
  RECT 1374.360 198.740 1375.220 199.020 ;
  LAYER VI2 ;
  RECT 1374.820 198.740 1375.020 198.940 ;
  LAYER VI2 ;
  RECT 1374.420 198.740 1374.620 198.940 ;
  LAYER VI3 ;
  RECT 1374.360 195.060 1375.220 195.340 ;
  LAYER VI3 ;
  RECT 1374.820 195.060 1375.020 195.260 ;
  LAYER VI3 ;
  RECT 1374.420 195.060 1374.620 195.260 ;
  LAYER VI2 ;
  RECT 1374.360 195.060 1375.220 195.340 ;
  LAYER VI2 ;
  RECT 1374.820 195.060 1375.020 195.260 ;
  LAYER VI2 ;
  RECT 1374.420 195.060 1374.620 195.260 ;
  LAYER VI3 ;
  RECT 1374.360 191.380 1375.220 191.660 ;
  LAYER VI3 ;
  RECT 1374.820 191.380 1375.020 191.580 ;
  LAYER VI3 ;
  RECT 1374.420 191.380 1374.620 191.580 ;
  LAYER VI2 ;
  RECT 1374.360 191.380 1375.220 191.660 ;
  LAYER VI2 ;
  RECT 1374.820 191.380 1375.020 191.580 ;
  LAYER VI2 ;
  RECT 1374.420 191.380 1374.620 191.580 ;
  LAYER VI3 ;
  RECT 1374.360 187.700 1375.220 187.980 ;
  LAYER VI3 ;
  RECT 1374.820 187.700 1375.020 187.900 ;
  LAYER VI3 ;
  RECT 1374.420 187.700 1374.620 187.900 ;
  LAYER VI2 ;
  RECT 1374.360 187.700 1375.220 187.980 ;
  LAYER VI2 ;
  RECT 1374.820 187.700 1375.020 187.900 ;
  LAYER VI2 ;
  RECT 1374.420 187.700 1374.620 187.900 ;
  LAYER VI3 ;
  RECT 1374.360 184.020 1375.220 184.300 ;
  LAYER VI3 ;
  RECT 1374.820 184.020 1375.020 184.220 ;
  LAYER VI3 ;
  RECT 1374.420 184.020 1374.620 184.220 ;
  LAYER VI2 ;
  RECT 1374.360 184.020 1375.220 184.300 ;
  LAYER VI2 ;
  RECT 1374.820 184.020 1375.020 184.220 ;
  LAYER VI2 ;
  RECT 1374.420 184.020 1374.620 184.220 ;
  LAYER VI3 ;
  RECT 1374.360 180.340 1375.220 180.620 ;
  LAYER VI3 ;
  RECT 1374.820 180.340 1375.020 180.540 ;
  LAYER VI3 ;
  RECT 1374.420 180.340 1374.620 180.540 ;
  LAYER VI2 ;
  RECT 1374.360 180.340 1375.220 180.620 ;
  LAYER VI2 ;
  RECT 1374.820 180.340 1375.020 180.540 ;
  LAYER VI2 ;
  RECT 1374.420 180.340 1374.620 180.540 ;
  LAYER VI3 ;
  RECT 1374.360 176.660 1375.220 176.940 ;
  LAYER VI3 ;
  RECT 1374.820 176.660 1375.020 176.860 ;
  LAYER VI3 ;
  RECT 1374.420 176.660 1374.620 176.860 ;
  LAYER VI2 ;
  RECT 1374.360 176.660 1375.220 176.940 ;
  LAYER VI2 ;
  RECT 1374.820 176.660 1375.020 176.860 ;
  LAYER VI2 ;
  RECT 1374.420 176.660 1374.620 176.860 ;
  LAYER VI3 ;
  RECT 1374.360 172.980 1375.220 173.260 ;
  LAYER VI3 ;
  RECT 1374.820 172.980 1375.020 173.180 ;
  LAYER VI3 ;
  RECT 1374.420 172.980 1374.620 173.180 ;
  LAYER VI2 ;
  RECT 1374.360 172.980 1375.220 173.260 ;
  LAYER VI2 ;
  RECT 1374.820 172.980 1375.020 173.180 ;
  LAYER VI2 ;
  RECT 1374.420 172.980 1374.620 173.180 ;
  LAYER VI3 ;
  RECT 1374.360 169.300 1375.220 169.580 ;
  LAYER VI3 ;
  RECT 1374.820 169.300 1375.020 169.500 ;
  LAYER VI3 ;
  RECT 1374.420 169.300 1374.620 169.500 ;
  LAYER VI2 ;
  RECT 1374.360 169.300 1375.220 169.580 ;
  LAYER VI2 ;
  RECT 1374.820 169.300 1375.020 169.500 ;
  LAYER VI2 ;
  RECT 1374.420 169.300 1374.620 169.500 ;
  LAYER VI3 ;
  RECT 1374.360 165.620 1375.220 165.900 ;
  LAYER VI3 ;
  RECT 1374.820 165.620 1375.020 165.820 ;
  LAYER VI3 ;
  RECT 1374.420 165.620 1374.620 165.820 ;
  LAYER VI2 ;
  RECT 1374.360 165.620 1375.220 165.900 ;
  LAYER VI2 ;
  RECT 1374.820 165.620 1375.020 165.820 ;
  LAYER VI2 ;
  RECT 1374.420 165.620 1374.620 165.820 ;
  LAYER VI3 ;
  RECT 1374.360 161.940 1375.220 162.220 ;
  LAYER VI3 ;
  RECT 1374.820 161.940 1375.020 162.140 ;
  LAYER VI3 ;
  RECT 1374.420 161.940 1374.620 162.140 ;
  LAYER VI2 ;
  RECT 1374.360 161.940 1375.220 162.220 ;
  LAYER VI2 ;
  RECT 1374.820 161.940 1375.020 162.140 ;
  LAYER VI2 ;
  RECT 1374.420 161.940 1374.620 162.140 ;
  LAYER VI3 ;
  RECT 1374.360 158.260 1375.220 158.540 ;
  LAYER VI3 ;
  RECT 1374.820 158.260 1375.020 158.460 ;
  LAYER VI3 ;
  RECT 1374.420 158.260 1374.620 158.460 ;
  LAYER VI2 ;
  RECT 1374.360 158.260 1375.220 158.540 ;
  LAYER VI2 ;
  RECT 1374.820 158.260 1375.020 158.460 ;
  LAYER VI2 ;
  RECT 1374.420 158.260 1374.620 158.460 ;
  LAYER VI3 ;
  RECT 1374.360 154.580 1375.220 154.860 ;
  LAYER VI3 ;
  RECT 1374.820 154.580 1375.020 154.780 ;
  LAYER VI3 ;
  RECT 1374.420 154.580 1374.620 154.780 ;
  LAYER VI2 ;
  RECT 1374.360 154.580 1375.220 154.860 ;
  LAYER VI2 ;
  RECT 1374.820 154.580 1375.020 154.780 ;
  LAYER VI2 ;
  RECT 1374.420 154.580 1374.620 154.780 ;
  LAYER VI3 ;
  RECT 1374.360 150.900 1375.220 151.180 ;
  LAYER VI3 ;
  RECT 1374.820 150.900 1375.020 151.100 ;
  LAYER VI3 ;
  RECT 1374.420 150.900 1374.620 151.100 ;
  LAYER VI2 ;
  RECT 1374.360 150.900 1375.220 151.180 ;
  LAYER VI2 ;
  RECT 1374.820 150.900 1375.020 151.100 ;
  LAYER VI2 ;
  RECT 1374.420 150.900 1374.620 151.100 ;
  LAYER VI3 ;
  RECT 1374.360 147.220 1375.220 147.500 ;
  LAYER VI3 ;
  RECT 1374.820 147.220 1375.020 147.420 ;
  LAYER VI3 ;
  RECT 1374.420 147.220 1374.620 147.420 ;
  LAYER VI2 ;
  RECT 1374.360 147.220 1375.220 147.500 ;
  LAYER VI2 ;
  RECT 1374.820 147.220 1375.020 147.420 ;
  LAYER VI2 ;
  RECT 1374.420 147.220 1374.620 147.420 ;
  LAYER VI3 ;
  RECT 1374.360 143.540 1375.220 143.820 ;
  LAYER VI3 ;
  RECT 1374.820 143.540 1375.020 143.740 ;
  LAYER VI3 ;
  RECT 1374.420 143.540 1374.620 143.740 ;
  LAYER VI2 ;
  RECT 1374.360 143.540 1375.220 143.820 ;
  LAYER VI2 ;
  RECT 1374.820 143.540 1375.020 143.740 ;
  LAYER VI2 ;
  RECT 1374.420 143.540 1374.620 143.740 ;
  LAYER VI3 ;
  RECT 1374.360 139.860 1375.220 140.140 ;
  LAYER VI3 ;
  RECT 1374.820 139.860 1375.020 140.060 ;
  LAYER VI3 ;
  RECT 1374.420 139.860 1374.620 140.060 ;
  LAYER VI2 ;
  RECT 1374.360 139.860 1375.220 140.140 ;
  LAYER VI2 ;
  RECT 1374.820 139.860 1375.020 140.060 ;
  LAYER VI2 ;
  RECT 1374.420 139.860 1374.620 140.060 ;
  LAYER VI3 ;
  RECT 1374.360 136.180 1375.220 136.460 ;
  LAYER VI3 ;
  RECT 1374.820 136.180 1375.020 136.380 ;
  LAYER VI3 ;
  RECT 1374.420 136.180 1374.620 136.380 ;
  LAYER VI2 ;
  RECT 1374.360 136.180 1375.220 136.460 ;
  LAYER VI2 ;
  RECT 1374.820 136.180 1375.020 136.380 ;
  LAYER VI2 ;
  RECT 1374.420 136.180 1374.620 136.380 ;
  LAYER VI3 ;
  RECT 1374.360 132.500 1375.220 132.780 ;
  LAYER VI3 ;
  RECT 1374.820 132.500 1375.020 132.700 ;
  LAYER VI3 ;
  RECT 1374.420 132.500 1374.620 132.700 ;
  LAYER VI2 ;
  RECT 1374.360 132.500 1375.220 132.780 ;
  LAYER VI2 ;
  RECT 1374.820 132.500 1375.020 132.700 ;
  LAYER VI2 ;
  RECT 1374.420 132.500 1374.620 132.700 ;
  LAYER VI3 ;
  RECT 1374.360 128.820 1375.220 129.100 ;
  LAYER VI3 ;
  RECT 1374.820 128.820 1375.020 129.020 ;
  LAYER VI3 ;
  RECT 1374.420 128.820 1374.620 129.020 ;
  LAYER VI2 ;
  RECT 1374.360 128.820 1375.220 129.100 ;
  LAYER VI2 ;
  RECT 1374.820 128.820 1375.020 129.020 ;
  LAYER VI2 ;
  RECT 1374.420 128.820 1374.620 129.020 ;
  LAYER VI3 ;
  RECT 1374.360 125.140 1375.220 125.420 ;
  LAYER VI3 ;
  RECT 1374.820 125.140 1375.020 125.340 ;
  LAYER VI3 ;
  RECT 1374.420 125.140 1374.620 125.340 ;
  LAYER VI2 ;
  RECT 1374.360 125.140 1375.220 125.420 ;
  LAYER VI2 ;
  RECT 1374.820 125.140 1375.020 125.340 ;
  LAYER VI2 ;
  RECT 1374.420 125.140 1374.620 125.340 ;
  LAYER VI3 ;
  RECT 1374.360 121.460 1375.220 121.740 ;
  LAYER VI3 ;
  RECT 1374.820 121.460 1375.020 121.660 ;
  LAYER VI3 ;
  RECT 1374.420 121.460 1374.620 121.660 ;
  LAYER VI2 ;
  RECT 1374.360 121.460 1375.220 121.740 ;
  LAYER VI2 ;
  RECT 1374.820 121.460 1375.020 121.660 ;
  LAYER VI2 ;
  RECT 1374.420 121.460 1374.620 121.660 ;
  LAYER VI3 ;
  RECT 1374.360 117.780 1375.220 118.060 ;
  LAYER VI3 ;
  RECT 1374.820 117.780 1375.020 117.980 ;
  LAYER VI3 ;
  RECT 1374.420 117.780 1374.620 117.980 ;
  LAYER VI2 ;
  RECT 1374.360 117.780 1375.220 118.060 ;
  LAYER VI2 ;
  RECT 1374.820 117.780 1375.020 117.980 ;
  LAYER VI2 ;
  RECT 1374.420 117.780 1374.620 117.980 ;
  LAYER VI3 ;
  RECT 1374.360 114.100 1375.220 114.380 ;
  LAYER VI3 ;
  RECT 1374.820 114.100 1375.020 114.300 ;
  LAYER VI3 ;
  RECT 1374.420 114.100 1374.620 114.300 ;
  LAYER VI2 ;
  RECT 1374.360 114.100 1375.220 114.380 ;
  LAYER VI2 ;
  RECT 1374.820 114.100 1375.020 114.300 ;
  LAYER VI2 ;
  RECT 1374.420 114.100 1374.620 114.300 ;
  LAYER VI3 ;
  RECT 1374.360 110.420 1375.220 110.700 ;
  LAYER VI3 ;
  RECT 1374.820 110.420 1375.020 110.620 ;
  LAYER VI3 ;
  RECT 1374.420 110.420 1374.620 110.620 ;
  LAYER VI2 ;
  RECT 1374.360 110.420 1375.220 110.700 ;
  LAYER VI2 ;
  RECT 1374.820 110.420 1375.020 110.620 ;
  LAYER VI2 ;
  RECT 1374.420 110.420 1374.620 110.620 ;
  LAYER VI3 ;
  RECT 1374.360 106.740 1375.220 107.020 ;
  LAYER VI3 ;
  RECT 1374.820 106.740 1375.020 106.940 ;
  LAYER VI3 ;
  RECT 1374.420 106.740 1374.620 106.940 ;
  LAYER VI2 ;
  RECT 1374.360 106.740 1375.220 107.020 ;
  LAYER VI2 ;
  RECT 1374.820 106.740 1375.020 106.940 ;
  LAYER VI2 ;
  RECT 1374.420 106.740 1374.620 106.940 ;
  LAYER VI3 ;
  RECT 1374.360 103.060 1375.220 103.340 ;
  LAYER VI3 ;
  RECT 1374.820 103.060 1375.020 103.260 ;
  LAYER VI3 ;
  RECT 1374.420 103.060 1374.620 103.260 ;
  LAYER VI2 ;
  RECT 1374.360 103.060 1375.220 103.340 ;
  LAYER VI2 ;
  RECT 1374.820 103.060 1375.020 103.260 ;
  LAYER VI2 ;
  RECT 1374.420 103.060 1374.620 103.260 ;
  LAYER VI3 ;
  RECT 1374.360 99.380 1375.220 99.660 ;
  LAYER VI3 ;
  RECT 1374.820 99.380 1375.020 99.580 ;
  LAYER VI3 ;
  RECT 1374.420 99.380 1374.620 99.580 ;
  LAYER VI2 ;
  RECT 1374.360 99.380 1375.220 99.660 ;
  LAYER VI2 ;
  RECT 1374.820 99.380 1375.020 99.580 ;
  LAYER VI2 ;
  RECT 1374.420 99.380 1374.620 99.580 ;
  LAYER VI3 ;
  RECT 1374.360 95.700 1375.220 95.980 ;
  LAYER VI3 ;
  RECT 1374.820 95.700 1375.020 95.900 ;
  LAYER VI3 ;
  RECT 1374.420 95.700 1374.620 95.900 ;
  LAYER VI2 ;
  RECT 1374.360 95.700 1375.220 95.980 ;
  LAYER VI2 ;
  RECT 1374.820 95.700 1375.020 95.900 ;
  LAYER VI2 ;
  RECT 1374.420 95.700 1374.620 95.900 ;
  LAYER VI3 ;
  RECT 1374.360 92.020 1375.220 92.300 ;
  LAYER VI3 ;
  RECT 1374.820 92.020 1375.020 92.220 ;
  LAYER VI3 ;
  RECT 1374.420 92.020 1374.620 92.220 ;
  LAYER VI2 ;
  RECT 1374.360 92.020 1375.220 92.300 ;
  LAYER VI2 ;
  RECT 1374.820 92.020 1375.020 92.220 ;
  LAYER VI2 ;
  RECT 1374.420 92.020 1374.620 92.220 ;
  LAYER VI3 ;
  RECT 1374.360 88.340 1375.220 88.620 ;
  LAYER VI3 ;
  RECT 1374.820 88.340 1375.020 88.540 ;
  LAYER VI3 ;
  RECT 1374.420 88.340 1374.620 88.540 ;
  LAYER VI2 ;
  RECT 1374.360 88.340 1375.220 88.620 ;
  LAYER VI2 ;
  RECT 1374.820 88.340 1375.020 88.540 ;
  LAYER VI2 ;
  RECT 1374.420 88.340 1374.620 88.540 ;
  LAYER VI3 ;
  RECT 1374.360 84.660 1375.220 84.940 ;
  LAYER VI3 ;
  RECT 1374.820 84.660 1375.020 84.860 ;
  LAYER VI3 ;
  RECT 1374.420 84.660 1374.620 84.860 ;
  LAYER VI2 ;
  RECT 1374.360 84.660 1375.220 84.940 ;
  LAYER VI2 ;
  RECT 1374.820 84.660 1375.020 84.860 ;
  LAYER VI2 ;
  RECT 1374.420 84.660 1374.620 84.860 ;
  LAYER VI3 ;
  RECT 1374.360 80.980 1375.220 81.260 ;
  LAYER VI3 ;
  RECT 1374.820 80.980 1375.020 81.180 ;
  LAYER VI3 ;
  RECT 1374.420 80.980 1374.620 81.180 ;
  LAYER VI2 ;
  RECT 1374.360 80.980 1375.220 81.260 ;
  LAYER VI2 ;
  RECT 1374.820 80.980 1375.020 81.180 ;
  LAYER VI2 ;
  RECT 1374.420 80.980 1374.620 81.180 ;
  LAYER VI3 ;
  RECT 1374.360 77.300 1375.220 77.580 ;
  LAYER VI3 ;
  RECT 1374.820 77.300 1375.020 77.500 ;
  LAYER VI3 ;
  RECT 1374.420 77.300 1374.620 77.500 ;
  LAYER VI2 ;
  RECT 1374.360 77.300 1375.220 77.580 ;
  LAYER VI2 ;
  RECT 1374.820 77.300 1375.020 77.500 ;
  LAYER VI2 ;
  RECT 1374.420 77.300 1374.620 77.500 ;
  LAYER VI3 ;
  RECT 1374.360 73.620 1375.220 73.900 ;
  LAYER VI3 ;
  RECT 1374.820 73.620 1375.020 73.820 ;
  LAYER VI3 ;
  RECT 1374.420 73.620 1374.620 73.820 ;
  LAYER VI2 ;
  RECT 1374.360 73.620 1375.220 73.900 ;
  LAYER VI2 ;
  RECT 1374.820 73.620 1375.020 73.820 ;
  LAYER VI2 ;
  RECT 1374.420 73.620 1374.620 73.820 ;
  LAYER VI3 ;
  RECT 1374.360 69.940 1375.220 70.220 ;
  LAYER VI3 ;
  RECT 1374.820 69.940 1375.020 70.140 ;
  LAYER VI3 ;
  RECT 1374.420 69.940 1374.620 70.140 ;
  LAYER VI2 ;
  RECT 1374.360 69.940 1375.220 70.220 ;
  LAYER VI2 ;
  RECT 1374.820 69.940 1375.020 70.140 ;
  LAYER VI2 ;
  RECT 1374.420 69.940 1374.620 70.140 ;
  LAYER VI3 ;
  RECT 1374.360 65.600 1375.220 65.980 ;
  LAYER VI3 ;
  RECT 1374.760 65.660 1374.960 65.860 ;
  LAYER VI3 ;
  RECT 1374.360 65.660 1374.560 65.860 ;
  LAYER VI2 ;
  RECT 1374.360 65.600 1375.220 65.980 ;
  LAYER VI2 ;
  RECT 1374.760 65.660 1374.960 65.860 ;
  LAYER VI2 ;
  RECT 1374.360 65.660 1374.560 65.860 ;
  LAYER VI3 ;
  RECT 718.100 546.070 718.350 546.930 ;
  LAYER VI3 ;
  RECT 718.100 546.530 718.300 546.730 ;
  LAYER VI3 ;
  RECT 718.100 546.130 718.300 546.330 ;
  LAYER VI2 ;
  RECT 718.100 546.070 718.350 546.930 ;
  LAYER VI2 ;
  RECT 718.100 546.530 718.300 546.730 ;
  LAYER VI2 ;
  RECT 718.100 546.130 718.300 546.330 ;
  LAYER VI3 ;
  RECT 759.020 546.070 759.270 546.930 ;
  LAYER VI3 ;
  RECT 759.020 546.530 759.220 546.730 ;
  LAYER VI3 ;
  RECT 759.020 546.130 759.220 546.330 ;
  LAYER VI2 ;
  RECT 759.020 546.070 759.270 546.930 ;
  LAYER VI2 ;
  RECT 759.020 546.530 759.220 546.730 ;
  LAYER VI2 ;
  RECT 759.020 546.130 759.220 546.330 ;
  LAYER VI3 ;
  RECT 799.940 546.070 800.190 546.930 ;
  LAYER VI3 ;
  RECT 799.940 546.530 800.140 546.730 ;
  LAYER VI3 ;
  RECT 799.940 546.130 800.140 546.330 ;
  LAYER VI2 ;
  RECT 799.940 546.070 800.190 546.930 ;
  LAYER VI2 ;
  RECT 799.940 546.530 800.140 546.730 ;
  LAYER VI2 ;
  RECT 799.940 546.130 800.140 546.330 ;
  LAYER VI3 ;
  RECT 840.860 546.070 841.110 546.930 ;
  LAYER VI3 ;
  RECT 840.860 546.530 841.060 546.730 ;
  LAYER VI3 ;
  RECT 840.860 546.130 841.060 546.330 ;
  LAYER VI2 ;
  RECT 840.860 546.070 841.110 546.930 ;
  LAYER VI2 ;
  RECT 840.860 546.530 841.060 546.730 ;
  LAYER VI2 ;
  RECT 840.860 546.130 841.060 546.330 ;
  LAYER VI3 ;
  RECT 881.780 546.070 882.030 546.930 ;
  LAYER VI3 ;
  RECT 881.780 546.530 881.980 546.730 ;
  LAYER VI3 ;
  RECT 881.780 546.130 881.980 546.330 ;
  LAYER VI2 ;
  RECT 881.780 546.070 882.030 546.930 ;
  LAYER VI2 ;
  RECT 881.780 546.530 881.980 546.730 ;
  LAYER VI2 ;
  RECT 881.780 546.130 881.980 546.330 ;
  LAYER VI3 ;
  RECT 922.700 546.070 922.950 546.930 ;
  LAYER VI3 ;
  RECT 922.700 546.530 922.900 546.730 ;
  LAYER VI3 ;
  RECT 922.700 546.130 922.900 546.330 ;
  LAYER VI2 ;
  RECT 922.700 546.070 922.950 546.930 ;
  LAYER VI2 ;
  RECT 922.700 546.530 922.900 546.730 ;
  LAYER VI2 ;
  RECT 922.700 546.130 922.900 546.330 ;
  LAYER VI3 ;
  RECT 963.620 546.070 963.870 546.930 ;
  LAYER VI3 ;
  RECT 963.620 546.530 963.820 546.730 ;
  LAYER VI3 ;
  RECT 963.620 546.130 963.820 546.330 ;
  LAYER VI2 ;
  RECT 963.620 546.070 963.870 546.930 ;
  LAYER VI2 ;
  RECT 963.620 546.530 963.820 546.730 ;
  LAYER VI2 ;
  RECT 963.620 546.130 963.820 546.330 ;
  LAYER VI3 ;
  RECT 1004.540 546.070 1004.790 546.930 ;
  LAYER VI3 ;
  RECT 1004.540 546.530 1004.740 546.730 ;
  LAYER VI3 ;
  RECT 1004.540 546.130 1004.740 546.330 ;
  LAYER VI2 ;
  RECT 1004.540 546.070 1004.790 546.930 ;
  LAYER VI2 ;
  RECT 1004.540 546.530 1004.740 546.730 ;
  LAYER VI2 ;
  RECT 1004.540 546.130 1004.740 546.330 ;
  LAYER VI3 ;
  RECT 1045.460 546.070 1045.710 546.930 ;
  LAYER VI3 ;
  RECT 1045.460 546.530 1045.660 546.730 ;
  LAYER VI3 ;
  RECT 1045.460 546.130 1045.660 546.330 ;
  LAYER VI2 ;
  RECT 1045.460 546.070 1045.710 546.930 ;
  LAYER VI2 ;
  RECT 1045.460 546.530 1045.660 546.730 ;
  LAYER VI2 ;
  RECT 1045.460 546.130 1045.660 546.330 ;
  LAYER VI3 ;
  RECT 1086.380 546.070 1086.630 546.930 ;
  LAYER VI3 ;
  RECT 1086.380 546.530 1086.580 546.730 ;
  LAYER VI3 ;
  RECT 1086.380 546.130 1086.580 546.330 ;
  LAYER VI2 ;
  RECT 1086.380 546.070 1086.630 546.930 ;
  LAYER VI2 ;
  RECT 1086.380 546.530 1086.580 546.730 ;
  LAYER VI2 ;
  RECT 1086.380 546.130 1086.580 546.330 ;
  LAYER VI3 ;
  RECT 1127.300 546.070 1127.550 546.930 ;
  LAYER VI3 ;
  RECT 1127.300 546.530 1127.500 546.730 ;
  LAYER VI3 ;
  RECT 1127.300 546.130 1127.500 546.330 ;
  LAYER VI2 ;
  RECT 1127.300 546.070 1127.550 546.930 ;
  LAYER VI2 ;
  RECT 1127.300 546.530 1127.500 546.730 ;
  LAYER VI2 ;
  RECT 1127.300 546.130 1127.500 546.330 ;
  LAYER VI3 ;
  RECT 1168.220 546.070 1168.470 546.930 ;
  LAYER VI3 ;
  RECT 1168.220 546.530 1168.420 546.730 ;
  LAYER VI3 ;
  RECT 1168.220 546.130 1168.420 546.330 ;
  LAYER VI2 ;
  RECT 1168.220 546.070 1168.470 546.930 ;
  LAYER VI2 ;
  RECT 1168.220 546.530 1168.420 546.730 ;
  LAYER VI2 ;
  RECT 1168.220 546.130 1168.420 546.330 ;
  LAYER VI3 ;
  RECT 1209.140 546.070 1209.390 546.930 ;
  LAYER VI3 ;
  RECT 1209.140 546.530 1209.340 546.730 ;
  LAYER VI3 ;
  RECT 1209.140 546.130 1209.340 546.330 ;
  LAYER VI2 ;
  RECT 1209.140 546.070 1209.390 546.930 ;
  LAYER VI2 ;
  RECT 1209.140 546.530 1209.340 546.730 ;
  LAYER VI2 ;
  RECT 1209.140 546.130 1209.340 546.330 ;
  LAYER VI3 ;
  RECT 1250.060 546.070 1250.310 546.930 ;
  LAYER VI3 ;
  RECT 1250.060 546.530 1250.260 546.730 ;
  LAYER VI3 ;
  RECT 1250.060 546.130 1250.260 546.330 ;
  LAYER VI2 ;
  RECT 1250.060 546.070 1250.310 546.930 ;
  LAYER VI2 ;
  RECT 1250.060 546.530 1250.260 546.730 ;
  LAYER VI2 ;
  RECT 1250.060 546.130 1250.260 546.330 ;
  LAYER VI3 ;
  RECT 1290.980 546.070 1291.230 546.930 ;
  LAYER VI3 ;
  RECT 1290.980 546.530 1291.180 546.730 ;
  LAYER VI3 ;
  RECT 1290.980 546.130 1291.180 546.330 ;
  LAYER VI2 ;
  RECT 1290.980 546.070 1291.230 546.930 ;
  LAYER VI2 ;
  RECT 1290.980 546.530 1291.180 546.730 ;
  LAYER VI2 ;
  RECT 1290.980 546.130 1291.180 546.330 ;
  LAYER VI3 ;
  RECT 1331.900 546.070 1332.150 546.930 ;
  LAYER VI3 ;
  RECT 1331.900 546.530 1332.100 546.730 ;
  LAYER VI3 ;
  RECT 1331.900 546.130 1332.100 546.330 ;
  LAYER VI2 ;
  RECT 1331.900 546.070 1332.150 546.930 ;
  LAYER VI2 ;
  RECT 1331.900 546.530 1332.100 546.730 ;
  LAYER VI2 ;
  RECT 1331.900 546.130 1332.100 546.330 ;
  LAYER VI3 ;
  RECT 701.090 546.070 703.600 546.930 ;
  LAYER VI3 ;
  RECT 703.090 546.530 703.290 546.730 ;
  LAYER VI3 ;
  RECT 703.090 546.130 703.290 546.330 ;
  LAYER VI3 ;
  RECT 702.690 546.530 702.890 546.730 ;
  LAYER VI3 ;
  RECT 702.690 546.130 702.890 546.330 ;
  LAYER VI3 ;
  RECT 702.290 546.530 702.490 546.730 ;
  LAYER VI3 ;
  RECT 702.290 546.130 702.490 546.330 ;
  LAYER VI3 ;
  RECT 701.890 546.530 702.090 546.730 ;
  LAYER VI3 ;
  RECT 701.890 546.130 702.090 546.330 ;
  LAYER VI3 ;
  RECT 701.490 546.530 701.690 546.730 ;
  LAYER VI3 ;
  RECT 701.490 546.130 701.690 546.330 ;
  LAYER VI3 ;
  RECT 701.090 546.530 701.290 546.730 ;
  LAYER VI3 ;
  RECT 701.090 546.130 701.290 546.330 ;
  LAYER VI2 ;
  RECT 701.090 546.070 703.600 546.930 ;
  LAYER VI2 ;
  RECT 703.090 546.530 703.290 546.730 ;
  LAYER VI2 ;
  RECT 703.090 546.130 703.290 546.330 ;
  LAYER VI2 ;
  RECT 702.690 546.530 702.890 546.730 ;
  LAYER VI2 ;
  RECT 702.690 546.130 702.890 546.330 ;
  LAYER VI2 ;
  RECT 702.290 546.530 702.490 546.730 ;
  LAYER VI2 ;
  RECT 702.290 546.130 702.490 546.330 ;
  LAYER VI2 ;
  RECT 701.890 546.530 702.090 546.730 ;
  LAYER VI2 ;
  RECT 701.890 546.130 702.090 546.330 ;
  LAYER VI2 ;
  RECT 701.490 546.530 701.690 546.730 ;
  LAYER VI2 ;
  RECT 701.490 546.130 701.690 546.330 ;
  LAYER VI2 ;
  RECT 701.090 546.530 701.290 546.730 ;
  LAYER VI2 ;
  RECT 701.090 546.130 701.290 546.330 ;
  LAYER VI3 ;
  RECT 688.670 546.070 691.060 546.930 ;
  LAYER VI3 ;
  RECT 690.670 546.530 690.870 546.730 ;
  LAYER VI3 ;
  RECT 690.670 546.130 690.870 546.330 ;
  LAYER VI3 ;
  RECT 690.270 546.530 690.470 546.730 ;
  LAYER VI3 ;
  RECT 690.270 546.130 690.470 546.330 ;
  LAYER VI3 ;
  RECT 689.870 546.530 690.070 546.730 ;
  LAYER VI3 ;
  RECT 689.870 546.130 690.070 546.330 ;
  LAYER VI3 ;
  RECT 689.470 546.530 689.670 546.730 ;
  LAYER VI3 ;
  RECT 689.470 546.130 689.670 546.330 ;
  LAYER VI3 ;
  RECT 689.070 546.530 689.270 546.730 ;
  LAYER VI3 ;
  RECT 689.070 546.130 689.270 546.330 ;
  LAYER VI3 ;
  RECT 688.670 546.530 688.870 546.730 ;
  LAYER VI3 ;
  RECT 688.670 546.130 688.870 546.330 ;
  LAYER VI2 ;
  RECT 688.670 546.070 691.060 546.930 ;
  LAYER VI2 ;
  RECT 690.670 546.530 690.870 546.730 ;
  LAYER VI2 ;
  RECT 690.670 546.130 690.870 546.330 ;
  LAYER VI2 ;
  RECT 690.270 546.530 690.470 546.730 ;
  LAYER VI2 ;
  RECT 690.270 546.130 690.470 546.330 ;
  LAYER VI2 ;
  RECT 689.870 546.530 690.070 546.730 ;
  LAYER VI2 ;
  RECT 689.870 546.130 690.070 546.330 ;
  LAYER VI2 ;
  RECT 689.470 546.530 689.670 546.730 ;
  LAYER VI2 ;
  RECT 689.470 546.130 689.670 546.330 ;
  LAYER VI2 ;
  RECT 689.070 546.530 689.270 546.730 ;
  LAYER VI2 ;
  RECT 689.070 546.130 689.270 546.330 ;
  LAYER VI2 ;
  RECT 688.670 546.530 688.870 546.730 ;
  LAYER VI2 ;
  RECT 688.670 546.130 688.870 546.330 ;
  LAYER VI3 ;
  RECT 681.160 546.070 684.220 546.930 ;
  LAYER VI3 ;
  RECT 683.960 546.530 684.160 546.730 ;
  LAYER VI3 ;
  RECT 683.960 546.130 684.160 546.330 ;
  LAYER VI3 ;
  RECT 683.560 546.530 683.760 546.730 ;
  LAYER VI3 ;
  RECT 683.560 546.130 683.760 546.330 ;
  LAYER VI3 ;
  RECT 683.160 546.530 683.360 546.730 ;
  LAYER VI3 ;
  RECT 683.160 546.130 683.360 546.330 ;
  LAYER VI3 ;
  RECT 682.760 546.530 682.960 546.730 ;
  LAYER VI3 ;
  RECT 682.760 546.130 682.960 546.330 ;
  LAYER VI3 ;
  RECT 682.360 546.530 682.560 546.730 ;
  LAYER VI3 ;
  RECT 682.360 546.130 682.560 546.330 ;
  LAYER VI3 ;
  RECT 681.960 546.530 682.160 546.730 ;
  LAYER VI3 ;
  RECT 681.960 546.130 682.160 546.330 ;
  LAYER VI3 ;
  RECT 681.560 546.530 681.760 546.730 ;
  LAYER VI3 ;
  RECT 681.560 546.130 681.760 546.330 ;
  LAYER VI3 ;
  RECT 681.160 546.530 681.360 546.730 ;
  LAYER VI3 ;
  RECT 681.160 546.130 681.360 546.330 ;
  LAYER VI2 ;
  RECT 681.160 546.070 684.220 546.930 ;
  LAYER VI2 ;
  RECT 683.960 546.530 684.160 546.730 ;
  LAYER VI2 ;
  RECT 683.960 546.130 684.160 546.330 ;
  LAYER VI2 ;
  RECT 683.560 546.530 683.760 546.730 ;
  LAYER VI2 ;
  RECT 683.560 546.130 683.760 546.330 ;
  LAYER VI2 ;
  RECT 683.160 546.530 683.360 546.730 ;
  LAYER VI2 ;
  RECT 683.160 546.130 683.360 546.330 ;
  LAYER VI2 ;
  RECT 682.760 546.530 682.960 546.730 ;
  LAYER VI2 ;
  RECT 682.760 546.130 682.960 546.330 ;
  LAYER VI2 ;
  RECT 682.360 546.530 682.560 546.730 ;
  LAYER VI2 ;
  RECT 682.360 546.130 682.560 546.330 ;
  LAYER VI2 ;
  RECT 681.960 546.530 682.160 546.730 ;
  LAYER VI2 ;
  RECT 681.960 546.130 682.160 546.330 ;
  LAYER VI2 ;
  RECT 681.560 546.530 681.760 546.730 ;
  LAYER VI2 ;
  RECT 681.560 546.130 681.760 546.330 ;
  LAYER VI2 ;
  RECT 681.160 546.530 681.360 546.730 ;
  LAYER VI2 ;
  RECT 681.160 546.130 681.360 546.330 ;
  LAYER VI3 ;
  RECT 705.340 546.070 708.190 546.930 ;
  LAYER VI3 ;
  RECT 707.740 546.530 707.940 546.730 ;
  LAYER VI3 ;
  RECT 707.740 546.130 707.940 546.330 ;
  LAYER VI3 ;
  RECT 707.340 546.530 707.540 546.730 ;
  LAYER VI3 ;
  RECT 707.340 546.130 707.540 546.330 ;
  LAYER VI3 ;
  RECT 706.940 546.530 707.140 546.730 ;
  LAYER VI3 ;
  RECT 706.940 546.130 707.140 546.330 ;
  LAYER VI3 ;
  RECT 706.540 546.530 706.740 546.730 ;
  LAYER VI3 ;
  RECT 706.540 546.130 706.740 546.330 ;
  LAYER VI3 ;
  RECT 706.140 546.530 706.340 546.730 ;
  LAYER VI3 ;
  RECT 706.140 546.130 706.340 546.330 ;
  LAYER VI3 ;
  RECT 705.740 546.530 705.940 546.730 ;
  LAYER VI3 ;
  RECT 705.740 546.130 705.940 546.330 ;
  LAYER VI3 ;
  RECT 705.340 546.530 705.540 546.730 ;
  LAYER VI3 ;
  RECT 705.340 546.130 705.540 546.330 ;
  LAYER VI2 ;
  RECT 705.340 546.070 708.190 546.930 ;
  LAYER VI2 ;
  RECT 707.740 546.530 707.940 546.730 ;
  LAYER VI2 ;
  RECT 707.740 546.130 707.940 546.330 ;
  LAYER VI2 ;
  RECT 707.340 546.530 707.540 546.730 ;
  LAYER VI2 ;
  RECT 707.340 546.130 707.540 546.330 ;
  LAYER VI2 ;
  RECT 706.940 546.530 707.140 546.730 ;
  LAYER VI2 ;
  RECT 706.940 546.130 707.140 546.330 ;
  LAYER VI2 ;
  RECT 706.540 546.530 706.740 546.730 ;
  LAYER VI2 ;
  RECT 706.540 546.130 706.740 546.330 ;
  LAYER VI2 ;
  RECT 706.140 546.530 706.340 546.730 ;
  LAYER VI2 ;
  RECT 706.140 546.130 706.340 546.330 ;
  LAYER VI2 ;
  RECT 705.740 546.530 705.940 546.730 ;
  LAYER VI2 ;
  RECT 705.740 546.130 705.940 546.330 ;
  LAYER VI2 ;
  RECT 705.340 546.530 705.540 546.730 ;
  LAYER VI2 ;
  RECT 705.340 546.130 705.540 546.330 ;
  LAYER VI3 ;
  RECT 709.640 546.070 712.890 546.930 ;
  LAYER VI3 ;
  RECT 712.440 546.530 712.640 546.730 ;
  LAYER VI3 ;
  RECT 712.440 546.130 712.640 546.330 ;
  LAYER VI3 ;
  RECT 712.040 546.530 712.240 546.730 ;
  LAYER VI3 ;
  RECT 712.040 546.130 712.240 546.330 ;
  LAYER VI3 ;
  RECT 711.640 546.530 711.840 546.730 ;
  LAYER VI3 ;
  RECT 711.640 546.130 711.840 546.330 ;
  LAYER VI3 ;
  RECT 711.240 546.530 711.440 546.730 ;
  LAYER VI3 ;
  RECT 711.240 546.130 711.440 546.330 ;
  LAYER VI3 ;
  RECT 710.840 546.530 711.040 546.730 ;
  LAYER VI3 ;
  RECT 710.840 546.130 711.040 546.330 ;
  LAYER VI3 ;
  RECT 710.440 546.530 710.640 546.730 ;
  LAYER VI3 ;
  RECT 710.440 546.130 710.640 546.330 ;
  LAYER VI3 ;
  RECT 710.040 546.530 710.240 546.730 ;
  LAYER VI3 ;
  RECT 710.040 546.130 710.240 546.330 ;
  LAYER VI3 ;
  RECT 709.640 546.530 709.840 546.730 ;
  LAYER VI3 ;
  RECT 709.640 546.130 709.840 546.330 ;
  LAYER VI2 ;
  RECT 709.640 546.070 712.890 546.930 ;
  LAYER VI2 ;
  RECT 712.440 546.530 712.640 546.730 ;
  LAYER VI2 ;
  RECT 712.440 546.130 712.640 546.330 ;
  LAYER VI2 ;
  RECT 712.040 546.530 712.240 546.730 ;
  LAYER VI2 ;
  RECT 712.040 546.130 712.240 546.330 ;
  LAYER VI2 ;
  RECT 711.640 546.530 711.840 546.730 ;
  LAYER VI2 ;
  RECT 711.640 546.130 711.840 546.330 ;
  LAYER VI2 ;
  RECT 711.240 546.530 711.440 546.730 ;
  LAYER VI2 ;
  RECT 711.240 546.130 711.440 546.330 ;
  LAYER VI2 ;
  RECT 710.840 546.530 711.040 546.730 ;
  LAYER VI2 ;
  RECT 710.840 546.130 711.040 546.330 ;
  LAYER VI2 ;
  RECT 710.440 546.530 710.640 546.730 ;
  LAYER VI2 ;
  RECT 710.440 546.130 710.640 546.330 ;
  LAYER VI2 ;
  RECT 710.040 546.530 710.240 546.730 ;
  LAYER VI2 ;
  RECT 710.040 546.130 710.240 546.330 ;
  LAYER VI2 ;
  RECT 709.640 546.530 709.840 546.730 ;
  LAYER VI2 ;
  RECT 709.640 546.130 709.840 546.330 ;
  LAYER VI3 ;
  RECT 678.440 546.070 680.200 546.930 ;
  LAYER VI3 ;
  RECT 679.640 546.530 679.840 546.730 ;
  LAYER VI3 ;
  RECT 679.640 546.130 679.840 546.330 ;
  LAYER VI3 ;
  RECT 679.240 546.530 679.440 546.730 ;
  LAYER VI3 ;
  RECT 679.240 546.130 679.440 546.330 ;
  LAYER VI3 ;
  RECT 678.840 546.530 679.040 546.730 ;
  LAYER VI3 ;
  RECT 678.840 546.130 679.040 546.330 ;
  LAYER VI3 ;
  RECT 678.440 546.530 678.640 546.730 ;
  LAYER VI3 ;
  RECT 678.440 546.130 678.640 546.330 ;
  LAYER VI2 ;
  RECT 678.440 546.070 680.200 546.930 ;
  LAYER VI2 ;
  RECT 679.640 546.530 679.840 546.730 ;
  LAYER VI2 ;
  RECT 679.640 546.130 679.840 546.330 ;
  LAYER VI2 ;
  RECT 679.240 546.530 679.440 546.730 ;
  LAYER VI2 ;
  RECT 679.240 546.130 679.440 546.330 ;
  LAYER VI2 ;
  RECT 678.840 546.530 679.040 546.730 ;
  LAYER VI2 ;
  RECT 678.840 546.130 679.040 546.330 ;
  LAYER VI2 ;
  RECT 678.440 546.530 678.640 546.730 ;
  LAYER VI2 ;
  RECT 678.440 546.130 678.640 546.330 ;
  LAYER VI3 ;
  RECT 673.100 546.070 674.860 546.930 ;
  LAYER VI3 ;
  RECT 674.300 546.530 674.500 546.730 ;
  LAYER VI3 ;
  RECT 674.300 546.130 674.500 546.330 ;
  LAYER VI3 ;
  RECT 673.900 546.530 674.100 546.730 ;
  LAYER VI3 ;
  RECT 673.900 546.130 674.100 546.330 ;
  LAYER VI3 ;
  RECT 673.500 546.530 673.700 546.730 ;
  LAYER VI3 ;
  RECT 673.500 546.130 673.700 546.330 ;
  LAYER VI3 ;
  RECT 673.100 546.530 673.300 546.730 ;
  LAYER VI3 ;
  RECT 673.100 546.130 673.300 546.330 ;
  LAYER VI2 ;
  RECT 673.100 546.070 674.860 546.930 ;
  LAYER VI2 ;
  RECT 674.300 546.530 674.500 546.730 ;
  LAYER VI2 ;
  RECT 674.300 546.130 674.500 546.330 ;
  LAYER VI2 ;
  RECT 673.900 546.530 674.100 546.730 ;
  LAYER VI2 ;
  RECT 673.900 546.130 674.100 546.330 ;
  LAYER VI2 ;
  RECT 673.500 546.530 673.700 546.730 ;
  LAYER VI2 ;
  RECT 673.500 546.130 673.700 546.330 ;
  LAYER VI2 ;
  RECT 673.100 546.530 673.300 546.730 ;
  LAYER VI2 ;
  RECT 673.100 546.130 673.300 546.330 ;
  LAYER VI3 ;
  RECT 669.100 546.070 670.860 546.930 ;
  LAYER VI3 ;
  RECT 670.300 546.530 670.500 546.730 ;
  LAYER VI3 ;
  RECT 670.300 546.130 670.500 546.330 ;
  LAYER VI3 ;
  RECT 669.900 546.530 670.100 546.730 ;
  LAYER VI3 ;
  RECT 669.900 546.130 670.100 546.330 ;
  LAYER VI3 ;
  RECT 669.500 546.530 669.700 546.730 ;
  LAYER VI3 ;
  RECT 669.500 546.130 669.700 546.330 ;
  LAYER VI3 ;
  RECT 669.100 546.530 669.300 546.730 ;
  LAYER VI3 ;
  RECT 669.100 546.130 669.300 546.330 ;
  LAYER VI2 ;
  RECT 669.100 546.070 670.860 546.930 ;
  LAYER VI2 ;
  RECT 670.300 546.530 670.500 546.730 ;
  LAYER VI2 ;
  RECT 670.300 546.130 670.500 546.330 ;
  LAYER VI2 ;
  RECT 669.900 546.530 670.100 546.730 ;
  LAYER VI2 ;
  RECT 669.900 546.130 670.100 546.330 ;
  LAYER VI2 ;
  RECT 669.500 546.530 669.700 546.730 ;
  LAYER VI2 ;
  RECT 669.500 546.130 669.700 546.330 ;
  LAYER VI2 ;
  RECT 669.100 546.530 669.300 546.730 ;
  LAYER VI2 ;
  RECT 669.100 546.130 669.300 546.330 ;
  LAYER VI3 ;
  RECT 665.100 546.070 666.860 546.930 ;
  LAYER VI3 ;
  RECT 666.300 546.530 666.500 546.730 ;
  LAYER VI3 ;
  RECT 666.300 546.130 666.500 546.330 ;
  LAYER VI3 ;
  RECT 665.900 546.530 666.100 546.730 ;
  LAYER VI3 ;
  RECT 665.900 546.130 666.100 546.330 ;
  LAYER VI3 ;
  RECT 665.500 546.530 665.700 546.730 ;
  LAYER VI3 ;
  RECT 665.500 546.130 665.700 546.330 ;
  LAYER VI3 ;
  RECT 665.100 546.530 665.300 546.730 ;
  LAYER VI3 ;
  RECT 665.100 546.130 665.300 546.330 ;
  LAYER VI2 ;
  RECT 665.100 546.070 666.860 546.930 ;
  LAYER VI2 ;
  RECT 666.300 546.530 666.500 546.730 ;
  LAYER VI2 ;
  RECT 666.300 546.130 666.500 546.330 ;
  LAYER VI2 ;
  RECT 665.900 546.530 666.100 546.730 ;
  LAYER VI2 ;
  RECT 665.900 546.130 666.100 546.330 ;
  LAYER VI2 ;
  RECT 665.500 546.530 665.700 546.730 ;
  LAYER VI2 ;
  RECT 665.500 546.130 665.700 546.330 ;
  LAYER VI2 ;
  RECT 665.100 546.530 665.300 546.730 ;
  LAYER VI2 ;
  RECT 665.100 546.130 665.300 546.330 ;
  LAYER VI3 ;
  RECT 4.280 65.600 5.140 65.980 ;
  LAYER VI3 ;
  RECT 4.680 65.660 4.880 65.860 ;
  LAYER VI3 ;
  RECT 4.280 65.660 4.480 65.860 ;
  LAYER VI2 ;
  RECT 4.280 65.600 5.140 65.980 ;
  LAYER VI2 ;
  RECT 4.680 65.660 4.880 65.860 ;
  LAYER VI2 ;
  RECT 4.280 65.660 4.480 65.860 ;
  LAYER VI3 ;
  RECT 4.280 69.940 5.140 70.220 ;
  LAYER VI3 ;
  RECT 4.740 69.940 4.940 70.140 ;
  LAYER VI3 ;
  RECT 4.340 69.940 4.540 70.140 ;
  LAYER VI2 ;
  RECT 4.280 69.940 5.140 70.220 ;
  LAYER VI2 ;
  RECT 4.740 69.940 4.940 70.140 ;
  LAYER VI2 ;
  RECT 4.340 69.940 4.540 70.140 ;
  LAYER VI3 ;
  RECT 4.280 73.620 5.140 73.900 ;
  LAYER VI3 ;
  RECT 4.740 73.620 4.940 73.820 ;
  LAYER VI3 ;
  RECT 4.340 73.620 4.540 73.820 ;
  LAYER VI2 ;
  RECT 4.280 73.620 5.140 73.900 ;
  LAYER VI2 ;
  RECT 4.740 73.620 4.940 73.820 ;
  LAYER VI2 ;
  RECT 4.340 73.620 4.540 73.820 ;
  LAYER VI3 ;
  RECT 4.280 77.300 5.140 77.580 ;
  LAYER VI3 ;
  RECT 4.740 77.300 4.940 77.500 ;
  LAYER VI3 ;
  RECT 4.340 77.300 4.540 77.500 ;
  LAYER VI2 ;
  RECT 4.280 77.300 5.140 77.580 ;
  LAYER VI2 ;
  RECT 4.740 77.300 4.940 77.500 ;
  LAYER VI2 ;
  RECT 4.340 77.300 4.540 77.500 ;
  LAYER VI3 ;
  RECT 4.280 80.980 5.140 81.260 ;
  LAYER VI3 ;
  RECT 4.740 80.980 4.940 81.180 ;
  LAYER VI3 ;
  RECT 4.340 80.980 4.540 81.180 ;
  LAYER VI2 ;
  RECT 4.280 80.980 5.140 81.260 ;
  LAYER VI2 ;
  RECT 4.740 80.980 4.940 81.180 ;
  LAYER VI2 ;
  RECT 4.340 80.980 4.540 81.180 ;
  LAYER VI3 ;
  RECT 4.280 84.660 5.140 84.940 ;
  LAYER VI3 ;
  RECT 4.740 84.660 4.940 84.860 ;
  LAYER VI3 ;
  RECT 4.340 84.660 4.540 84.860 ;
  LAYER VI2 ;
  RECT 4.280 84.660 5.140 84.940 ;
  LAYER VI2 ;
  RECT 4.740 84.660 4.940 84.860 ;
  LAYER VI2 ;
  RECT 4.340 84.660 4.540 84.860 ;
  LAYER VI3 ;
  RECT 4.280 88.340 5.140 88.620 ;
  LAYER VI3 ;
  RECT 4.740 88.340 4.940 88.540 ;
  LAYER VI3 ;
  RECT 4.340 88.340 4.540 88.540 ;
  LAYER VI2 ;
  RECT 4.280 88.340 5.140 88.620 ;
  LAYER VI2 ;
  RECT 4.740 88.340 4.940 88.540 ;
  LAYER VI2 ;
  RECT 4.340 88.340 4.540 88.540 ;
  LAYER VI3 ;
  RECT 4.280 92.020 5.140 92.300 ;
  LAYER VI3 ;
  RECT 4.740 92.020 4.940 92.220 ;
  LAYER VI3 ;
  RECT 4.340 92.020 4.540 92.220 ;
  LAYER VI2 ;
  RECT 4.280 92.020 5.140 92.300 ;
  LAYER VI2 ;
  RECT 4.740 92.020 4.940 92.220 ;
  LAYER VI2 ;
  RECT 4.340 92.020 4.540 92.220 ;
  LAYER VI3 ;
  RECT 4.280 95.700 5.140 95.980 ;
  LAYER VI3 ;
  RECT 4.740 95.700 4.940 95.900 ;
  LAYER VI3 ;
  RECT 4.340 95.700 4.540 95.900 ;
  LAYER VI2 ;
  RECT 4.280 95.700 5.140 95.980 ;
  LAYER VI2 ;
  RECT 4.740 95.700 4.940 95.900 ;
  LAYER VI2 ;
  RECT 4.340 95.700 4.540 95.900 ;
  LAYER VI3 ;
  RECT 4.280 99.380 5.140 99.660 ;
  LAYER VI3 ;
  RECT 4.740 99.380 4.940 99.580 ;
  LAYER VI3 ;
  RECT 4.340 99.380 4.540 99.580 ;
  LAYER VI2 ;
  RECT 4.280 99.380 5.140 99.660 ;
  LAYER VI2 ;
  RECT 4.740 99.380 4.940 99.580 ;
  LAYER VI2 ;
  RECT 4.340 99.380 4.540 99.580 ;
  LAYER VI3 ;
  RECT 4.280 103.060 5.140 103.340 ;
  LAYER VI3 ;
  RECT 4.740 103.060 4.940 103.260 ;
  LAYER VI3 ;
  RECT 4.340 103.060 4.540 103.260 ;
  LAYER VI2 ;
  RECT 4.280 103.060 5.140 103.340 ;
  LAYER VI2 ;
  RECT 4.740 103.060 4.940 103.260 ;
  LAYER VI2 ;
  RECT 4.340 103.060 4.540 103.260 ;
  LAYER VI3 ;
  RECT 4.280 106.740 5.140 107.020 ;
  LAYER VI3 ;
  RECT 4.740 106.740 4.940 106.940 ;
  LAYER VI3 ;
  RECT 4.340 106.740 4.540 106.940 ;
  LAYER VI2 ;
  RECT 4.280 106.740 5.140 107.020 ;
  LAYER VI2 ;
  RECT 4.740 106.740 4.940 106.940 ;
  LAYER VI2 ;
  RECT 4.340 106.740 4.540 106.940 ;
  LAYER VI3 ;
  RECT 4.280 110.420 5.140 110.700 ;
  LAYER VI3 ;
  RECT 4.740 110.420 4.940 110.620 ;
  LAYER VI3 ;
  RECT 4.340 110.420 4.540 110.620 ;
  LAYER VI2 ;
  RECT 4.280 110.420 5.140 110.700 ;
  LAYER VI2 ;
  RECT 4.740 110.420 4.940 110.620 ;
  LAYER VI2 ;
  RECT 4.340 110.420 4.540 110.620 ;
  LAYER VI3 ;
  RECT 4.280 114.100 5.140 114.380 ;
  LAYER VI3 ;
  RECT 4.740 114.100 4.940 114.300 ;
  LAYER VI3 ;
  RECT 4.340 114.100 4.540 114.300 ;
  LAYER VI2 ;
  RECT 4.280 114.100 5.140 114.380 ;
  LAYER VI2 ;
  RECT 4.740 114.100 4.940 114.300 ;
  LAYER VI2 ;
  RECT 4.340 114.100 4.540 114.300 ;
  LAYER VI3 ;
  RECT 4.280 117.780 5.140 118.060 ;
  LAYER VI3 ;
  RECT 4.740 117.780 4.940 117.980 ;
  LAYER VI3 ;
  RECT 4.340 117.780 4.540 117.980 ;
  LAYER VI2 ;
  RECT 4.280 117.780 5.140 118.060 ;
  LAYER VI2 ;
  RECT 4.740 117.780 4.940 117.980 ;
  LAYER VI2 ;
  RECT 4.340 117.780 4.540 117.980 ;
  LAYER VI3 ;
  RECT 4.280 121.460 5.140 121.740 ;
  LAYER VI3 ;
  RECT 4.740 121.460 4.940 121.660 ;
  LAYER VI3 ;
  RECT 4.340 121.460 4.540 121.660 ;
  LAYER VI2 ;
  RECT 4.280 121.460 5.140 121.740 ;
  LAYER VI2 ;
  RECT 4.740 121.460 4.940 121.660 ;
  LAYER VI2 ;
  RECT 4.340 121.460 4.540 121.660 ;
  LAYER VI3 ;
  RECT 4.280 125.140 5.140 125.420 ;
  LAYER VI3 ;
  RECT 4.740 125.140 4.940 125.340 ;
  LAYER VI3 ;
  RECT 4.340 125.140 4.540 125.340 ;
  LAYER VI2 ;
  RECT 4.280 125.140 5.140 125.420 ;
  LAYER VI2 ;
  RECT 4.740 125.140 4.940 125.340 ;
  LAYER VI2 ;
  RECT 4.340 125.140 4.540 125.340 ;
  LAYER VI3 ;
  RECT 4.280 128.820 5.140 129.100 ;
  LAYER VI3 ;
  RECT 4.740 128.820 4.940 129.020 ;
  LAYER VI3 ;
  RECT 4.340 128.820 4.540 129.020 ;
  LAYER VI2 ;
  RECT 4.280 128.820 5.140 129.100 ;
  LAYER VI2 ;
  RECT 4.740 128.820 4.940 129.020 ;
  LAYER VI2 ;
  RECT 4.340 128.820 4.540 129.020 ;
  LAYER VI3 ;
  RECT 4.280 132.500 5.140 132.780 ;
  LAYER VI3 ;
  RECT 4.740 132.500 4.940 132.700 ;
  LAYER VI3 ;
  RECT 4.340 132.500 4.540 132.700 ;
  LAYER VI2 ;
  RECT 4.280 132.500 5.140 132.780 ;
  LAYER VI2 ;
  RECT 4.740 132.500 4.940 132.700 ;
  LAYER VI2 ;
  RECT 4.340 132.500 4.540 132.700 ;
  LAYER VI3 ;
  RECT 4.280 136.180 5.140 136.460 ;
  LAYER VI3 ;
  RECT 4.740 136.180 4.940 136.380 ;
  LAYER VI3 ;
  RECT 4.340 136.180 4.540 136.380 ;
  LAYER VI2 ;
  RECT 4.280 136.180 5.140 136.460 ;
  LAYER VI2 ;
  RECT 4.740 136.180 4.940 136.380 ;
  LAYER VI2 ;
  RECT 4.340 136.180 4.540 136.380 ;
  LAYER VI3 ;
  RECT 4.280 139.860 5.140 140.140 ;
  LAYER VI3 ;
  RECT 4.740 139.860 4.940 140.060 ;
  LAYER VI3 ;
  RECT 4.340 139.860 4.540 140.060 ;
  LAYER VI2 ;
  RECT 4.280 139.860 5.140 140.140 ;
  LAYER VI2 ;
  RECT 4.740 139.860 4.940 140.060 ;
  LAYER VI2 ;
  RECT 4.340 139.860 4.540 140.060 ;
  LAYER VI3 ;
  RECT 4.280 143.540 5.140 143.820 ;
  LAYER VI3 ;
  RECT 4.740 143.540 4.940 143.740 ;
  LAYER VI3 ;
  RECT 4.340 143.540 4.540 143.740 ;
  LAYER VI2 ;
  RECT 4.280 143.540 5.140 143.820 ;
  LAYER VI2 ;
  RECT 4.740 143.540 4.940 143.740 ;
  LAYER VI2 ;
  RECT 4.340 143.540 4.540 143.740 ;
  LAYER VI3 ;
  RECT 4.280 147.220 5.140 147.500 ;
  LAYER VI3 ;
  RECT 4.740 147.220 4.940 147.420 ;
  LAYER VI3 ;
  RECT 4.340 147.220 4.540 147.420 ;
  LAYER VI2 ;
  RECT 4.280 147.220 5.140 147.500 ;
  LAYER VI2 ;
  RECT 4.740 147.220 4.940 147.420 ;
  LAYER VI2 ;
  RECT 4.340 147.220 4.540 147.420 ;
  LAYER VI3 ;
  RECT 4.280 150.900 5.140 151.180 ;
  LAYER VI3 ;
  RECT 4.740 150.900 4.940 151.100 ;
  LAYER VI3 ;
  RECT 4.340 150.900 4.540 151.100 ;
  LAYER VI2 ;
  RECT 4.280 150.900 5.140 151.180 ;
  LAYER VI2 ;
  RECT 4.740 150.900 4.940 151.100 ;
  LAYER VI2 ;
  RECT 4.340 150.900 4.540 151.100 ;
  LAYER VI3 ;
  RECT 4.280 154.580 5.140 154.860 ;
  LAYER VI3 ;
  RECT 4.740 154.580 4.940 154.780 ;
  LAYER VI3 ;
  RECT 4.340 154.580 4.540 154.780 ;
  LAYER VI2 ;
  RECT 4.280 154.580 5.140 154.860 ;
  LAYER VI2 ;
  RECT 4.740 154.580 4.940 154.780 ;
  LAYER VI2 ;
  RECT 4.340 154.580 4.540 154.780 ;
  LAYER VI3 ;
  RECT 4.280 158.260 5.140 158.540 ;
  LAYER VI3 ;
  RECT 4.740 158.260 4.940 158.460 ;
  LAYER VI3 ;
  RECT 4.340 158.260 4.540 158.460 ;
  LAYER VI2 ;
  RECT 4.280 158.260 5.140 158.540 ;
  LAYER VI2 ;
  RECT 4.740 158.260 4.940 158.460 ;
  LAYER VI2 ;
  RECT 4.340 158.260 4.540 158.460 ;
  LAYER VI3 ;
  RECT 4.280 161.940 5.140 162.220 ;
  LAYER VI3 ;
  RECT 4.740 161.940 4.940 162.140 ;
  LAYER VI3 ;
  RECT 4.340 161.940 4.540 162.140 ;
  LAYER VI2 ;
  RECT 4.280 161.940 5.140 162.220 ;
  LAYER VI2 ;
  RECT 4.740 161.940 4.940 162.140 ;
  LAYER VI2 ;
  RECT 4.340 161.940 4.540 162.140 ;
  LAYER VI3 ;
  RECT 4.280 165.620 5.140 165.900 ;
  LAYER VI3 ;
  RECT 4.740 165.620 4.940 165.820 ;
  LAYER VI3 ;
  RECT 4.340 165.620 4.540 165.820 ;
  LAYER VI2 ;
  RECT 4.280 165.620 5.140 165.900 ;
  LAYER VI2 ;
  RECT 4.740 165.620 4.940 165.820 ;
  LAYER VI2 ;
  RECT 4.340 165.620 4.540 165.820 ;
  LAYER VI3 ;
  RECT 4.280 169.300 5.140 169.580 ;
  LAYER VI3 ;
  RECT 4.740 169.300 4.940 169.500 ;
  LAYER VI3 ;
  RECT 4.340 169.300 4.540 169.500 ;
  LAYER VI2 ;
  RECT 4.280 169.300 5.140 169.580 ;
  LAYER VI2 ;
  RECT 4.740 169.300 4.940 169.500 ;
  LAYER VI2 ;
  RECT 4.340 169.300 4.540 169.500 ;
  LAYER VI3 ;
  RECT 4.280 172.980 5.140 173.260 ;
  LAYER VI3 ;
  RECT 4.740 172.980 4.940 173.180 ;
  LAYER VI3 ;
  RECT 4.340 172.980 4.540 173.180 ;
  LAYER VI2 ;
  RECT 4.280 172.980 5.140 173.260 ;
  LAYER VI2 ;
  RECT 4.740 172.980 4.940 173.180 ;
  LAYER VI2 ;
  RECT 4.340 172.980 4.540 173.180 ;
  LAYER VI3 ;
  RECT 4.280 176.660 5.140 176.940 ;
  LAYER VI3 ;
  RECT 4.740 176.660 4.940 176.860 ;
  LAYER VI3 ;
  RECT 4.340 176.660 4.540 176.860 ;
  LAYER VI2 ;
  RECT 4.280 176.660 5.140 176.940 ;
  LAYER VI2 ;
  RECT 4.740 176.660 4.940 176.860 ;
  LAYER VI2 ;
  RECT 4.340 176.660 4.540 176.860 ;
  LAYER VI3 ;
  RECT 4.280 180.340 5.140 180.620 ;
  LAYER VI3 ;
  RECT 4.740 180.340 4.940 180.540 ;
  LAYER VI3 ;
  RECT 4.340 180.340 4.540 180.540 ;
  LAYER VI2 ;
  RECT 4.280 180.340 5.140 180.620 ;
  LAYER VI2 ;
  RECT 4.740 180.340 4.940 180.540 ;
  LAYER VI2 ;
  RECT 4.340 180.340 4.540 180.540 ;
  LAYER VI3 ;
  RECT 4.280 184.020 5.140 184.300 ;
  LAYER VI3 ;
  RECT 4.740 184.020 4.940 184.220 ;
  LAYER VI3 ;
  RECT 4.340 184.020 4.540 184.220 ;
  LAYER VI2 ;
  RECT 4.280 184.020 5.140 184.300 ;
  LAYER VI2 ;
  RECT 4.740 184.020 4.940 184.220 ;
  LAYER VI2 ;
  RECT 4.340 184.020 4.540 184.220 ;
  LAYER VI3 ;
  RECT 4.280 187.700 5.140 187.980 ;
  LAYER VI3 ;
  RECT 4.740 187.700 4.940 187.900 ;
  LAYER VI3 ;
  RECT 4.340 187.700 4.540 187.900 ;
  LAYER VI2 ;
  RECT 4.280 187.700 5.140 187.980 ;
  LAYER VI2 ;
  RECT 4.740 187.700 4.940 187.900 ;
  LAYER VI2 ;
  RECT 4.340 187.700 4.540 187.900 ;
  LAYER VI3 ;
  RECT 4.280 191.380 5.140 191.660 ;
  LAYER VI3 ;
  RECT 4.740 191.380 4.940 191.580 ;
  LAYER VI3 ;
  RECT 4.340 191.380 4.540 191.580 ;
  LAYER VI2 ;
  RECT 4.280 191.380 5.140 191.660 ;
  LAYER VI2 ;
  RECT 4.740 191.380 4.940 191.580 ;
  LAYER VI2 ;
  RECT 4.340 191.380 4.540 191.580 ;
  LAYER VI3 ;
  RECT 4.280 195.060 5.140 195.340 ;
  LAYER VI3 ;
  RECT 4.740 195.060 4.940 195.260 ;
  LAYER VI3 ;
  RECT 4.340 195.060 4.540 195.260 ;
  LAYER VI2 ;
  RECT 4.280 195.060 5.140 195.340 ;
  LAYER VI2 ;
  RECT 4.740 195.060 4.940 195.260 ;
  LAYER VI2 ;
  RECT 4.340 195.060 4.540 195.260 ;
  LAYER VI3 ;
  RECT 4.280 198.740 5.140 199.020 ;
  LAYER VI3 ;
  RECT 4.740 198.740 4.940 198.940 ;
  LAYER VI3 ;
  RECT 4.340 198.740 4.540 198.940 ;
  LAYER VI2 ;
  RECT 4.280 198.740 5.140 199.020 ;
  LAYER VI2 ;
  RECT 4.740 198.740 4.940 198.940 ;
  LAYER VI2 ;
  RECT 4.340 198.740 4.540 198.940 ;
  LAYER VI3 ;
  RECT 4.280 202.420 5.140 202.700 ;
  LAYER VI3 ;
  RECT 4.740 202.420 4.940 202.620 ;
  LAYER VI3 ;
  RECT 4.340 202.420 4.540 202.620 ;
  LAYER VI2 ;
  RECT 4.280 202.420 5.140 202.700 ;
  LAYER VI2 ;
  RECT 4.740 202.420 4.940 202.620 ;
  LAYER VI2 ;
  RECT 4.340 202.420 4.540 202.620 ;
  LAYER VI3 ;
  RECT 4.280 206.100 5.140 206.380 ;
  LAYER VI3 ;
  RECT 4.740 206.100 4.940 206.300 ;
  LAYER VI3 ;
  RECT 4.340 206.100 4.540 206.300 ;
  LAYER VI2 ;
  RECT 4.280 206.100 5.140 206.380 ;
  LAYER VI2 ;
  RECT 4.740 206.100 4.940 206.300 ;
  LAYER VI2 ;
  RECT 4.340 206.100 4.540 206.300 ;
  LAYER VI3 ;
  RECT 4.280 209.780 5.140 210.060 ;
  LAYER VI3 ;
  RECT 4.740 209.780 4.940 209.980 ;
  LAYER VI3 ;
  RECT 4.340 209.780 4.540 209.980 ;
  LAYER VI2 ;
  RECT 4.280 209.780 5.140 210.060 ;
  LAYER VI2 ;
  RECT 4.740 209.780 4.940 209.980 ;
  LAYER VI2 ;
  RECT 4.340 209.780 4.540 209.980 ;
  LAYER VI3 ;
  RECT 4.280 213.460 5.140 213.740 ;
  LAYER VI3 ;
  RECT 4.740 213.460 4.940 213.660 ;
  LAYER VI3 ;
  RECT 4.340 213.460 4.540 213.660 ;
  LAYER VI2 ;
  RECT 4.280 213.460 5.140 213.740 ;
  LAYER VI2 ;
  RECT 4.740 213.460 4.940 213.660 ;
  LAYER VI2 ;
  RECT 4.340 213.460 4.540 213.660 ;
  LAYER VI3 ;
  RECT 4.280 217.140 5.140 217.420 ;
  LAYER VI3 ;
  RECT 4.740 217.140 4.940 217.340 ;
  LAYER VI3 ;
  RECT 4.340 217.140 4.540 217.340 ;
  LAYER VI2 ;
  RECT 4.280 217.140 5.140 217.420 ;
  LAYER VI2 ;
  RECT 4.740 217.140 4.940 217.340 ;
  LAYER VI2 ;
  RECT 4.340 217.140 4.540 217.340 ;
  LAYER VI3 ;
  RECT 4.280 220.820 5.140 221.100 ;
  LAYER VI3 ;
  RECT 4.740 220.820 4.940 221.020 ;
  LAYER VI3 ;
  RECT 4.340 220.820 4.540 221.020 ;
  LAYER VI2 ;
  RECT 4.280 220.820 5.140 221.100 ;
  LAYER VI2 ;
  RECT 4.740 220.820 4.940 221.020 ;
  LAYER VI2 ;
  RECT 4.340 220.820 4.540 221.020 ;
  LAYER VI3 ;
  RECT 4.280 224.500 5.140 224.780 ;
  LAYER VI3 ;
  RECT 4.740 224.500 4.940 224.700 ;
  LAYER VI3 ;
  RECT 4.340 224.500 4.540 224.700 ;
  LAYER VI2 ;
  RECT 4.280 224.500 5.140 224.780 ;
  LAYER VI2 ;
  RECT 4.740 224.500 4.940 224.700 ;
  LAYER VI2 ;
  RECT 4.340 224.500 4.540 224.700 ;
  LAYER VI3 ;
  RECT 4.280 228.180 5.140 228.460 ;
  LAYER VI3 ;
  RECT 4.740 228.180 4.940 228.380 ;
  LAYER VI3 ;
  RECT 4.340 228.180 4.540 228.380 ;
  LAYER VI2 ;
  RECT 4.280 228.180 5.140 228.460 ;
  LAYER VI2 ;
  RECT 4.740 228.180 4.940 228.380 ;
  LAYER VI2 ;
  RECT 4.340 228.180 4.540 228.380 ;
  LAYER VI3 ;
  RECT 4.280 231.860 5.140 232.140 ;
  LAYER VI3 ;
  RECT 4.740 231.860 4.940 232.060 ;
  LAYER VI3 ;
  RECT 4.340 231.860 4.540 232.060 ;
  LAYER VI2 ;
  RECT 4.280 231.860 5.140 232.140 ;
  LAYER VI2 ;
  RECT 4.740 231.860 4.940 232.060 ;
  LAYER VI2 ;
  RECT 4.340 231.860 4.540 232.060 ;
  LAYER VI3 ;
  RECT 4.280 235.540 5.140 235.820 ;
  LAYER VI3 ;
  RECT 4.740 235.540 4.940 235.740 ;
  LAYER VI3 ;
  RECT 4.340 235.540 4.540 235.740 ;
  LAYER VI2 ;
  RECT 4.280 235.540 5.140 235.820 ;
  LAYER VI2 ;
  RECT 4.740 235.540 4.940 235.740 ;
  LAYER VI2 ;
  RECT 4.340 235.540 4.540 235.740 ;
  LAYER VI3 ;
  RECT 4.280 239.220 5.140 239.500 ;
  LAYER VI3 ;
  RECT 4.740 239.220 4.940 239.420 ;
  LAYER VI3 ;
  RECT 4.340 239.220 4.540 239.420 ;
  LAYER VI2 ;
  RECT 4.280 239.220 5.140 239.500 ;
  LAYER VI2 ;
  RECT 4.740 239.220 4.940 239.420 ;
  LAYER VI2 ;
  RECT 4.340 239.220 4.540 239.420 ;
  LAYER VI3 ;
  RECT 4.280 242.900 5.140 243.180 ;
  LAYER VI3 ;
  RECT 4.740 242.900 4.940 243.100 ;
  LAYER VI3 ;
  RECT 4.340 242.900 4.540 243.100 ;
  LAYER VI2 ;
  RECT 4.280 242.900 5.140 243.180 ;
  LAYER VI2 ;
  RECT 4.740 242.900 4.940 243.100 ;
  LAYER VI2 ;
  RECT 4.340 242.900 4.540 243.100 ;
  LAYER VI3 ;
  RECT 4.280 246.580 5.140 246.860 ;
  LAYER VI3 ;
  RECT 4.740 246.580 4.940 246.780 ;
  LAYER VI3 ;
  RECT 4.340 246.580 4.540 246.780 ;
  LAYER VI2 ;
  RECT 4.280 246.580 5.140 246.860 ;
  LAYER VI2 ;
  RECT 4.740 246.580 4.940 246.780 ;
  LAYER VI2 ;
  RECT 4.340 246.580 4.540 246.780 ;
  LAYER VI3 ;
  RECT 4.280 250.260 5.140 250.540 ;
  LAYER VI3 ;
  RECT 4.740 250.260 4.940 250.460 ;
  LAYER VI3 ;
  RECT 4.340 250.260 4.540 250.460 ;
  LAYER VI2 ;
  RECT 4.280 250.260 5.140 250.540 ;
  LAYER VI2 ;
  RECT 4.740 250.260 4.940 250.460 ;
  LAYER VI2 ;
  RECT 4.340 250.260 4.540 250.460 ;
  LAYER VI3 ;
  RECT 4.280 253.940 5.140 254.220 ;
  LAYER VI3 ;
  RECT 4.740 253.940 4.940 254.140 ;
  LAYER VI3 ;
  RECT 4.340 253.940 4.540 254.140 ;
  LAYER VI2 ;
  RECT 4.280 253.940 5.140 254.220 ;
  LAYER VI2 ;
  RECT 4.740 253.940 4.940 254.140 ;
  LAYER VI2 ;
  RECT 4.340 253.940 4.540 254.140 ;
  LAYER VI3 ;
  RECT 4.280 257.620 5.140 257.900 ;
  LAYER VI3 ;
  RECT 4.740 257.620 4.940 257.820 ;
  LAYER VI3 ;
  RECT 4.340 257.620 4.540 257.820 ;
  LAYER VI2 ;
  RECT 4.280 257.620 5.140 257.900 ;
  LAYER VI2 ;
  RECT 4.740 257.620 4.940 257.820 ;
  LAYER VI2 ;
  RECT 4.340 257.620 4.540 257.820 ;
  LAYER VI3 ;
  RECT 4.280 261.300 5.140 261.580 ;
  LAYER VI3 ;
  RECT 4.740 261.300 4.940 261.500 ;
  LAYER VI3 ;
  RECT 4.340 261.300 4.540 261.500 ;
  LAYER VI2 ;
  RECT 4.280 261.300 5.140 261.580 ;
  LAYER VI2 ;
  RECT 4.740 261.300 4.940 261.500 ;
  LAYER VI2 ;
  RECT 4.340 261.300 4.540 261.500 ;
  LAYER VI3 ;
  RECT 4.280 264.980 5.140 265.260 ;
  LAYER VI3 ;
  RECT 4.740 264.980 4.940 265.180 ;
  LAYER VI3 ;
  RECT 4.340 264.980 4.540 265.180 ;
  LAYER VI2 ;
  RECT 4.280 264.980 5.140 265.260 ;
  LAYER VI2 ;
  RECT 4.740 264.980 4.940 265.180 ;
  LAYER VI2 ;
  RECT 4.340 264.980 4.540 265.180 ;
  LAYER VI3 ;
  RECT 4.280 268.660 5.140 268.940 ;
  LAYER VI3 ;
  RECT 4.740 268.660 4.940 268.860 ;
  LAYER VI3 ;
  RECT 4.340 268.660 4.540 268.860 ;
  LAYER VI2 ;
  RECT 4.280 268.660 5.140 268.940 ;
  LAYER VI2 ;
  RECT 4.740 268.660 4.940 268.860 ;
  LAYER VI2 ;
  RECT 4.340 268.660 4.540 268.860 ;
  LAYER VI3 ;
  RECT 4.280 272.340 5.140 272.620 ;
  LAYER VI3 ;
  RECT 4.740 272.340 4.940 272.540 ;
  LAYER VI3 ;
  RECT 4.340 272.340 4.540 272.540 ;
  LAYER VI2 ;
  RECT 4.280 272.340 5.140 272.620 ;
  LAYER VI2 ;
  RECT 4.740 272.340 4.940 272.540 ;
  LAYER VI2 ;
  RECT 4.340 272.340 4.540 272.540 ;
  LAYER VI3 ;
  RECT 4.280 276.020 5.140 276.300 ;
  LAYER VI3 ;
  RECT 4.740 276.020 4.940 276.220 ;
  LAYER VI3 ;
  RECT 4.340 276.020 4.540 276.220 ;
  LAYER VI2 ;
  RECT 4.280 276.020 5.140 276.300 ;
  LAYER VI2 ;
  RECT 4.740 276.020 4.940 276.220 ;
  LAYER VI2 ;
  RECT 4.340 276.020 4.540 276.220 ;
  LAYER VI3 ;
  RECT 4.280 279.700 5.140 279.980 ;
  LAYER VI3 ;
  RECT 4.740 279.700 4.940 279.900 ;
  LAYER VI3 ;
  RECT 4.340 279.700 4.540 279.900 ;
  LAYER VI2 ;
  RECT 4.280 279.700 5.140 279.980 ;
  LAYER VI2 ;
  RECT 4.740 279.700 4.940 279.900 ;
  LAYER VI2 ;
  RECT 4.340 279.700 4.540 279.900 ;
  LAYER VI3 ;
  RECT 4.280 283.380 5.140 283.660 ;
  LAYER VI3 ;
  RECT 4.740 283.380 4.940 283.580 ;
  LAYER VI3 ;
  RECT 4.340 283.380 4.540 283.580 ;
  LAYER VI2 ;
  RECT 4.280 283.380 5.140 283.660 ;
  LAYER VI2 ;
  RECT 4.740 283.380 4.940 283.580 ;
  LAYER VI2 ;
  RECT 4.340 283.380 4.540 283.580 ;
  LAYER VI3 ;
  RECT 4.280 287.060 5.140 287.340 ;
  LAYER VI3 ;
  RECT 4.740 287.060 4.940 287.260 ;
  LAYER VI3 ;
  RECT 4.340 287.060 4.540 287.260 ;
  LAYER VI2 ;
  RECT 4.280 287.060 5.140 287.340 ;
  LAYER VI2 ;
  RECT 4.740 287.060 4.940 287.260 ;
  LAYER VI2 ;
  RECT 4.340 287.060 4.540 287.260 ;
  LAYER VI3 ;
  RECT 4.280 290.740 5.140 291.020 ;
  LAYER VI3 ;
  RECT 4.740 290.740 4.940 290.940 ;
  LAYER VI3 ;
  RECT 4.340 290.740 4.540 290.940 ;
  LAYER VI2 ;
  RECT 4.280 290.740 5.140 291.020 ;
  LAYER VI2 ;
  RECT 4.740 290.740 4.940 290.940 ;
  LAYER VI2 ;
  RECT 4.340 290.740 4.540 290.940 ;
  LAYER VI3 ;
  RECT 4.280 294.420 5.140 294.700 ;
  LAYER VI3 ;
  RECT 4.740 294.420 4.940 294.620 ;
  LAYER VI3 ;
  RECT 4.340 294.420 4.540 294.620 ;
  LAYER VI2 ;
  RECT 4.280 294.420 5.140 294.700 ;
  LAYER VI2 ;
  RECT 4.740 294.420 4.940 294.620 ;
  LAYER VI2 ;
  RECT 4.340 294.420 4.540 294.620 ;
  LAYER VI3 ;
  RECT 4.280 298.100 5.140 298.380 ;
  LAYER VI3 ;
  RECT 4.740 298.100 4.940 298.300 ;
  LAYER VI3 ;
  RECT 4.340 298.100 4.540 298.300 ;
  LAYER VI2 ;
  RECT 4.280 298.100 5.140 298.380 ;
  LAYER VI2 ;
  RECT 4.740 298.100 4.940 298.300 ;
  LAYER VI2 ;
  RECT 4.340 298.100 4.540 298.300 ;
  LAYER VI3 ;
  RECT 4.280 301.780 5.140 302.060 ;
  LAYER VI3 ;
  RECT 4.740 301.780 4.940 301.980 ;
  LAYER VI3 ;
  RECT 4.340 301.780 4.540 301.980 ;
  LAYER VI2 ;
  RECT 4.280 301.780 5.140 302.060 ;
  LAYER VI2 ;
  RECT 4.740 301.780 4.940 301.980 ;
  LAYER VI2 ;
  RECT 4.340 301.780 4.540 301.980 ;
  LAYER VI3 ;
  RECT 4.280 305.460 5.140 305.740 ;
  LAYER VI3 ;
  RECT 4.740 305.460 4.940 305.660 ;
  LAYER VI3 ;
  RECT 4.340 305.460 4.540 305.660 ;
  LAYER VI2 ;
  RECT 4.280 305.460 5.140 305.740 ;
  LAYER VI2 ;
  RECT 4.740 305.460 4.940 305.660 ;
  LAYER VI2 ;
  RECT 4.340 305.460 4.540 305.660 ;
  LAYER VI3 ;
  RECT 4.280 309.140 5.140 309.420 ;
  LAYER VI3 ;
  RECT 4.740 309.140 4.940 309.340 ;
  LAYER VI3 ;
  RECT 4.340 309.140 4.540 309.340 ;
  LAYER VI2 ;
  RECT 4.280 309.140 5.140 309.420 ;
  LAYER VI2 ;
  RECT 4.740 309.140 4.940 309.340 ;
  LAYER VI2 ;
  RECT 4.340 309.140 4.540 309.340 ;
  LAYER VI3 ;
  RECT 4.280 312.820 5.140 313.100 ;
  LAYER VI3 ;
  RECT 4.740 312.820 4.940 313.020 ;
  LAYER VI3 ;
  RECT 4.340 312.820 4.540 313.020 ;
  LAYER VI2 ;
  RECT 4.280 312.820 5.140 313.100 ;
  LAYER VI2 ;
  RECT 4.740 312.820 4.940 313.020 ;
  LAYER VI2 ;
  RECT 4.340 312.820 4.540 313.020 ;
  LAYER VI3 ;
  RECT 4.280 316.500 5.140 316.780 ;
  LAYER VI3 ;
  RECT 4.740 316.500 4.940 316.700 ;
  LAYER VI3 ;
  RECT 4.340 316.500 4.540 316.700 ;
  LAYER VI2 ;
  RECT 4.280 316.500 5.140 316.780 ;
  LAYER VI2 ;
  RECT 4.740 316.500 4.940 316.700 ;
  LAYER VI2 ;
  RECT 4.340 316.500 4.540 316.700 ;
  LAYER VI3 ;
  RECT 4.280 320.180 5.140 320.460 ;
  LAYER VI3 ;
  RECT 4.740 320.180 4.940 320.380 ;
  LAYER VI3 ;
  RECT 4.340 320.180 4.540 320.380 ;
  LAYER VI2 ;
  RECT 4.280 320.180 5.140 320.460 ;
  LAYER VI2 ;
  RECT 4.740 320.180 4.940 320.380 ;
  LAYER VI2 ;
  RECT 4.340 320.180 4.540 320.380 ;
  LAYER VI3 ;
  RECT 4.280 323.860 5.140 324.140 ;
  LAYER VI3 ;
  RECT 4.740 323.860 4.940 324.060 ;
  LAYER VI3 ;
  RECT 4.340 323.860 4.540 324.060 ;
  LAYER VI2 ;
  RECT 4.280 323.860 5.140 324.140 ;
  LAYER VI2 ;
  RECT 4.740 323.860 4.940 324.060 ;
  LAYER VI2 ;
  RECT 4.340 323.860 4.540 324.060 ;
  LAYER VI3 ;
  RECT 4.280 327.540 5.140 327.820 ;
  LAYER VI3 ;
  RECT 4.740 327.540 4.940 327.740 ;
  LAYER VI3 ;
  RECT 4.340 327.540 4.540 327.740 ;
  LAYER VI2 ;
  RECT 4.280 327.540 5.140 327.820 ;
  LAYER VI2 ;
  RECT 4.740 327.540 4.940 327.740 ;
  LAYER VI2 ;
  RECT 4.340 327.540 4.540 327.740 ;
  LAYER VI3 ;
  RECT 4.280 331.220 5.140 331.500 ;
  LAYER VI3 ;
  RECT 4.740 331.220 4.940 331.420 ;
  LAYER VI3 ;
  RECT 4.340 331.220 4.540 331.420 ;
  LAYER VI2 ;
  RECT 4.280 331.220 5.140 331.500 ;
  LAYER VI2 ;
  RECT 4.740 331.220 4.940 331.420 ;
  LAYER VI2 ;
  RECT 4.340 331.220 4.540 331.420 ;
  LAYER VI3 ;
  RECT 4.280 334.900 5.140 335.180 ;
  LAYER VI3 ;
  RECT 4.740 334.900 4.940 335.100 ;
  LAYER VI3 ;
  RECT 4.340 334.900 4.540 335.100 ;
  LAYER VI2 ;
  RECT 4.280 334.900 5.140 335.180 ;
  LAYER VI2 ;
  RECT 4.740 334.900 4.940 335.100 ;
  LAYER VI2 ;
  RECT 4.340 334.900 4.540 335.100 ;
  LAYER VI3 ;
  RECT 4.280 338.580 5.140 338.860 ;
  LAYER VI3 ;
  RECT 4.740 338.580 4.940 338.780 ;
  LAYER VI3 ;
  RECT 4.340 338.580 4.540 338.780 ;
  LAYER VI2 ;
  RECT 4.280 338.580 5.140 338.860 ;
  LAYER VI2 ;
  RECT 4.740 338.580 4.940 338.780 ;
  LAYER VI2 ;
  RECT 4.340 338.580 4.540 338.780 ;
  LAYER VI3 ;
  RECT 4.280 342.260 5.140 342.540 ;
  LAYER VI3 ;
  RECT 4.740 342.260 4.940 342.460 ;
  LAYER VI3 ;
  RECT 4.340 342.260 4.540 342.460 ;
  LAYER VI2 ;
  RECT 4.280 342.260 5.140 342.540 ;
  LAYER VI2 ;
  RECT 4.740 342.260 4.940 342.460 ;
  LAYER VI2 ;
  RECT 4.340 342.260 4.540 342.460 ;
  LAYER VI3 ;
  RECT 4.280 345.940 5.140 346.220 ;
  LAYER VI3 ;
  RECT 4.740 345.940 4.940 346.140 ;
  LAYER VI3 ;
  RECT 4.340 345.940 4.540 346.140 ;
  LAYER VI2 ;
  RECT 4.280 345.940 5.140 346.220 ;
  LAYER VI2 ;
  RECT 4.740 345.940 4.940 346.140 ;
  LAYER VI2 ;
  RECT 4.340 345.940 4.540 346.140 ;
  LAYER VI3 ;
  RECT 4.280 349.620 5.140 349.900 ;
  LAYER VI3 ;
  RECT 4.740 349.620 4.940 349.820 ;
  LAYER VI3 ;
  RECT 4.340 349.620 4.540 349.820 ;
  LAYER VI2 ;
  RECT 4.280 349.620 5.140 349.900 ;
  LAYER VI2 ;
  RECT 4.740 349.620 4.940 349.820 ;
  LAYER VI2 ;
  RECT 4.340 349.620 4.540 349.820 ;
  LAYER VI3 ;
  RECT 4.280 353.300 5.140 353.580 ;
  LAYER VI3 ;
  RECT 4.740 353.300 4.940 353.500 ;
  LAYER VI3 ;
  RECT 4.340 353.300 4.540 353.500 ;
  LAYER VI2 ;
  RECT 4.280 353.300 5.140 353.580 ;
  LAYER VI2 ;
  RECT 4.740 353.300 4.940 353.500 ;
  LAYER VI2 ;
  RECT 4.340 353.300 4.540 353.500 ;
  LAYER VI3 ;
  RECT 4.280 356.980 5.140 357.260 ;
  LAYER VI3 ;
  RECT 4.740 356.980 4.940 357.180 ;
  LAYER VI3 ;
  RECT 4.340 356.980 4.540 357.180 ;
  LAYER VI2 ;
  RECT 4.280 356.980 5.140 357.260 ;
  LAYER VI2 ;
  RECT 4.740 356.980 4.940 357.180 ;
  LAYER VI2 ;
  RECT 4.340 356.980 4.540 357.180 ;
  LAYER VI3 ;
  RECT 4.280 360.660 5.140 360.940 ;
  LAYER VI3 ;
  RECT 4.740 360.660 4.940 360.860 ;
  LAYER VI3 ;
  RECT 4.340 360.660 4.540 360.860 ;
  LAYER VI2 ;
  RECT 4.280 360.660 5.140 360.940 ;
  LAYER VI2 ;
  RECT 4.740 360.660 4.940 360.860 ;
  LAYER VI2 ;
  RECT 4.340 360.660 4.540 360.860 ;
  LAYER VI3 ;
  RECT 4.280 364.340 5.140 364.620 ;
  LAYER VI3 ;
  RECT 4.740 364.340 4.940 364.540 ;
  LAYER VI3 ;
  RECT 4.340 364.340 4.540 364.540 ;
  LAYER VI2 ;
  RECT 4.280 364.340 5.140 364.620 ;
  LAYER VI2 ;
  RECT 4.740 364.340 4.940 364.540 ;
  LAYER VI2 ;
  RECT 4.340 364.340 4.540 364.540 ;
  LAYER VI3 ;
  RECT 4.280 368.020 5.140 368.300 ;
  LAYER VI3 ;
  RECT 4.740 368.020 4.940 368.220 ;
  LAYER VI3 ;
  RECT 4.340 368.020 4.540 368.220 ;
  LAYER VI2 ;
  RECT 4.280 368.020 5.140 368.300 ;
  LAYER VI2 ;
  RECT 4.740 368.020 4.940 368.220 ;
  LAYER VI2 ;
  RECT 4.340 368.020 4.540 368.220 ;
  LAYER VI3 ;
  RECT 4.280 371.700 5.140 371.980 ;
  LAYER VI3 ;
  RECT 4.740 371.700 4.940 371.900 ;
  LAYER VI3 ;
  RECT 4.340 371.700 4.540 371.900 ;
  LAYER VI2 ;
  RECT 4.280 371.700 5.140 371.980 ;
  LAYER VI2 ;
  RECT 4.740 371.700 4.940 371.900 ;
  LAYER VI2 ;
  RECT 4.340 371.700 4.540 371.900 ;
  LAYER VI3 ;
  RECT 4.280 375.380 5.140 375.660 ;
  LAYER VI3 ;
  RECT 4.740 375.380 4.940 375.580 ;
  LAYER VI3 ;
  RECT 4.340 375.380 4.540 375.580 ;
  LAYER VI2 ;
  RECT 4.280 375.380 5.140 375.660 ;
  LAYER VI2 ;
  RECT 4.740 375.380 4.940 375.580 ;
  LAYER VI2 ;
  RECT 4.340 375.380 4.540 375.580 ;
  LAYER VI3 ;
  RECT 4.280 379.060 5.140 379.340 ;
  LAYER VI3 ;
  RECT 4.740 379.060 4.940 379.260 ;
  LAYER VI3 ;
  RECT 4.340 379.060 4.540 379.260 ;
  LAYER VI2 ;
  RECT 4.280 379.060 5.140 379.340 ;
  LAYER VI2 ;
  RECT 4.740 379.060 4.940 379.260 ;
  LAYER VI2 ;
  RECT 4.340 379.060 4.540 379.260 ;
  LAYER VI3 ;
  RECT 4.280 382.740 5.140 383.020 ;
  LAYER VI3 ;
  RECT 4.740 382.740 4.940 382.940 ;
  LAYER VI3 ;
  RECT 4.340 382.740 4.540 382.940 ;
  LAYER VI2 ;
  RECT 4.280 382.740 5.140 383.020 ;
  LAYER VI2 ;
  RECT 4.740 382.740 4.940 382.940 ;
  LAYER VI2 ;
  RECT 4.340 382.740 4.540 382.940 ;
  LAYER VI3 ;
  RECT 4.280 386.420 5.140 386.700 ;
  LAYER VI3 ;
  RECT 4.740 386.420 4.940 386.620 ;
  LAYER VI3 ;
  RECT 4.340 386.420 4.540 386.620 ;
  LAYER VI2 ;
  RECT 4.280 386.420 5.140 386.700 ;
  LAYER VI2 ;
  RECT 4.740 386.420 4.940 386.620 ;
  LAYER VI2 ;
  RECT 4.340 386.420 4.540 386.620 ;
  LAYER VI3 ;
  RECT 4.280 390.100 5.140 390.380 ;
  LAYER VI3 ;
  RECT 4.740 390.100 4.940 390.300 ;
  LAYER VI3 ;
  RECT 4.340 390.100 4.540 390.300 ;
  LAYER VI2 ;
  RECT 4.280 390.100 5.140 390.380 ;
  LAYER VI2 ;
  RECT 4.740 390.100 4.940 390.300 ;
  LAYER VI2 ;
  RECT 4.340 390.100 4.540 390.300 ;
  LAYER VI3 ;
  RECT 4.280 393.780 5.140 394.060 ;
  LAYER VI3 ;
  RECT 4.740 393.780 4.940 393.980 ;
  LAYER VI3 ;
  RECT 4.340 393.780 4.540 393.980 ;
  LAYER VI2 ;
  RECT 4.280 393.780 5.140 394.060 ;
  LAYER VI2 ;
  RECT 4.740 393.780 4.940 393.980 ;
  LAYER VI2 ;
  RECT 4.340 393.780 4.540 393.980 ;
  LAYER VI3 ;
  RECT 4.280 397.460 5.140 397.740 ;
  LAYER VI3 ;
  RECT 4.740 397.460 4.940 397.660 ;
  LAYER VI3 ;
  RECT 4.340 397.460 4.540 397.660 ;
  LAYER VI2 ;
  RECT 4.280 397.460 5.140 397.740 ;
  LAYER VI2 ;
  RECT 4.740 397.460 4.940 397.660 ;
  LAYER VI2 ;
  RECT 4.340 397.460 4.540 397.660 ;
  LAYER VI3 ;
  RECT 4.280 401.140 5.140 401.420 ;
  LAYER VI3 ;
  RECT 4.740 401.140 4.940 401.340 ;
  LAYER VI3 ;
  RECT 4.340 401.140 4.540 401.340 ;
  LAYER VI2 ;
  RECT 4.280 401.140 5.140 401.420 ;
  LAYER VI2 ;
  RECT 4.740 401.140 4.940 401.340 ;
  LAYER VI2 ;
  RECT 4.340 401.140 4.540 401.340 ;
  LAYER VI3 ;
  RECT 4.280 404.820 5.140 405.100 ;
  LAYER VI3 ;
  RECT 4.740 404.820 4.940 405.020 ;
  LAYER VI3 ;
  RECT 4.340 404.820 4.540 405.020 ;
  LAYER VI2 ;
  RECT 4.280 404.820 5.140 405.100 ;
  LAYER VI2 ;
  RECT 4.740 404.820 4.940 405.020 ;
  LAYER VI2 ;
  RECT 4.340 404.820 4.540 405.020 ;
  LAYER VI3 ;
  RECT 4.280 408.500 5.140 408.780 ;
  LAYER VI3 ;
  RECT 4.740 408.500 4.940 408.700 ;
  LAYER VI3 ;
  RECT 4.340 408.500 4.540 408.700 ;
  LAYER VI2 ;
  RECT 4.280 408.500 5.140 408.780 ;
  LAYER VI2 ;
  RECT 4.740 408.500 4.940 408.700 ;
  LAYER VI2 ;
  RECT 4.340 408.500 4.540 408.700 ;
  LAYER VI3 ;
  RECT 4.280 412.180 5.140 412.460 ;
  LAYER VI3 ;
  RECT 4.740 412.180 4.940 412.380 ;
  LAYER VI3 ;
  RECT 4.340 412.180 4.540 412.380 ;
  LAYER VI2 ;
  RECT 4.280 412.180 5.140 412.460 ;
  LAYER VI2 ;
  RECT 4.740 412.180 4.940 412.380 ;
  LAYER VI2 ;
  RECT 4.340 412.180 4.540 412.380 ;
  LAYER VI3 ;
  RECT 4.280 415.860 5.140 416.140 ;
  LAYER VI3 ;
  RECT 4.740 415.860 4.940 416.060 ;
  LAYER VI3 ;
  RECT 4.340 415.860 4.540 416.060 ;
  LAYER VI2 ;
  RECT 4.280 415.860 5.140 416.140 ;
  LAYER VI2 ;
  RECT 4.740 415.860 4.940 416.060 ;
  LAYER VI2 ;
  RECT 4.340 415.860 4.540 416.060 ;
  LAYER VI3 ;
  RECT 4.280 419.540 5.140 419.820 ;
  LAYER VI3 ;
  RECT 4.740 419.540 4.940 419.740 ;
  LAYER VI3 ;
  RECT 4.340 419.540 4.540 419.740 ;
  LAYER VI2 ;
  RECT 4.280 419.540 5.140 419.820 ;
  LAYER VI2 ;
  RECT 4.740 419.540 4.940 419.740 ;
  LAYER VI2 ;
  RECT 4.340 419.540 4.540 419.740 ;
  LAYER VI3 ;
  RECT 4.280 423.220 5.140 423.500 ;
  LAYER VI3 ;
  RECT 4.740 423.220 4.940 423.420 ;
  LAYER VI3 ;
  RECT 4.340 423.220 4.540 423.420 ;
  LAYER VI2 ;
  RECT 4.280 423.220 5.140 423.500 ;
  LAYER VI2 ;
  RECT 4.740 423.220 4.940 423.420 ;
  LAYER VI2 ;
  RECT 4.340 423.220 4.540 423.420 ;
  LAYER VI3 ;
  RECT 4.280 426.900 5.140 427.180 ;
  LAYER VI3 ;
  RECT 4.740 426.900 4.940 427.100 ;
  LAYER VI3 ;
  RECT 4.340 426.900 4.540 427.100 ;
  LAYER VI2 ;
  RECT 4.280 426.900 5.140 427.180 ;
  LAYER VI2 ;
  RECT 4.740 426.900 4.940 427.100 ;
  LAYER VI2 ;
  RECT 4.340 426.900 4.540 427.100 ;
  LAYER VI3 ;
  RECT 4.280 430.580 5.140 430.860 ;
  LAYER VI3 ;
  RECT 4.740 430.580 4.940 430.780 ;
  LAYER VI3 ;
  RECT 4.340 430.580 4.540 430.780 ;
  LAYER VI2 ;
  RECT 4.280 430.580 5.140 430.860 ;
  LAYER VI2 ;
  RECT 4.740 430.580 4.940 430.780 ;
  LAYER VI2 ;
  RECT 4.340 430.580 4.540 430.780 ;
  LAYER VI3 ;
  RECT 4.280 434.260 5.140 434.540 ;
  LAYER VI3 ;
  RECT 4.740 434.260 4.940 434.460 ;
  LAYER VI3 ;
  RECT 4.340 434.260 4.540 434.460 ;
  LAYER VI2 ;
  RECT 4.280 434.260 5.140 434.540 ;
  LAYER VI2 ;
  RECT 4.740 434.260 4.940 434.460 ;
  LAYER VI2 ;
  RECT 4.340 434.260 4.540 434.460 ;
  LAYER VI3 ;
  RECT 4.280 437.940 5.140 438.220 ;
  LAYER VI3 ;
  RECT 4.740 437.940 4.940 438.140 ;
  LAYER VI3 ;
  RECT 4.340 437.940 4.540 438.140 ;
  LAYER VI2 ;
  RECT 4.280 437.940 5.140 438.220 ;
  LAYER VI2 ;
  RECT 4.740 437.940 4.940 438.140 ;
  LAYER VI2 ;
  RECT 4.340 437.940 4.540 438.140 ;
  LAYER VI3 ;
  RECT 4.280 441.620 5.140 441.900 ;
  LAYER VI3 ;
  RECT 4.740 441.620 4.940 441.820 ;
  LAYER VI3 ;
  RECT 4.340 441.620 4.540 441.820 ;
  LAYER VI2 ;
  RECT 4.280 441.620 5.140 441.900 ;
  LAYER VI2 ;
  RECT 4.740 441.620 4.940 441.820 ;
  LAYER VI2 ;
  RECT 4.340 441.620 4.540 441.820 ;
  LAYER VI3 ;
  RECT 4.280 445.300 5.140 445.580 ;
  LAYER VI3 ;
  RECT 4.740 445.300 4.940 445.500 ;
  LAYER VI3 ;
  RECT 4.340 445.300 4.540 445.500 ;
  LAYER VI2 ;
  RECT 4.280 445.300 5.140 445.580 ;
  LAYER VI2 ;
  RECT 4.740 445.300 4.940 445.500 ;
  LAYER VI2 ;
  RECT 4.340 445.300 4.540 445.500 ;
  LAYER VI3 ;
  RECT 4.280 448.980 5.140 449.260 ;
  LAYER VI3 ;
  RECT 4.740 448.980 4.940 449.180 ;
  LAYER VI3 ;
  RECT 4.340 448.980 4.540 449.180 ;
  LAYER VI2 ;
  RECT 4.280 448.980 5.140 449.260 ;
  LAYER VI2 ;
  RECT 4.740 448.980 4.940 449.180 ;
  LAYER VI2 ;
  RECT 4.340 448.980 4.540 449.180 ;
  LAYER VI3 ;
  RECT 4.280 452.660 5.140 452.940 ;
  LAYER VI3 ;
  RECT 4.740 452.660 4.940 452.860 ;
  LAYER VI3 ;
  RECT 4.340 452.660 4.540 452.860 ;
  LAYER VI2 ;
  RECT 4.280 452.660 5.140 452.940 ;
  LAYER VI2 ;
  RECT 4.740 452.660 4.940 452.860 ;
  LAYER VI2 ;
  RECT 4.340 452.660 4.540 452.860 ;
  LAYER VI3 ;
  RECT 4.280 456.340 5.140 456.620 ;
  LAYER VI3 ;
  RECT 4.740 456.340 4.940 456.540 ;
  LAYER VI3 ;
  RECT 4.340 456.340 4.540 456.540 ;
  LAYER VI2 ;
  RECT 4.280 456.340 5.140 456.620 ;
  LAYER VI2 ;
  RECT 4.740 456.340 4.940 456.540 ;
  LAYER VI2 ;
  RECT 4.340 456.340 4.540 456.540 ;
  LAYER VI3 ;
  RECT 4.280 460.020 5.140 460.300 ;
  LAYER VI3 ;
  RECT 4.740 460.020 4.940 460.220 ;
  LAYER VI3 ;
  RECT 4.340 460.020 4.540 460.220 ;
  LAYER VI2 ;
  RECT 4.280 460.020 5.140 460.300 ;
  LAYER VI2 ;
  RECT 4.740 460.020 4.940 460.220 ;
  LAYER VI2 ;
  RECT 4.340 460.020 4.540 460.220 ;
  LAYER VI3 ;
  RECT 4.280 463.700 5.140 463.980 ;
  LAYER VI3 ;
  RECT 4.740 463.700 4.940 463.900 ;
  LAYER VI3 ;
  RECT 4.340 463.700 4.540 463.900 ;
  LAYER VI2 ;
  RECT 4.280 463.700 5.140 463.980 ;
  LAYER VI2 ;
  RECT 4.740 463.700 4.940 463.900 ;
  LAYER VI2 ;
  RECT 4.340 463.700 4.540 463.900 ;
  LAYER VI3 ;
  RECT 4.280 467.380 5.140 467.660 ;
  LAYER VI3 ;
  RECT 4.740 467.380 4.940 467.580 ;
  LAYER VI3 ;
  RECT 4.340 467.380 4.540 467.580 ;
  LAYER VI2 ;
  RECT 4.280 467.380 5.140 467.660 ;
  LAYER VI2 ;
  RECT 4.740 467.380 4.940 467.580 ;
  LAYER VI2 ;
  RECT 4.340 467.380 4.540 467.580 ;
  LAYER VI3 ;
  RECT 4.280 471.060 5.140 471.340 ;
  LAYER VI3 ;
  RECT 4.740 471.060 4.940 471.260 ;
  LAYER VI3 ;
  RECT 4.340 471.060 4.540 471.260 ;
  LAYER VI2 ;
  RECT 4.280 471.060 5.140 471.340 ;
  LAYER VI2 ;
  RECT 4.740 471.060 4.940 471.260 ;
  LAYER VI2 ;
  RECT 4.340 471.060 4.540 471.260 ;
  LAYER VI3 ;
  RECT 4.280 474.740 5.140 475.020 ;
  LAYER VI3 ;
  RECT 4.740 474.740 4.940 474.940 ;
  LAYER VI3 ;
  RECT 4.340 474.740 4.540 474.940 ;
  LAYER VI2 ;
  RECT 4.280 474.740 5.140 475.020 ;
  LAYER VI2 ;
  RECT 4.740 474.740 4.940 474.940 ;
  LAYER VI2 ;
  RECT 4.340 474.740 4.540 474.940 ;
  LAYER VI3 ;
  RECT 4.280 478.420 5.140 478.700 ;
  LAYER VI3 ;
  RECT 4.740 478.420 4.940 478.620 ;
  LAYER VI3 ;
  RECT 4.340 478.420 4.540 478.620 ;
  LAYER VI2 ;
  RECT 4.280 478.420 5.140 478.700 ;
  LAYER VI2 ;
  RECT 4.740 478.420 4.940 478.620 ;
  LAYER VI2 ;
  RECT 4.340 478.420 4.540 478.620 ;
  LAYER VI3 ;
  RECT 4.280 482.100 5.140 482.380 ;
  LAYER VI3 ;
  RECT 4.740 482.100 4.940 482.300 ;
  LAYER VI3 ;
  RECT 4.340 482.100 4.540 482.300 ;
  LAYER VI2 ;
  RECT 4.280 482.100 5.140 482.380 ;
  LAYER VI2 ;
  RECT 4.740 482.100 4.940 482.300 ;
  LAYER VI2 ;
  RECT 4.340 482.100 4.540 482.300 ;
  LAYER VI3 ;
  RECT 4.280 485.780 5.140 486.060 ;
  LAYER VI3 ;
  RECT 4.740 485.780 4.940 485.980 ;
  LAYER VI3 ;
  RECT 4.340 485.780 4.540 485.980 ;
  LAYER VI2 ;
  RECT 4.280 485.780 5.140 486.060 ;
  LAYER VI2 ;
  RECT 4.740 485.780 4.940 485.980 ;
  LAYER VI2 ;
  RECT 4.340 485.780 4.540 485.980 ;
  LAYER VI3 ;
  RECT 4.280 489.460 5.140 489.740 ;
  LAYER VI3 ;
  RECT 4.740 489.460 4.940 489.660 ;
  LAYER VI3 ;
  RECT 4.340 489.460 4.540 489.660 ;
  LAYER VI2 ;
  RECT 4.280 489.460 5.140 489.740 ;
  LAYER VI2 ;
  RECT 4.740 489.460 4.940 489.660 ;
  LAYER VI2 ;
  RECT 4.340 489.460 4.540 489.660 ;
  LAYER VI3 ;
  RECT 4.280 493.140 5.140 493.420 ;
  LAYER VI3 ;
  RECT 4.740 493.140 4.940 493.340 ;
  LAYER VI3 ;
  RECT 4.340 493.140 4.540 493.340 ;
  LAYER VI2 ;
  RECT 4.280 493.140 5.140 493.420 ;
  LAYER VI2 ;
  RECT 4.740 493.140 4.940 493.340 ;
  LAYER VI2 ;
  RECT 4.340 493.140 4.540 493.340 ;
  LAYER VI3 ;
  RECT 4.280 496.820 5.140 497.100 ;
  LAYER VI3 ;
  RECT 4.740 496.820 4.940 497.020 ;
  LAYER VI3 ;
  RECT 4.340 496.820 4.540 497.020 ;
  LAYER VI2 ;
  RECT 4.280 496.820 5.140 497.100 ;
  LAYER VI2 ;
  RECT 4.740 496.820 4.940 497.020 ;
  LAYER VI2 ;
  RECT 4.340 496.820 4.540 497.020 ;
  LAYER VI3 ;
  RECT 4.280 500.500 5.140 500.780 ;
  LAYER VI3 ;
  RECT 4.740 500.500 4.940 500.700 ;
  LAYER VI3 ;
  RECT 4.340 500.500 4.540 500.700 ;
  LAYER VI2 ;
  RECT 4.280 500.500 5.140 500.780 ;
  LAYER VI2 ;
  RECT 4.740 500.500 4.940 500.700 ;
  LAYER VI2 ;
  RECT 4.340 500.500 4.540 500.700 ;
  LAYER VI3 ;
  RECT 4.280 504.180 5.140 504.460 ;
  LAYER VI3 ;
  RECT 4.740 504.180 4.940 504.380 ;
  LAYER VI3 ;
  RECT 4.340 504.180 4.540 504.380 ;
  LAYER VI2 ;
  RECT 4.280 504.180 5.140 504.460 ;
  LAYER VI2 ;
  RECT 4.740 504.180 4.940 504.380 ;
  LAYER VI2 ;
  RECT 4.340 504.180 4.540 504.380 ;
  LAYER VI3 ;
  RECT 4.280 507.860 5.140 508.140 ;
  LAYER VI3 ;
  RECT 4.740 507.860 4.940 508.060 ;
  LAYER VI3 ;
  RECT 4.340 507.860 4.540 508.060 ;
  LAYER VI2 ;
  RECT 4.280 507.860 5.140 508.140 ;
  LAYER VI2 ;
  RECT 4.740 507.860 4.940 508.060 ;
  LAYER VI2 ;
  RECT 4.340 507.860 4.540 508.060 ;
  LAYER VI3 ;
  RECT 4.280 511.540 5.140 511.820 ;
  LAYER VI3 ;
  RECT 4.740 511.540 4.940 511.740 ;
  LAYER VI3 ;
  RECT 4.340 511.540 4.540 511.740 ;
  LAYER VI2 ;
  RECT 4.280 511.540 5.140 511.820 ;
  LAYER VI2 ;
  RECT 4.740 511.540 4.940 511.740 ;
  LAYER VI2 ;
  RECT 4.340 511.540 4.540 511.740 ;
  LAYER VI3 ;
  RECT 4.280 515.220 5.140 515.500 ;
  LAYER VI3 ;
  RECT 4.740 515.220 4.940 515.420 ;
  LAYER VI3 ;
  RECT 4.340 515.220 4.540 515.420 ;
  LAYER VI2 ;
  RECT 4.280 515.220 5.140 515.500 ;
  LAYER VI2 ;
  RECT 4.740 515.220 4.940 515.420 ;
  LAYER VI2 ;
  RECT 4.340 515.220 4.540 515.420 ;
  LAYER VI3 ;
  RECT 4.280 518.900 5.140 519.180 ;
  LAYER VI3 ;
  RECT 4.740 518.900 4.940 519.100 ;
  LAYER VI3 ;
  RECT 4.340 518.900 4.540 519.100 ;
  LAYER VI2 ;
  RECT 4.280 518.900 5.140 519.180 ;
  LAYER VI2 ;
  RECT 4.740 518.900 4.940 519.100 ;
  LAYER VI2 ;
  RECT 4.340 518.900 4.540 519.100 ;
  LAYER VI3 ;
  RECT 4.280 522.580 5.140 522.860 ;
  LAYER VI3 ;
  RECT 4.740 522.580 4.940 522.780 ;
  LAYER VI3 ;
  RECT 4.340 522.580 4.540 522.780 ;
  LAYER VI2 ;
  RECT 4.280 522.580 5.140 522.860 ;
  LAYER VI2 ;
  RECT 4.740 522.580 4.940 522.780 ;
  LAYER VI2 ;
  RECT 4.340 522.580 4.540 522.780 ;
  LAYER VI3 ;
  RECT 4.280 526.260 5.140 526.540 ;
  LAYER VI3 ;
  RECT 4.740 526.260 4.940 526.460 ;
  LAYER VI3 ;
  RECT 4.340 526.260 4.540 526.460 ;
  LAYER VI2 ;
  RECT 4.280 526.260 5.140 526.540 ;
  LAYER VI2 ;
  RECT 4.740 526.260 4.940 526.460 ;
  LAYER VI2 ;
  RECT 4.340 526.260 4.540 526.460 ;
  LAYER VI3 ;
  RECT 4.280 529.940 5.140 530.220 ;
  LAYER VI3 ;
  RECT 4.740 529.940 4.940 530.140 ;
  LAYER VI3 ;
  RECT 4.340 529.940 4.540 530.140 ;
  LAYER VI2 ;
  RECT 4.280 529.940 5.140 530.220 ;
  LAYER VI2 ;
  RECT 4.740 529.940 4.940 530.140 ;
  LAYER VI2 ;
  RECT 4.340 529.940 4.540 530.140 ;
  LAYER VI3 ;
  RECT 4.280 533.620 5.140 533.900 ;
  LAYER VI3 ;
  RECT 4.740 533.620 4.940 533.820 ;
  LAYER VI3 ;
  RECT 4.340 533.620 4.540 533.820 ;
  LAYER VI2 ;
  RECT 4.280 533.620 5.140 533.900 ;
  LAYER VI2 ;
  RECT 4.740 533.620 4.940 533.820 ;
  LAYER VI2 ;
  RECT 4.340 533.620 4.540 533.820 ;
  LAYER VI3 ;
  RECT 4.280 537.300 5.140 537.580 ;
  LAYER VI3 ;
  RECT 4.740 537.300 4.940 537.500 ;
  LAYER VI3 ;
  RECT 4.340 537.300 4.540 537.500 ;
  LAYER VI2 ;
  RECT 4.280 537.300 5.140 537.580 ;
  LAYER VI2 ;
  RECT 4.740 537.300 4.940 537.500 ;
  LAYER VI2 ;
  RECT 4.340 537.300 4.540 537.500 ;
  LAYER VI3 ;
  RECT 4.280 545.220 5.140 545.600 ;
  LAYER VI3 ;
  RECT 4.680 545.280 4.880 545.480 ;
  LAYER VI3 ;
  RECT 4.280 545.280 4.480 545.480 ;
  LAYER VI2 ;
  RECT 4.280 545.220 5.140 545.600 ;
  LAYER VI2 ;
  RECT 4.680 545.280 4.880 545.480 ;
  LAYER VI2 ;
  RECT 4.280 545.280 4.480 545.480 ;
  LAYER VI3 ;
  RECT 47.350 546.070 47.600 546.930 ;
  LAYER VI3 ;
  RECT 47.350 546.530 47.550 546.730 ;
  LAYER VI3 ;
  RECT 47.350 546.130 47.550 546.330 ;
  LAYER VI2 ;
  RECT 47.350 546.070 47.600 546.930 ;
  LAYER VI2 ;
  RECT 47.350 546.530 47.550 546.730 ;
  LAYER VI2 ;
  RECT 47.350 546.130 47.550 546.330 ;
  LAYER VI3 ;
  RECT 88.270 546.070 88.520 546.930 ;
  LAYER VI3 ;
  RECT 88.270 546.530 88.470 546.730 ;
  LAYER VI3 ;
  RECT 88.270 546.130 88.470 546.330 ;
  LAYER VI2 ;
  RECT 88.270 546.070 88.520 546.930 ;
  LAYER VI2 ;
  RECT 88.270 546.530 88.470 546.730 ;
  LAYER VI2 ;
  RECT 88.270 546.130 88.470 546.330 ;
  LAYER VI3 ;
  RECT 129.190 546.070 129.440 546.930 ;
  LAYER VI3 ;
  RECT 129.190 546.530 129.390 546.730 ;
  LAYER VI3 ;
  RECT 129.190 546.130 129.390 546.330 ;
  LAYER VI2 ;
  RECT 129.190 546.070 129.440 546.930 ;
  LAYER VI2 ;
  RECT 129.190 546.530 129.390 546.730 ;
  LAYER VI2 ;
  RECT 129.190 546.130 129.390 546.330 ;
  LAYER VI3 ;
  RECT 170.110 546.070 170.360 546.930 ;
  LAYER VI3 ;
  RECT 170.110 546.530 170.310 546.730 ;
  LAYER VI3 ;
  RECT 170.110 546.130 170.310 546.330 ;
  LAYER VI2 ;
  RECT 170.110 546.070 170.360 546.930 ;
  LAYER VI2 ;
  RECT 170.110 546.530 170.310 546.730 ;
  LAYER VI2 ;
  RECT 170.110 546.130 170.310 546.330 ;
  LAYER VI3 ;
  RECT 211.030 546.070 211.280 546.930 ;
  LAYER VI3 ;
  RECT 211.030 546.530 211.230 546.730 ;
  LAYER VI3 ;
  RECT 211.030 546.130 211.230 546.330 ;
  LAYER VI2 ;
  RECT 211.030 546.070 211.280 546.930 ;
  LAYER VI2 ;
  RECT 211.030 546.530 211.230 546.730 ;
  LAYER VI2 ;
  RECT 211.030 546.130 211.230 546.330 ;
  LAYER VI3 ;
  RECT 251.950 546.070 252.200 546.930 ;
  LAYER VI3 ;
  RECT 251.950 546.530 252.150 546.730 ;
  LAYER VI3 ;
  RECT 251.950 546.130 252.150 546.330 ;
  LAYER VI2 ;
  RECT 251.950 546.070 252.200 546.930 ;
  LAYER VI2 ;
  RECT 251.950 546.530 252.150 546.730 ;
  LAYER VI2 ;
  RECT 251.950 546.130 252.150 546.330 ;
  LAYER VI3 ;
  RECT 292.870 546.070 293.120 546.930 ;
  LAYER VI3 ;
  RECT 292.870 546.530 293.070 546.730 ;
  LAYER VI3 ;
  RECT 292.870 546.130 293.070 546.330 ;
  LAYER VI2 ;
  RECT 292.870 546.070 293.120 546.930 ;
  LAYER VI2 ;
  RECT 292.870 546.530 293.070 546.730 ;
  LAYER VI2 ;
  RECT 292.870 546.130 293.070 546.330 ;
  LAYER VI3 ;
  RECT 333.790 546.070 334.040 546.930 ;
  LAYER VI3 ;
  RECT 333.790 546.530 333.990 546.730 ;
  LAYER VI3 ;
  RECT 333.790 546.130 333.990 546.330 ;
  LAYER VI2 ;
  RECT 333.790 546.070 334.040 546.930 ;
  LAYER VI2 ;
  RECT 333.790 546.530 333.990 546.730 ;
  LAYER VI2 ;
  RECT 333.790 546.130 333.990 546.330 ;
  LAYER VI3 ;
  RECT 374.710 546.070 374.960 546.930 ;
  LAYER VI3 ;
  RECT 374.710 546.530 374.910 546.730 ;
  LAYER VI3 ;
  RECT 374.710 546.130 374.910 546.330 ;
  LAYER VI2 ;
  RECT 374.710 546.070 374.960 546.930 ;
  LAYER VI2 ;
  RECT 374.710 546.530 374.910 546.730 ;
  LAYER VI2 ;
  RECT 374.710 546.130 374.910 546.330 ;
  LAYER VI3 ;
  RECT 415.630 546.070 415.880 546.930 ;
  LAYER VI3 ;
  RECT 415.630 546.530 415.830 546.730 ;
  LAYER VI3 ;
  RECT 415.630 546.130 415.830 546.330 ;
  LAYER VI2 ;
  RECT 415.630 546.070 415.880 546.930 ;
  LAYER VI2 ;
  RECT 415.630 546.530 415.830 546.730 ;
  LAYER VI2 ;
  RECT 415.630 546.130 415.830 546.330 ;
  LAYER VI3 ;
  RECT 456.550 546.070 456.800 546.930 ;
  LAYER VI3 ;
  RECT 456.550 546.530 456.750 546.730 ;
  LAYER VI3 ;
  RECT 456.550 546.130 456.750 546.330 ;
  LAYER VI2 ;
  RECT 456.550 546.070 456.800 546.930 ;
  LAYER VI2 ;
  RECT 456.550 546.530 456.750 546.730 ;
  LAYER VI2 ;
  RECT 456.550 546.130 456.750 546.330 ;
  LAYER VI3 ;
  RECT 497.470 546.070 497.720 546.930 ;
  LAYER VI3 ;
  RECT 497.470 546.530 497.670 546.730 ;
  LAYER VI3 ;
  RECT 497.470 546.130 497.670 546.330 ;
  LAYER VI2 ;
  RECT 497.470 546.070 497.720 546.930 ;
  LAYER VI2 ;
  RECT 497.470 546.530 497.670 546.730 ;
  LAYER VI2 ;
  RECT 497.470 546.130 497.670 546.330 ;
  LAYER VI3 ;
  RECT 538.390 546.070 538.640 546.930 ;
  LAYER VI3 ;
  RECT 538.390 546.530 538.590 546.730 ;
  LAYER VI3 ;
  RECT 538.390 546.130 538.590 546.330 ;
  LAYER VI2 ;
  RECT 538.390 546.070 538.640 546.930 ;
  LAYER VI2 ;
  RECT 538.390 546.530 538.590 546.730 ;
  LAYER VI2 ;
  RECT 538.390 546.130 538.590 546.330 ;
  LAYER VI3 ;
  RECT 579.310 546.070 579.560 546.930 ;
  LAYER VI3 ;
  RECT 579.310 546.530 579.510 546.730 ;
  LAYER VI3 ;
  RECT 579.310 546.130 579.510 546.330 ;
  LAYER VI2 ;
  RECT 579.310 546.070 579.560 546.930 ;
  LAYER VI2 ;
  RECT 579.310 546.530 579.510 546.730 ;
  LAYER VI2 ;
  RECT 579.310 546.130 579.510 546.330 ;
  LAYER VI3 ;
  RECT 620.230 546.070 620.480 546.930 ;
  LAYER VI3 ;
  RECT 620.230 546.530 620.430 546.730 ;
  LAYER VI3 ;
  RECT 620.230 546.130 620.430 546.330 ;
  LAYER VI2 ;
  RECT 620.230 546.070 620.480 546.930 ;
  LAYER VI2 ;
  RECT 620.230 546.530 620.430 546.730 ;
  LAYER VI2 ;
  RECT 620.230 546.130 620.430 546.330 ;
END
END SHKD110_4096X8X8BM1
END LIBRARY





