`timescale 1ns / 1ps

    // L2Cache_dataSRAM u_L2Cache_dataSRAM (
    //     .clka   (w_cfifo2_fire), 
    //     .ena    (1'b1),      
    //     .wea    (r_read_or_write_dataSRAM),     
    //     .addra  (r_dataSRAM_addr_10),  
    //     .dina   (r_dataSRAM_in_32B),   
    //     .douta  ({w_dataSRAM_out_way7_32B, w_dataSRAM_out_way6_32B, w_dataSRAM_out_way5_32B, w_dataSRAM_out_way4_32B, w_dataSRAM_out_way3_32B, w_dataSRAM_out_way2_32B, w_dataSRAM_out_way1_32B, w_dataSRAM_out_way0_32B})
    // );

module L2Cache_dataSRAM(
    input wire clka,ena,wea,  // fire ʹ��1 ��д01  // ena û����
    input wire [9:0] addra,   // ��ַ [9:3]:Ƭ��    [2:0]:Ƭѡ
    input wire [255:0] dina,
    output wire [2047:0] douta
);

    wire [6:0] RAM_addr;    // Ƭ��
    reg  [15:0] w_sel_SRAM_16;   // Ƭѡ
    wire [255:0] w_datain_256;

    wire [255:0] RAM7_data_in,  RAM6_data_in,  RAM5_data_in,  RAM4_data_in,  RAM3_data_in,  RAM2_data_in,  RAM1_data_in, RAM0_data_in;
    wire [255:0] RAM15_data_in, RAM14_data_in, RAM13_data_in, RAM12_data_in, RAM11_data_in, RAM10_data_in, RAM9_data_in, RAM8_data_in;
    
    wire [255:0] RAM7_data_out,  RAM6_data_out,  RAM5_data_out,  RAM4_data_out,  RAM3_data_out,  RAM2_data_out,  RAM1_data_out, RAM0_data_out;
    wire [255:0] RAM15_data_out, RAM14_data_out, RAM13_data_out, RAM12_data_out, RAM11_data_out, RAM10_data_out, RAM9_data_out, RAM8_data_out;

    assign RAM_addr = addra[9:3];   // Ƭ�ڵ�ַ

    assign w_datain_256 = dina;

    assign RAM15_data_in = {w_datain_256[255:128], 128'b0 };
    assign RAM14_data_in = { 128'b0, w_datain_256[127:0]};
    assign RAM13_data_in = {w_datain_256[255:128], 128'b0 };
    assign RAM12_data_in = { 128'b0, w_datain_256[127:0]};
    assign RAM11_data_in = {w_datain_256[255:128], 128'b0 };
    assign RAM10_data_in = { 128'b0, w_datain_256[127:0]};
    assign  RAM9_data_in = {w_datain_256[255:128], 128'b0 };
    assign  RAM8_data_in = { 128'b0, w_datain_256[127:0]};
    assign  RAM7_data_in = {w_datain_256[255:128], 128'b0 };
    assign  RAM6_data_in = { 128'b0, w_datain_256[127:0]};
    assign  RAM5_data_in = {w_datain_256[255:128], 128'b0 };
    assign  RAM4_data_in = { 128'b0, w_datain_256[127:0]};
    assign  RAM3_data_in = {w_datain_256[255:128], 128'b0 };
    assign  RAM2_data_in = { 128'b0, w_datain_256[127:0]};
    assign  RAM1_data_in = {w_datain_256[255:128], 128'b0 };
    assign  RAM0_data_in = { 128'b0, w_datain_256[127:0]};

    assign douta = {RAM15_data_out[255:128], RAM14_data_out[127:0], RAM13_data_out[255:128], RAM12_data_out[127:0], RAM11_data_out[255:128], RAM10_data_out[127:0], RAM9_data_out[255:128], RAM8_data_out[127:0], 
                    RAM7_data_out[255:128],  RAM6_data_out[127:0],  RAM5_data_out[255:128],  RAM4_data_out[127:0],  RAM3_data_out[255:128],  RAM2_data_out[127:0],  RAM1_data_out[255:128], RAM0_data_out[127:0]};

    wire [7:0]  w_WEB0_8, w_WEB1_8, w_WEB2_8, w_WEB3_8, w_WEB4_8, w_WEB5_8, w_WEB6_8, w_WEB7_8;
    wire [7:0]  w_WEB8_8, w_WEB9_8, w_WEB10_8, w_WEB11_8, w_WEB12_8, w_WEB13_8, w_WEB14_8, w_WEB15_8;

    // Ƭѡ
    always @( *) begin
        case (addra[2:0])
            3'b000:begin
              w_sel_SRAM_16 = 16'b0000000000000011;
            end
            3'b001:begin
              w_sel_SRAM_16 = 16'b0000000000001100;
            end 
            3'b010:begin
              w_sel_SRAM_16 = 16'b0000000000110000;
            end 
            3'b011:begin
              w_sel_SRAM_16 = 16'b0000000011000000;
            end 
            3'b100:begin
              w_sel_SRAM_16 = 16'b0000001100000000;
            end 
            3'b101:begin
              w_sel_SRAM_16 = 16'b0000110000000000;
            end 
            3'b110:begin
              w_sel_SRAM_16 = 16'b0011000000000000;
            end
            default:begin
              w_sel_SRAM_16 = 16'b1100000000000000;
            end  
            // default:begin
            //   w_sel_SRAM_16 = 16'b0000000000000000;
            // end
        endcase
    end

    assign w_WEB0_8[7:0] = { 8{wea & w_sel_SRAM_16[0]} };
    assign w_WEB1_8[7:0] = { 8{wea & w_sel_SRAM_16[1]} };

    assign w_WEB2_8[7:0] = { 8{wea & w_sel_SRAM_16[2]} };
    assign w_WEB3_8[7:0] = { 8{wea & w_sel_SRAM_16[3]} };

    assign w_WEB4_8[7:0] = { 8{wea & w_sel_SRAM_16[4]} };
    assign w_WEB5_8[7:0] = { 8{wea & w_sel_SRAM_16[5]} };

    assign w_WEB6_8[7:0] = { 8{wea & w_sel_SRAM_16[6]} };
    assign w_WEB7_8[7:0] = { 8{wea & w_sel_SRAM_16[7]} };

    assign w_WEB8_8[7:0] = { 8{wea & w_sel_SRAM_16[8]} };
    assign w_WEB9_8[7:0] = { 8{wea & w_sel_SRAM_16[9]} };

    assign w_WEB10_8[7:0] = { 8{wea & w_sel_SRAM_16[10]} };
    assign w_WEB11_8[7:0] = { 8{wea & w_sel_SRAM_16[11]} };

    assign w_WEB12_8[7:0] = { 8{wea & w_sel_SRAM_16[12]} };
    assign w_WEB13_8[7:0] = { 8{wea & w_sel_SRAM_16[13]} };

    assign w_WEB14_8[7:0] = { 8{wea & w_sel_SRAM_16[14]} };
    assign w_WEB15_8[7:0] = { 8{wea & w_sel_SRAM_16[15]} };

SYKB110_128X16X8CM2 u_L2data0_SYKB110_128X16X8CM2(
    .DO0   (RAM0_data_out[0  ] ),    .DO1   (RAM0_data_out[1  ] ),    .DO2   (RAM0_data_out[2  ] ),    .DO3   (RAM0_data_out[3  ] ),
    .DO4   (RAM0_data_out[4  ] ),    .DO5   (RAM0_data_out[5  ] ),    .DO6   (RAM0_data_out[6  ] ),    .DO7   (RAM0_data_out[7  ] ),
    .DO8   (RAM0_data_out[8  ] ),    .DO9   (RAM0_data_out[9  ] ),    .DO10  (RAM0_data_out[10 ] ),    .DO11  (RAM0_data_out[11 ] ),
    .DO12  (RAM0_data_out[12 ] ),    .DO13  (RAM0_data_out[13 ] ),    .DO14  (RAM0_data_out[14 ] ),    .DO15  (RAM0_data_out[15 ] ),
    .DO16  (RAM0_data_out[16 ] ),    .DO17  (RAM0_data_out[17 ] ),    .DO18  (RAM0_data_out[18 ] ),    .DO19  (RAM0_data_out[19 ] ),
    .DO20  (RAM0_data_out[20 ] ),    .DO21  (RAM0_data_out[21 ] ),    .DO22  (RAM0_data_out[22 ] ),    .DO23  (RAM0_data_out[23 ] ),
    .DO24  (RAM0_data_out[24 ] ),    .DO25  (RAM0_data_out[25 ] ),    .DO26  (RAM0_data_out[26 ] ),    .DO27  (RAM0_data_out[27 ] ),
    .DO28  (RAM0_data_out[28 ] ),    .DO29  (RAM0_data_out[29 ] ),    .DO30  (RAM0_data_out[30 ] ),    .DO31  (RAM0_data_out[31 ] ),
    .DO32  (RAM0_data_out[32 ] ),    .DO33  (RAM0_data_out[33 ] ),    .DO34  (RAM0_data_out[34 ] ),    .DO35  (RAM0_data_out[35 ] ),
    .DO36  (RAM0_data_out[36 ] ),    .DO37  (RAM0_data_out[37 ] ),    .DO38  (RAM0_data_out[38 ] ),    .DO39  (RAM0_data_out[39 ] ),
    .DO40  (RAM0_data_out[40 ] ),    .DO41  (RAM0_data_out[41 ] ),    .DO42  (RAM0_data_out[42 ] ),    .DO43  (RAM0_data_out[43 ] ),
    .DO44  (RAM0_data_out[44 ] ),    .DO45  (RAM0_data_out[45 ] ),    .DO46  (RAM0_data_out[46 ] ),    .DO47  (RAM0_data_out[47 ] ),
    .DO48  (RAM0_data_out[48 ] ),    .DO49  (RAM0_data_out[49 ] ),    .DO50  (RAM0_data_out[50 ] ),    .DO51  (RAM0_data_out[51 ] ),
    .DO52  (RAM0_data_out[52 ] ),    .DO53  (RAM0_data_out[53 ] ),    .DO54  (RAM0_data_out[54 ] ),    .DO55  (RAM0_data_out[55 ] ),
    .DO56  (RAM0_data_out[56 ] ),    .DO57  (RAM0_data_out[57 ] ),    .DO58  (RAM0_data_out[58 ] ),    .DO59  (RAM0_data_out[59 ] ),
    .DO60  (RAM0_data_out[60 ] ),    .DO61  (RAM0_data_out[61 ] ),    .DO62  (RAM0_data_out[62 ] ),    .DO63  (RAM0_data_out[63 ] ),
    .DO64  (RAM0_data_out[64 ] ),    .DO65  (RAM0_data_out[65 ] ),    .DO66  (RAM0_data_out[66 ] ),    .DO67  (RAM0_data_out[67 ] ),
    .DO68  (RAM0_data_out[68 ] ),    .DO69  (RAM0_data_out[69 ] ),    .DO70  (RAM0_data_out[70 ] ),    .DO71  (RAM0_data_out[71 ] ),
    .DO72  (RAM0_data_out[72 ] ),    .DO73  (RAM0_data_out[73 ] ),    .DO74  (RAM0_data_out[74 ] ),    .DO75  (RAM0_data_out[75 ] ),
    .DO76  (RAM0_data_out[76 ] ),    .DO77  (RAM0_data_out[77 ] ),    .DO78  (RAM0_data_out[78 ] ),    .DO79  (RAM0_data_out[79 ] ),
    .DO80  (RAM0_data_out[80 ] ),    .DO81  (RAM0_data_out[81 ] ),    .DO82  (RAM0_data_out[82 ] ),    .DO83  (RAM0_data_out[83 ] ),
    .DO84  (RAM0_data_out[84 ] ),    .DO85  (RAM0_data_out[85 ] ),    .DO86  (RAM0_data_out[86 ] ),    .DO87  (RAM0_data_out[87 ] ),
    .DO88  (RAM0_data_out[88 ] ),    .DO89  (RAM0_data_out[89 ] ),    .DO90  (RAM0_data_out[90 ] ),    .DO91  (RAM0_data_out[91 ] ),
    .DO92  (RAM0_data_out[92 ] ),    .DO93  (RAM0_data_out[93 ] ),    .DO94  (RAM0_data_out[94 ] ),    .DO95  (RAM0_data_out[95 ] ),
    .DO96  (RAM0_data_out[96 ] ),    .DO97  (RAM0_data_out[97 ] ),    .DO98  (RAM0_data_out[98 ] ),    .DO99  (RAM0_data_out[99 ] ),
    .DO100 (RAM0_data_out[100] ),    .DO101 (RAM0_data_out[101] ),    .DO102 (RAM0_data_out[102] ),    .DO103 (RAM0_data_out[103] ),
    .DO104 (RAM0_data_out[104] ),    .DO105 (RAM0_data_out[105] ),    .DO106 (RAM0_data_out[106] ),    .DO107 (RAM0_data_out[107] ),
    .DO108 (RAM0_data_out[108] ),    .DO109 (RAM0_data_out[109] ),    .DO110 (RAM0_data_out[110] ),    .DO111 (RAM0_data_out[111] ),
    .DO112 (RAM0_data_out[112] ),    .DO113 (RAM0_data_out[113] ),    .DO114 (RAM0_data_out[114] ),    .DO115 (RAM0_data_out[115] ),
    .DO116 (RAM0_data_out[116] ),    .DO117 (RAM0_data_out[117] ),    .DO118 (RAM0_data_out[118] ),    .DO119 (RAM0_data_out[119] ),
    .DO120 (RAM0_data_out[120] ),    .DO121 (RAM0_data_out[121] ),    .DO122 (RAM0_data_out[122] ),    .DO123 (RAM0_data_out[123] ),
    .DO124 (RAM0_data_out[124] ),    .DO125 (RAM0_data_out[125] ),    .DO126 (RAM0_data_out[126] ),    .DO127 (RAM0_data_out[127] ),

    .DI0   (RAM0_data_in[0  ] ),    .DI1   (RAM0_data_in[1  ] ),    .DI2   (RAM0_data_in[2  ] ),    .DI3   (RAM0_data_in[3  ] ),
    .DI4   (RAM0_data_in[4  ] ),    .DI5   (RAM0_data_in[5  ] ),    .DI6   (RAM0_data_in[6  ] ),    .DI7   (RAM0_data_in[7  ] ),
    .DI8   (RAM0_data_in[8  ] ),    .DI9   (RAM0_data_in[9  ] ),    .DI10  (RAM0_data_in[10 ] ),    .DI11  (RAM0_data_in[11 ] ),
    .DI12  (RAM0_data_in[12 ] ),    .DI13  (RAM0_data_in[13 ] ),    .DI14  (RAM0_data_in[14 ] ),    .DI15  (RAM0_data_in[15 ] ),
    .DI16  (RAM0_data_in[16 ] ),    .DI17  (RAM0_data_in[17 ] ),    .DI18  (RAM0_data_in[18 ] ),    .DI19  (RAM0_data_in[19 ] ),
    .DI20  (RAM0_data_in[20 ] ),    .DI21  (RAM0_data_in[21 ] ),    .DI22  (RAM0_data_in[22 ] ),    .DI23  (RAM0_data_in[23 ] ),
    .DI24  (RAM0_data_in[24 ] ),    .DI25  (RAM0_data_in[25 ] ),    .DI26  (RAM0_data_in[26 ] ),    .DI27  (RAM0_data_in[27 ] ),
    .DI28  (RAM0_data_in[28 ] ),    .DI29  (RAM0_data_in[29 ] ),    .DI30  (RAM0_data_in[30 ] ),    .DI31  (RAM0_data_in[31 ] ),
    .DI32  (RAM0_data_in[32 ] ),    .DI33  (RAM0_data_in[33 ] ),    .DI34  (RAM0_data_in[34 ] ),    .DI35  (RAM0_data_in[35 ] ),
    .DI36  (RAM0_data_in[36 ] ),    .DI37  (RAM0_data_in[37 ] ),    .DI38  (RAM0_data_in[38 ] ),    .DI39  (RAM0_data_in[39 ] ),
    .DI40  (RAM0_data_in[40 ] ),    .DI41  (RAM0_data_in[41 ] ),    .DI42  (RAM0_data_in[42 ] ),    .DI43  (RAM0_data_in[43 ] ),
    .DI44  (RAM0_data_in[44 ] ),    .DI45  (RAM0_data_in[45 ] ),    .DI46  (RAM0_data_in[46 ] ),    .DI47  (RAM0_data_in[47 ] ),
    .DI48  (RAM0_data_in[48 ] ),    .DI49  (RAM0_data_in[49 ] ),    .DI50  (RAM0_data_in[50 ] ),    .DI51  (RAM0_data_in[51 ] ),
    .DI52  (RAM0_data_in[52 ] ),    .DI53  (RAM0_data_in[53 ] ),    .DI54  (RAM0_data_in[54 ] ),    .DI55  (RAM0_data_in[55 ] ),
    .DI56  (RAM0_data_in[56 ] ),    .DI57  (RAM0_data_in[57 ] ),    .DI58  (RAM0_data_in[58 ] ),    .DI59  (RAM0_data_in[59 ] ),
    .DI60  (RAM0_data_in[60 ] ),    .DI61  (RAM0_data_in[61 ] ),    .DI62  (RAM0_data_in[62 ] ),    .DI63  (RAM0_data_in[63 ] ),
    .DI64  (RAM0_data_in[64 ] ),    .DI65  (RAM0_data_in[65 ] ),    .DI66  (RAM0_data_in[66 ] ),    .DI67  (RAM0_data_in[67 ] ),
    .DI68  (RAM0_data_in[68 ] ),    .DI69  (RAM0_data_in[69 ] ),    .DI70  (RAM0_data_in[70 ] ),    .DI71  (RAM0_data_in[71 ] ),
    .DI72  (RAM0_data_in[72 ] ),    .DI73  (RAM0_data_in[73 ] ),    .DI74  (RAM0_data_in[74 ] ),    .DI75  (RAM0_data_in[75 ] ),
    .DI76  (RAM0_data_in[76 ] ),    .DI77  (RAM0_data_in[77 ] ),    .DI78  (RAM0_data_in[78 ] ),    .DI79  (RAM0_data_in[79 ] ),
    .DI80  (RAM0_data_in[80 ] ),    .DI81  (RAM0_data_in[81 ] ),    .DI82  (RAM0_data_in[82 ] ),    .DI83  (RAM0_data_in[83 ] ),
    .DI84  (RAM0_data_in[84 ] ),    .DI85  (RAM0_data_in[85 ] ),    .DI86  (RAM0_data_in[86 ] ),    .DI87  (RAM0_data_in[87 ] ),
    .DI88  (RAM0_data_in[88 ] ),    .DI89  (RAM0_data_in[89 ] ),    .DI90  (RAM0_data_in[90 ] ),    .DI91  (RAM0_data_in[91 ] ),
    .DI92  (RAM0_data_in[92 ] ),    .DI93  (RAM0_data_in[93 ] ),    .DI94  (RAM0_data_in[94 ] ),    .DI95  (RAM0_data_in[95 ] ),
    .DI96  (RAM0_data_in[96 ] ),    .DI97  (RAM0_data_in[97 ] ),    .DI98  (RAM0_data_in[98 ] ),    .DI99  (RAM0_data_in[99 ] ),
    .DI100 (RAM0_data_in[100] ),    .DI101 (RAM0_data_in[101] ),    .DI102 (RAM0_data_in[102] ),    .DI103 (RAM0_data_in[103] ),
    .DI104 (RAM0_data_in[104] ),    .DI105 (RAM0_data_in[105] ),    .DI106 (RAM0_data_in[106] ),    .DI107 (RAM0_data_in[107] ),
    .DI108 (RAM0_data_in[108] ),    .DI109 (RAM0_data_in[109] ),    .DI110 (RAM0_data_in[110] ),    .DI111 (RAM0_data_in[111] ),
    .DI112 (RAM0_data_in[112] ),    .DI113 (RAM0_data_in[113] ),    .DI114 (RAM0_data_in[114] ),    .DI115 (RAM0_data_in[115] ),
    .DI116 (RAM0_data_in[116] ),    .DI117 (RAM0_data_in[117] ),    .DI118 (RAM0_data_in[118] ),    .DI119 (RAM0_data_in[119] ),
    .DI120 (RAM0_data_in[120] ),    .DI121 (RAM0_data_in[121] ),    .DI122 (RAM0_data_in[122] ),    .DI123 (RAM0_data_in[123] ),
    .DI124 (RAM0_data_in[124] ),    .DI125 (RAM0_data_in[125] ),    .DI126 (RAM0_data_in[126] ),    .DI127 (RAM0_data_in[127] ),

    .A0   (RAM_addr[0]   ),.A1   (RAM_addr[1]   ),.A2   (RAM_addr[2]   ),.A3   (RAM_addr[3]   ),.A4   (RAM_addr[4]   ),.A5   (RAM_addr[5]   ),.A6   (RAM_addr[6]   ),
    .DVSE (1'b0  ),.DVS0 (1'b0  ),.DVS1 (1'b0  ),.DVS2 (1'b0  ),.DVS3 (1'b0  ),
    .WEB0 (~w_WEB0_8[0] ),.WEB1 (~w_WEB0_8[1] ),.WEB2 (~w_WEB0_8[2] ),.WEB3 (~w_WEB0_8[3] ),
    .WEB4 (~w_WEB0_8[4] ),.WEB5 (~w_WEB0_8[5] ),.WEB6 (~w_WEB0_8[6] ),.WEB7 (~w_WEB0_8[7] ),

    .CK    (clka   ),
    .CSB   (1'b0   )
);

SYKB110_128X16X8CM2 u_L2data1_SYKB110_128X16X8CM2(
    .DO0   (RAM1_data_out[128] ),    .DO1   (RAM1_data_out[129] ),    .DO2   (RAM1_data_out[130] ),    .DO3   (RAM1_data_out[131] ),
    .DO4   (RAM1_data_out[132] ),    .DO5   (RAM1_data_out[133] ),    .DO6   (RAM1_data_out[134] ),    .DO7   (RAM1_data_out[135] ),
    .DO8   (RAM1_data_out[136] ),    .DO9   (RAM1_data_out[137] ),    .DO10  (RAM1_data_out[138] ),    .DO11  (RAM1_data_out[139] ),
    .DO12  (RAM1_data_out[140] ),    .DO13  (RAM1_data_out[141] ),    .DO14  (RAM1_data_out[142] ),    .DO15  (RAM1_data_out[143] ),
    .DO16  (RAM1_data_out[144] ),    .DO17  (RAM1_data_out[145] ),    .DO18  (RAM1_data_out[146] ),    .DO19  (RAM1_data_out[147] ),
    .DO20  (RAM1_data_out[148] ),    .DO21  (RAM1_data_out[149] ),    .DO22  (RAM1_data_out[150] ),    .DO23  (RAM1_data_out[151] ),
    .DO24  (RAM1_data_out[152] ),    .DO25  (RAM1_data_out[153] ),    .DO26  (RAM1_data_out[154] ),    .DO27  (RAM1_data_out[155] ),
    .DO28  (RAM1_data_out[156] ),    .DO29  (RAM1_data_out[157] ),    .DO30  (RAM1_data_out[158] ),    .DO31  (RAM1_data_out[159] ),
    .DO32  (RAM1_data_out[160] ),    .DO33  (RAM1_data_out[161] ),    .DO34  (RAM1_data_out[162] ),    .DO35  (RAM1_data_out[163] ),
    .DO36  (RAM1_data_out[164] ),    .DO37  (RAM1_data_out[165] ),    .DO38  (RAM1_data_out[166] ),    .DO39  (RAM1_data_out[167] ),
    .DO40  (RAM1_data_out[168] ),    .DO41  (RAM1_data_out[169] ),    .DO42  (RAM1_data_out[170] ),    .DO43  (RAM1_data_out[171] ),
    .DO44  (RAM1_data_out[172] ),    .DO45  (RAM1_data_out[173] ),    .DO46  (RAM1_data_out[174] ),    .DO47  (RAM1_data_out[175] ),
    .DO48  (RAM1_data_out[176] ),    .DO49  (RAM1_data_out[177] ),    .DO50  (RAM1_data_out[178] ),    .DO51  (RAM1_data_out[179] ),
    .DO52  (RAM1_data_out[180] ),    .DO53  (RAM1_data_out[181] ),    .DO54  (RAM1_data_out[182] ),    .DO55  (RAM1_data_out[183] ),
    .DO56  (RAM1_data_out[184] ),    .DO57  (RAM1_data_out[185] ),    .DO58  (RAM1_data_out[186] ),    .DO59  (RAM1_data_out[187] ),
    .DO60  (RAM1_data_out[188] ),    .DO61  (RAM1_data_out[189] ),    .DO62  (RAM1_data_out[190] ),    .DO63  (RAM1_data_out[191] ),
    .DO64  (RAM1_data_out[192] ),    .DO65  (RAM1_data_out[193] ),    .DO66  (RAM1_data_out[194] ),    .DO67  (RAM1_data_out[195] ),
    .DO68  (RAM1_data_out[196] ),    .DO69  (RAM1_data_out[197] ),    .DO70  (RAM1_data_out[198] ),    .DO71  (RAM1_data_out[199] ),
    .DO72  (RAM1_data_out[200] ),    .DO73  (RAM1_data_out[201] ),    .DO74  (RAM1_data_out[202] ),    .DO75  (RAM1_data_out[203] ),
    .DO76  (RAM1_data_out[204] ),    .DO77  (RAM1_data_out[205] ),    .DO78  (RAM1_data_out[206] ),    .DO79  (RAM1_data_out[207] ),
    .DO80  (RAM1_data_out[208] ),    .DO81  (RAM1_data_out[209] ),    .DO82  (RAM1_data_out[210] ),    .DO83  (RAM1_data_out[211] ),
    .DO84  (RAM1_data_out[212] ),    .DO85  (RAM1_data_out[213] ),    .DO86  (RAM1_data_out[214] ),    .DO87  (RAM1_data_out[215] ),
    .DO88  (RAM1_data_out[216] ),    .DO89  (RAM1_data_out[217] ),    .DO90  (RAM1_data_out[218] ),    .DO91  (RAM1_data_out[219] ),
    .DO92  (RAM1_data_out[220] ),    .DO93  (RAM1_data_out[221] ),    .DO94  (RAM1_data_out[222] ),    .DO95  (RAM1_data_out[223] ),
    .DO96  (RAM1_data_out[224] ),    .DO97  (RAM1_data_out[225] ),    .DO98  (RAM1_data_out[226] ),    .DO99  (RAM1_data_out[227] ),
    .DO100 (RAM1_data_out[228] ),    .DO101 (RAM1_data_out[229] ),    .DO102 (RAM1_data_out[230] ),    .DO103 (RAM1_data_out[231] ),
    .DO104 (RAM1_data_out[232] ),    .DO105 (RAM1_data_out[233] ),    .DO106 (RAM1_data_out[234] ),    .DO107 (RAM1_data_out[235] ),
    .DO108 (RAM1_data_out[236] ),    .DO109 (RAM1_data_out[237] ),    .DO110 (RAM1_data_out[238] ),    .DO111 (RAM1_data_out[239] ),
    .DO112 (RAM1_data_out[240] ),    .DO113 (RAM1_data_out[241] ),    .DO114 (RAM1_data_out[242] ),    .DO115 (RAM1_data_out[243] ),
    .DO116 (RAM1_data_out[244] ),    .DO117 (RAM1_data_out[245] ),    .DO118 (RAM1_data_out[246] ),    .DO119 (RAM1_data_out[247] ),
    .DO120 (RAM1_data_out[248] ),    .DO121 (RAM1_data_out[249] ),    .DO122 (RAM1_data_out[250] ),    .DO123 (RAM1_data_out[251] ),
    .DO124 (RAM1_data_out[252] ),    .DO125 (RAM1_data_out[253] ),    .DO126 (RAM1_data_out[254] ),    .DO127 (RAM1_data_out[255] ),

    .DI0   (RAM1_data_in[128] ),    .DI1   (RAM1_data_in[129] ),    .DI2   (RAM1_data_in[130] ),    .DI3   (RAM1_data_in[131] ),
    .DI4   (RAM1_data_in[132] ),    .DI5   (RAM1_data_in[133] ),    .DI6   (RAM1_data_in[134] ),    .DI7   (RAM1_data_in[135] ),
    .DI8   (RAM1_data_in[136] ),    .DI9   (RAM1_data_in[137] ),    .DI10  (RAM1_data_in[138] ),    .DI11  (RAM1_data_in[139] ),
    .DI12  (RAM1_data_in[140] ),    .DI13  (RAM1_data_in[141] ),    .DI14  (RAM1_data_in[142] ),    .DI15  (RAM1_data_in[143] ),
    .DI16  (RAM1_data_in[144] ),    .DI17  (RAM1_data_in[145] ),    .DI18  (RAM1_data_in[146] ),    .DI19  (RAM1_data_in[147] ),
    .DI20  (RAM1_data_in[148] ),    .DI21  (RAM1_data_in[149] ),    .DI22  (RAM1_data_in[150] ),    .DI23  (RAM1_data_in[151] ),
    .DI24  (RAM1_data_in[152] ),    .DI25  (RAM1_data_in[153] ),    .DI26  (RAM1_data_in[154] ),    .DI27  (RAM1_data_in[155] ),
    .DI28  (RAM1_data_in[156] ),    .DI29  (RAM1_data_in[157] ),    .DI30  (RAM1_data_in[158] ),    .DI31  (RAM1_data_in[159] ),
    .DI32  (RAM1_data_in[160] ),    .DI33  (RAM1_data_in[161] ),    .DI34  (RAM1_data_in[162] ),    .DI35  (RAM1_data_in[163] ),
    .DI36  (RAM1_data_in[164] ),    .DI37  (RAM1_data_in[165] ),    .DI38  (RAM1_data_in[166] ),    .DI39  (RAM1_data_in[167] ),
    .DI40  (RAM1_data_in[168] ),    .DI41  (RAM1_data_in[169] ),    .DI42  (RAM1_data_in[170] ),    .DI43  (RAM1_data_in[171] ),
    .DI44  (RAM1_data_in[172] ),    .DI45  (RAM1_data_in[173] ),    .DI46  (RAM1_data_in[174] ),    .DI47  (RAM1_data_in[175] ),
    .DI48  (RAM1_data_in[176] ),    .DI49  (RAM1_data_in[177] ),    .DI50  (RAM1_data_in[178] ),    .DI51  (RAM1_data_in[179] ),
    .DI52  (RAM1_data_in[180] ),    .DI53  (RAM1_data_in[181] ),    .DI54  (RAM1_data_in[182] ),    .DI55  (RAM1_data_in[183] ),
    .DI56  (RAM1_data_in[184] ),    .DI57  (RAM1_data_in[185] ),    .DI58  (RAM1_data_in[186] ),    .DI59  (RAM1_data_in[187] ),
    .DI60  (RAM1_data_in[188] ),    .DI61  (RAM1_data_in[189] ),    .DI62  (RAM1_data_in[190] ),    .DI63  (RAM1_data_in[191] ),
    .DI64  (RAM1_data_in[192] ),    .DI65  (RAM1_data_in[193] ),    .DI66  (RAM1_data_in[194] ),    .DI67  (RAM1_data_in[195] ),
    .DI68  (RAM1_data_in[196] ),    .DI69  (RAM1_data_in[197] ),    .DI70  (RAM1_data_in[198] ),    .DI71  (RAM1_data_in[199] ),
    .DI72  (RAM1_data_in[200] ),    .DI73  (RAM1_data_in[201] ),    .DI74  (RAM1_data_in[202] ),    .DI75  (RAM1_data_in[203] ),
    .DI76  (RAM1_data_in[204] ),    .DI77  (RAM1_data_in[205] ),    .DI78  (RAM1_data_in[206] ),    .DI79  (RAM1_data_in[207] ),
    .DI80  (RAM1_data_in[208] ),    .DI81  (RAM1_data_in[209] ),    .DI82  (RAM1_data_in[210] ),    .DI83  (RAM1_data_in[211] ),
    .DI84  (RAM1_data_in[212] ),    .DI85  (RAM1_data_in[213] ),    .DI86  (RAM1_data_in[214] ),    .DI87  (RAM1_data_in[215] ),
    .DI88  (RAM1_data_in[216] ),    .DI89  (RAM1_data_in[217] ),    .DI90  (RAM1_data_in[218] ),    .DI91  (RAM1_data_in[219] ),
    .DI92  (RAM1_data_in[220] ),    .DI93  (RAM1_data_in[221] ),    .DI94  (RAM1_data_in[222] ),    .DI95  (RAM1_data_in[223] ),
    .DI96  (RAM1_data_in[224] ),    .DI97  (RAM1_data_in[225] ),    .DI98  (RAM1_data_in[226] ),    .DI99  (RAM1_data_in[227] ),
    .DI100 (RAM1_data_in[228] ),    .DI101 (RAM1_data_in[229] ),    .DI102 (RAM1_data_in[230] ),    .DI103 (RAM1_data_in[231] ),
    .DI104 (RAM1_data_in[232] ),    .DI105 (RAM1_data_in[233] ),    .DI106 (RAM1_data_in[234] ),    .DI107 (RAM1_data_in[235] ),
    .DI108 (RAM1_data_in[236] ),    .DI109 (RAM1_data_in[237] ),    .DI110 (RAM1_data_in[238] ),    .DI111 (RAM1_data_in[239] ),
    .DI112 (RAM1_data_in[240] ),    .DI113 (RAM1_data_in[241] ),    .DI114 (RAM1_data_in[242] ),    .DI115 (RAM1_data_in[243] ),
    .DI116 (RAM1_data_in[244] ),    .DI117 (RAM1_data_in[245] ),    .DI118 (RAM1_data_in[246] ),    .DI119 (RAM1_data_in[247] ),
    .DI120 (RAM1_data_in[248] ),    .DI121 (RAM1_data_in[249] ),    .DI122 (RAM1_data_in[250] ),    .DI123 (RAM1_data_in[251] ),
    .DI124 (RAM1_data_in[252] ),    .DI125 (RAM1_data_in[253] ),    .DI126 (RAM1_data_in[254] ),    .DI127 (RAM1_data_in[255] ),

    .A0   (RAM_addr[0]   ),.A1   (RAM_addr[1]   ),.A2   (RAM_addr[2]   ),.A3   (RAM_addr[3]   ),.A4   (RAM_addr[4]   ),.A5   (RAM_addr[5]   ),.A6   (RAM_addr[6]   ),
    .DVSE (1'b0  ),.DVS0 (1'b0  ),.DVS1 (1'b0  ),.DVS2 (1'b0  ),.DVS3 (1'b0  ),
    .WEB0 (~w_WEB1_8[0] ),.WEB1 (~w_WEB1_8[1] ),.WEB2 (~w_WEB1_8[2] ),.WEB3 (~w_WEB1_8[3] ),
    .WEB4 (~w_WEB1_8[4] ),.WEB5 (~w_WEB1_8[5] ),.WEB6 (~w_WEB1_8[6] ),.WEB7 (~w_WEB1_8[7] ),

    .CK    (clka   ),
    .CSB   (1'b0   )
);


SYKB110_128X16X8CM2 u_L2data2_SYKB110_128X16X8CM2(
    .DO0   (RAM2_data_out[0  ] ),    .DO1   (RAM2_data_out[1  ] ),    .DO2   (RAM2_data_out[2  ] ),    .DO3   (RAM2_data_out[3  ] ),
    .DO4   (RAM2_data_out[4  ] ),    .DO5   (RAM2_data_out[5  ] ),    .DO6   (RAM2_data_out[6  ] ),    .DO7   (RAM2_data_out[7  ] ),
    .DO8   (RAM2_data_out[8  ] ),    .DO9   (RAM2_data_out[9  ] ),    .DO10  (RAM2_data_out[10 ] ),    .DO11  (RAM2_data_out[11 ] ),
    .DO12  (RAM2_data_out[12 ] ),    .DO13  (RAM2_data_out[13 ] ),    .DO14  (RAM2_data_out[14 ] ),    .DO15  (RAM2_data_out[15 ] ),
    .DO16  (RAM2_data_out[16 ] ),    .DO17  (RAM2_data_out[17 ] ),    .DO18  (RAM2_data_out[18 ] ),    .DO19  (RAM2_data_out[19 ] ),
    .DO20  (RAM2_data_out[20 ] ),    .DO21  (RAM2_data_out[21 ] ),    .DO22  (RAM2_data_out[22 ] ),    .DO23  (RAM2_data_out[23 ] ),
    .DO24  (RAM2_data_out[24 ] ),    .DO25  (RAM2_data_out[25 ] ),    .DO26  (RAM2_data_out[26 ] ),    .DO27  (RAM2_data_out[27 ] ),
    .DO28  (RAM2_data_out[28 ] ),    .DO29  (RAM2_data_out[29 ] ),    .DO30  (RAM2_data_out[30 ] ),    .DO31  (RAM2_data_out[31 ] ),
    .DO32  (RAM2_data_out[32 ] ),    .DO33  (RAM2_data_out[33 ] ),    .DO34  (RAM2_data_out[34 ] ),    .DO35  (RAM2_data_out[35 ] ),
    .DO36  (RAM2_data_out[36 ] ),    .DO37  (RAM2_data_out[37 ] ),    .DO38  (RAM2_data_out[38 ] ),    .DO39  (RAM2_data_out[39 ] ),
    .DO40  (RAM2_data_out[40 ] ),    .DO41  (RAM2_data_out[41 ] ),    .DO42  (RAM2_data_out[42 ] ),    .DO43  (RAM2_data_out[43 ] ),
    .DO44  (RAM2_data_out[44 ] ),    .DO45  (RAM2_data_out[45 ] ),    .DO46  (RAM2_data_out[46 ] ),    .DO47  (RAM2_data_out[47 ] ),
    .DO48  (RAM2_data_out[48 ] ),    .DO49  (RAM2_data_out[49 ] ),    .DO50  (RAM2_data_out[50 ] ),    .DO51  (RAM2_data_out[51 ] ),
    .DO52  (RAM2_data_out[52 ] ),    .DO53  (RAM2_data_out[53 ] ),    .DO54  (RAM2_data_out[54 ] ),    .DO55  (RAM2_data_out[55 ] ),
    .DO56  (RAM2_data_out[56 ] ),    .DO57  (RAM2_data_out[57 ] ),    .DO58  (RAM2_data_out[58 ] ),    .DO59  (RAM2_data_out[59 ] ),
    .DO60  (RAM2_data_out[60 ] ),    .DO61  (RAM2_data_out[61 ] ),    .DO62  (RAM2_data_out[62 ] ),    .DO63  (RAM2_data_out[63 ] ),
    .DO64  (RAM2_data_out[64 ] ),    .DO65  (RAM2_data_out[65 ] ),    .DO66  (RAM2_data_out[66 ] ),    .DO67  (RAM2_data_out[67 ] ),
    .DO68  (RAM2_data_out[68 ] ),    .DO69  (RAM2_data_out[69 ] ),    .DO70  (RAM2_data_out[70 ] ),    .DO71  (RAM2_data_out[71 ] ),
    .DO72  (RAM2_data_out[72 ] ),    .DO73  (RAM2_data_out[73 ] ),    .DO74  (RAM2_data_out[74 ] ),    .DO75  (RAM2_data_out[75 ] ),
    .DO76  (RAM2_data_out[76 ] ),    .DO77  (RAM2_data_out[77 ] ),    .DO78  (RAM2_data_out[78 ] ),    .DO79  (RAM2_data_out[79 ] ),
    .DO80  (RAM2_data_out[80 ] ),    .DO81  (RAM2_data_out[81 ] ),    .DO82  (RAM2_data_out[82 ] ),    .DO83  (RAM2_data_out[83 ] ),
    .DO84  (RAM2_data_out[84 ] ),    .DO85  (RAM2_data_out[85 ] ),    .DO86  (RAM2_data_out[86 ] ),    .DO87  (RAM2_data_out[87 ] ),
    .DO88  (RAM2_data_out[88 ] ),    .DO89  (RAM2_data_out[89 ] ),    .DO90  (RAM2_data_out[90 ] ),    .DO91  (RAM2_data_out[91 ] ),
    .DO92  (RAM2_data_out[92 ] ),    .DO93  (RAM2_data_out[93 ] ),    .DO94  (RAM2_data_out[94 ] ),    .DO95  (RAM2_data_out[95 ] ),
    .DO96  (RAM2_data_out[96 ] ),    .DO97  (RAM2_data_out[97 ] ),    .DO98  (RAM2_data_out[98 ] ),    .DO99  (RAM2_data_out[99 ] ),
    .DO100 (RAM2_data_out[100] ),    .DO101 (RAM2_data_out[101] ),    .DO102 (RAM2_data_out[102] ),    .DO103 (RAM2_data_out[103] ),
    .DO104 (RAM2_data_out[104] ),    .DO105 (RAM2_data_out[105] ),    .DO106 (RAM2_data_out[106] ),    .DO107 (RAM2_data_out[107] ),
    .DO108 (RAM2_data_out[108] ),    .DO109 (RAM2_data_out[109] ),    .DO110 (RAM2_data_out[110] ),    .DO111 (RAM2_data_out[111] ),
    .DO112 (RAM2_data_out[112] ),    .DO113 (RAM2_data_out[113] ),    .DO114 (RAM2_data_out[114] ),    .DO115 (RAM2_data_out[115] ),
    .DO116 (RAM2_data_out[116] ),    .DO117 (RAM2_data_out[117] ),    .DO118 (RAM2_data_out[118] ),    .DO119 (RAM2_data_out[119] ),
    .DO120 (RAM2_data_out[120] ),    .DO121 (RAM2_data_out[121] ),    .DO122 (RAM2_data_out[122] ),    .DO123 (RAM2_data_out[123] ),
    .DO124 (RAM2_data_out[124] ),    .DO125 (RAM2_data_out[125] ),    .DO126 (RAM2_data_out[126] ),    .DO127 (RAM2_data_out[127] ),

    .DI0   (RAM2_data_in[0  ] ),    .DI1   (RAM2_data_in[1  ] ),    .DI2   (RAM2_data_in[2  ] ),    .DI3   (RAM2_data_in[3  ] ),
    .DI4   (RAM2_data_in[4  ] ),    .DI5   (RAM2_data_in[5  ] ),    .DI6   (RAM2_data_in[6  ] ),    .DI7   (RAM2_data_in[7  ] ),
    .DI8   (RAM2_data_in[8  ] ),    .DI9   (RAM2_data_in[9  ] ),    .DI10  (RAM2_data_in[10 ] ),    .DI11  (RAM2_data_in[11 ] ),
    .DI12  (RAM2_data_in[12 ] ),    .DI13  (RAM2_data_in[13 ] ),    .DI14  (RAM2_data_in[14 ] ),    .DI15  (RAM2_data_in[15 ] ),
    .DI16  (RAM2_data_in[16 ] ),    .DI17  (RAM2_data_in[17 ] ),    .DI18  (RAM2_data_in[18 ] ),    .DI19  (RAM2_data_in[19 ] ),
    .DI20  (RAM2_data_in[20 ] ),    .DI21  (RAM2_data_in[21 ] ),    .DI22  (RAM2_data_in[22 ] ),    .DI23  (RAM2_data_in[23 ] ),
    .DI24  (RAM2_data_in[24 ] ),    .DI25  (RAM2_data_in[25 ] ),    .DI26  (RAM2_data_in[26 ] ),    .DI27  (RAM2_data_in[27 ] ),
    .DI28  (RAM2_data_in[28 ] ),    .DI29  (RAM2_data_in[29 ] ),    .DI30  (RAM2_data_in[30 ] ),    .DI31  (RAM2_data_in[31 ] ),
    .DI32  (RAM2_data_in[32 ] ),    .DI33  (RAM2_data_in[33 ] ),    .DI34  (RAM2_data_in[34 ] ),    .DI35  (RAM2_data_in[35 ] ),
    .DI36  (RAM2_data_in[36 ] ),    .DI37  (RAM2_data_in[37 ] ),    .DI38  (RAM2_data_in[38 ] ),    .DI39  (RAM2_data_in[39 ] ),
    .DI40  (RAM2_data_in[40 ] ),    .DI41  (RAM2_data_in[41 ] ),    .DI42  (RAM2_data_in[42 ] ),    .DI43  (RAM2_data_in[43 ] ),
    .DI44  (RAM2_data_in[44 ] ),    .DI45  (RAM2_data_in[45 ] ),    .DI46  (RAM2_data_in[46 ] ),    .DI47  (RAM2_data_in[47 ] ),
    .DI48  (RAM2_data_in[48 ] ),    .DI49  (RAM2_data_in[49 ] ),    .DI50  (RAM2_data_in[50 ] ),    .DI51  (RAM2_data_in[51 ] ),
    .DI52  (RAM2_data_in[52 ] ),    .DI53  (RAM2_data_in[53 ] ),    .DI54  (RAM2_data_in[54 ] ),    .DI55  (RAM2_data_in[55 ] ),
    .DI56  (RAM2_data_in[56 ] ),    .DI57  (RAM2_data_in[57 ] ),    .DI58  (RAM2_data_in[58 ] ),    .DI59  (RAM2_data_in[59 ] ),
    .DI60  (RAM2_data_in[60 ] ),    .DI61  (RAM2_data_in[61 ] ),    .DI62  (RAM2_data_in[62 ] ),    .DI63  (RAM2_data_in[63 ] ),
    .DI64  (RAM2_data_in[64 ] ),    .DI65  (RAM2_data_in[65 ] ),    .DI66  (RAM2_data_in[66 ] ),    .DI67  (RAM2_data_in[67 ] ),
    .DI68  (RAM2_data_in[68 ] ),    .DI69  (RAM2_data_in[69 ] ),    .DI70  (RAM2_data_in[70 ] ),    .DI71  (RAM2_data_in[71 ] ),
    .DI72  (RAM2_data_in[72 ] ),    .DI73  (RAM2_data_in[73 ] ),    .DI74  (RAM2_data_in[74 ] ),    .DI75  (RAM2_data_in[75 ] ),
    .DI76  (RAM2_data_in[76 ] ),    .DI77  (RAM2_data_in[77 ] ),    .DI78  (RAM2_data_in[78 ] ),    .DI79  (RAM2_data_in[79 ] ),
    .DI80  (RAM2_data_in[80 ] ),    .DI81  (RAM2_data_in[81 ] ),    .DI82  (RAM2_data_in[82 ] ),    .DI83  (RAM2_data_in[83 ] ),
    .DI84  (RAM2_data_in[84 ] ),    .DI85  (RAM2_data_in[85 ] ),    .DI86  (RAM2_data_in[86 ] ),    .DI87  (RAM2_data_in[87 ] ),
    .DI88  (RAM2_data_in[88 ] ),    .DI89  (RAM2_data_in[89 ] ),    .DI90  (RAM2_data_in[90 ] ),    .DI91  (RAM2_data_in[91 ] ),
    .DI92  (RAM2_data_in[92 ] ),    .DI93  (RAM2_data_in[93 ] ),    .DI94  (RAM2_data_in[94 ] ),    .DI95  (RAM2_data_in[95 ] ),
    .DI96  (RAM2_data_in[96 ] ),    .DI97  (RAM2_data_in[97 ] ),    .DI98  (RAM2_data_in[98 ] ),    .DI99  (RAM2_data_in[99 ] ),
    .DI100 (RAM2_data_in[100] ),    .DI101 (RAM2_data_in[101] ),    .DI102 (RAM2_data_in[102] ),    .DI103 (RAM2_data_in[103] ),
    .DI104 (RAM2_data_in[104] ),    .DI105 (RAM2_data_in[105] ),    .DI106 (RAM2_data_in[106] ),    .DI107 (RAM2_data_in[107] ),
    .DI108 (RAM2_data_in[108] ),    .DI109 (RAM2_data_in[109] ),    .DI110 (RAM2_data_in[110] ),    .DI111 (RAM2_data_in[111] ),
    .DI112 (RAM2_data_in[112] ),    .DI113 (RAM2_data_in[113] ),    .DI114 (RAM2_data_in[114] ),    .DI115 (RAM2_data_in[115] ),
    .DI116 (RAM2_data_in[116] ),    .DI117 (RAM2_data_in[117] ),    .DI118 (RAM2_data_in[118] ),    .DI119 (RAM2_data_in[119] ),
    .DI120 (RAM2_data_in[120] ),    .DI121 (RAM2_data_in[121] ),    .DI122 (RAM2_data_in[122] ),    .DI123 (RAM2_data_in[123] ),
    .DI124 (RAM2_data_in[124] ),    .DI125 (RAM2_data_in[125] ),    .DI126 (RAM2_data_in[126] ),    .DI127 (RAM2_data_in[127] ),

    .A0   (RAM_addr[0]   ),.A1   (RAM_addr[1]   ),.A2   (RAM_addr[2]   ),.A3   (RAM_addr[3]   ),.A4   (RAM_addr[4]   ),.A5   (RAM_addr[5]   ),.A6   (RAM_addr[6]   ),
    .DVSE (1'b0  ),.DVS0 (1'b0  ),.DVS1 (1'b0  ),.DVS2 (1'b0  ),.DVS3 (1'b0  ),
    .WEB0 (~w_WEB2_8[0] ),.WEB1 (~w_WEB2_8[1] ),.WEB2 (~w_WEB2_8[2] ),.WEB3 (~w_WEB2_8[3] ),
    .WEB4 (~w_WEB2_8[4] ),.WEB5 (~w_WEB2_8[5] ),.WEB6 (~w_WEB2_8[6] ),.WEB7 (~w_WEB2_8[7] ),

    .CK    (clka   ),
    .CSB   (1'b0   )
);


SYKB110_128X16X8CM2 u_L2data3_SYKB110_128X16X8CM2(
    .DO0   (RAM3_data_out[128] ),    .DO1   (RAM3_data_out[129] ),    .DO2   (RAM3_data_out[130] ),    .DO3   (RAM3_data_out[131] ),
    .DO4   (RAM3_data_out[132] ),    .DO5   (RAM3_data_out[133] ),    .DO6   (RAM3_data_out[134] ),    .DO7   (RAM3_data_out[135] ),
    .DO8   (RAM3_data_out[136] ),    .DO9   (RAM3_data_out[137] ),    .DO10  (RAM3_data_out[138] ),    .DO11  (RAM3_data_out[139] ),
    .DO12  (RAM3_data_out[140] ),    .DO13  (RAM3_data_out[141] ),    .DO14  (RAM3_data_out[142] ),    .DO15  (RAM3_data_out[143] ),
    .DO16  (RAM3_data_out[144] ),    .DO17  (RAM3_data_out[145] ),    .DO18  (RAM3_data_out[146] ),    .DO19  (RAM3_data_out[147] ),
    .DO20  (RAM3_data_out[148] ),    .DO21  (RAM3_data_out[149] ),    .DO22  (RAM3_data_out[150] ),    .DO23  (RAM3_data_out[151] ),
    .DO24  (RAM3_data_out[152] ),    .DO25  (RAM3_data_out[153] ),    .DO26  (RAM3_data_out[154] ),    .DO27  (RAM3_data_out[155] ),
    .DO28  (RAM3_data_out[156] ),    .DO29  (RAM3_data_out[157] ),    .DO30  (RAM3_data_out[158] ),    .DO31  (RAM3_data_out[159] ),
    .DO32  (RAM3_data_out[160] ),    .DO33  (RAM3_data_out[161] ),    .DO34  (RAM3_data_out[162] ),    .DO35  (RAM3_data_out[163] ),
    .DO36  (RAM3_data_out[164] ),    .DO37  (RAM3_data_out[165] ),    .DO38  (RAM3_data_out[166] ),    .DO39  (RAM3_data_out[167] ),
    .DO40  (RAM3_data_out[168] ),    .DO41  (RAM3_data_out[169] ),    .DO42  (RAM3_data_out[170] ),    .DO43  (RAM3_data_out[171] ),
    .DO44  (RAM3_data_out[172] ),    .DO45  (RAM3_data_out[173] ),    .DO46  (RAM3_data_out[174] ),    .DO47  (RAM3_data_out[175] ),
    .DO48  (RAM3_data_out[176] ),    .DO49  (RAM3_data_out[177] ),    .DO50  (RAM3_data_out[178] ),    .DO51  (RAM3_data_out[179] ),
    .DO52  (RAM3_data_out[180] ),    .DO53  (RAM3_data_out[181] ),    .DO54  (RAM3_data_out[182] ),    .DO55  (RAM3_data_out[183] ),
    .DO56  (RAM3_data_out[184] ),    .DO57  (RAM3_data_out[185] ),    .DO58  (RAM3_data_out[186] ),    .DO59  (RAM3_data_out[187] ),
    .DO60  (RAM3_data_out[188] ),    .DO61  (RAM3_data_out[189] ),    .DO62  (RAM3_data_out[190] ),    .DO63  (RAM3_data_out[191] ),
    .DO64  (RAM3_data_out[192] ),    .DO65  (RAM3_data_out[193] ),    .DO66  (RAM3_data_out[194] ),    .DO67  (RAM3_data_out[195] ),
    .DO68  (RAM3_data_out[196] ),    .DO69  (RAM3_data_out[197] ),    .DO70  (RAM3_data_out[198] ),    .DO71  (RAM3_data_out[199] ),
    .DO72  (RAM3_data_out[200] ),    .DO73  (RAM3_data_out[201] ),    .DO74  (RAM3_data_out[202] ),    .DO75  (RAM3_data_out[203] ),
    .DO76  (RAM3_data_out[204] ),    .DO77  (RAM3_data_out[205] ),    .DO78  (RAM3_data_out[206] ),    .DO79  (RAM3_data_out[207] ),
    .DO80  (RAM3_data_out[208] ),    .DO81  (RAM3_data_out[209] ),    .DO82  (RAM3_data_out[210] ),    .DO83  (RAM3_data_out[211] ),
    .DO84  (RAM3_data_out[212] ),    .DO85  (RAM3_data_out[213] ),    .DO86  (RAM3_data_out[214] ),    .DO87  (RAM3_data_out[215] ),
    .DO88  (RAM3_data_out[216] ),    .DO89  (RAM3_data_out[217] ),    .DO90  (RAM3_data_out[218] ),    .DO91  (RAM3_data_out[219] ),
    .DO92  (RAM3_data_out[220] ),    .DO93  (RAM3_data_out[221] ),    .DO94  (RAM3_data_out[222] ),    .DO95  (RAM3_data_out[223] ),
    .DO96  (RAM3_data_out[224] ),    .DO97  (RAM3_data_out[225] ),    .DO98  (RAM3_data_out[226] ),    .DO99  (RAM3_data_out[227] ),
    .DO100 (RAM3_data_out[228] ),    .DO101 (RAM3_data_out[229] ),    .DO102 (RAM3_data_out[230] ),    .DO103 (RAM3_data_out[231] ),
    .DO104 (RAM3_data_out[232] ),    .DO105 (RAM3_data_out[233] ),    .DO106 (RAM3_data_out[234] ),    .DO107 (RAM3_data_out[235] ),
    .DO108 (RAM3_data_out[236] ),    .DO109 (RAM3_data_out[237] ),    .DO110 (RAM3_data_out[238] ),    .DO111 (RAM3_data_out[239] ),
    .DO112 (RAM3_data_out[240] ),    .DO113 (RAM3_data_out[241] ),    .DO114 (RAM3_data_out[242] ),    .DO115 (RAM3_data_out[243] ),
    .DO116 (RAM3_data_out[244] ),    .DO117 (RAM3_data_out[245] ),    .DO118 (RAM3_data_out[246] ),    .DO119 (RAM3_data_out[247] ),
    .DO120 (RAM3_data_out[248] ),    .DO121 (RAM3_data_out[249] ),    .DO122 (RAM3_data_out[250] ),    .DO123 (RAM3_data_out[251] ),
    .DO124 (RAM3_data_out[252] ),    .DO125 (RAM3_data_out[253] ),    .DO126 (RAM3_data_out[254] ),    .DO127 (RAM3_data_out[255] ),

    .DI0   (RAM3_data_in[128] ),    .DI1   (RAM3_data_in[129] ),    .DI2   (RAM3_data_in[130] ),    .DI3   (RAM3_data_in[131] ),
    .DI4   (RAM3_data_in[132] ),    .DI5   (RAM3_data_in[133] ),    .DI6   (RAM3_data_in[134] ),    .DI7   (RAM3_data_in[135] ),
    .DI8   (RAM3_data_in[136] ),    .DI9   (RAM3_data_in[137] ),    .DI10  (RAM3_data_in[138] ),    .DI11  (RAM3_data_in[139] ),
    .DI12  (RAM3_data_in[140] ),    .DI13  (RAM3_data_in[141] ),    .DI14  (RAM3_data_in[142] ),    .DI15  (RAM3_data_in[143] ),
    .DI16  (RAM3_data_in[144] ),    .DI17  (RAM3_data_in[145] ),    .DI18  (RAM3_data_in[146] ),    .DI19  (RAM3_data_in[147] ),
    .DI20  (RAM3_data_in[148] ),    .DI21  (RAM3_data_in[149] ),    .DI22  (RAM3_data_in[150] ),    .DI23  (RAM3_data_in[151] ),
    .DI24  (RAM3_data_in[152] ),    .DI25  (RAM3_data_in[153] ),    .DI26  (RAM3_data_in[154] ),    .DI27  (RAM3_data_in[155] ),
    .DI28  (RAM3_data_in[156] ),    .DI29  (RAM3_data_in[157] ),    .DI30  (RAM3_data_in[158] ),    .DI31  (RAM3_data_in[159] ),
    .DI32  (RAM3_data_in[160] ),    .DI33  (RAM3_data_in[161] ),    .DI34  (RAM3_data_in[162] ),    .DI35  (RAM3_data_in[163] ),
    .DI36  (RAM3_data_in[164] ),    .DI37  (RAM3_data_in[165] ),    .DI38  (RAM3_data_in[166] ),    .DI39  (RAM3_data_in[167] ),
    .DI40  (RAM3_data_in[168] ),    .DI41  (RAM3_data_in[169] ),    .DI42  (RAM3_data_in[170] ),    .DI43  (RAM3_data_in[171] ),
    .DI44  (RAM3_data_in[172] ),    .DI45  (RAM3_data_in[173] ),    .DI46  (RAM3_data_in[174] ),    .DI47  (RAM3_data_in[175] ),
    .DI48  (RAM3_data_in[176] ),    .DI49  (RAM3_data_in[177] ),    .DI50  (RAM3_data_in[178] ),    .DI51  (RAM3_data_in[179] ),
    .DI52  (RAM3_data_in[180] ),    .DI53  (RAM3_data_in[181] ),    .DI54  (RAM3_data_in[182] ),    .DI55  (RAM3_data_in[183] ),
    .DI56  (RAM3_data_in[184] ),    .DI57  (RAM3_data_in[185] ),    .DI58  (RAM3_data_in[186] ),    .DI59  (RAM3_data_in[187] ),
    .DI60  (RAM3_data_in[188] ),    .DI61  (RAM3_data_in[189] ),    .DI62  (RAM3_data_in[190] ),    .DI63  (RAM3_data_in[191] ),
    .DI64  (RAM3_data_in[192] ),    .DI65  (RAM3_data_in[193] ),    .DI66  (RAM3_data_in[194] ),    .DI67  (RAM3_data_in[195] ),
    .DI68  (RAM3_data_in[196] ),    .DI69  (RAM3_data_in[197] ),    .DI70  (RAM3_data_in[198] ),    .DI71  (RAM3_data_in[199] ),
    .DI72  (RAM3_data_in[200] ),    .DI73  (RAM3_data_in[201] ),    .DI74  (RAM3_data_in[202] ),    .DI75  (RAM3_data_in[203] ),
    .DI76  (RAM3_data_in[204] ),    .DI77  (RAM3_data_in[205] ),    .DI78  (RAM3_data_in[206] ),    .DI79  (RAM3_data_in[207] ),
    .DI80  (RAM3_data_in[208] ),    .DI81  (RAM3_data_in[209] ),    .DI82  (RAM3_data_in[210] ),    .DI83  (RAM3_data_in[211] ),
    .DI84  (RAM3_data_in[212] ),    .DI85  (RAM3_data_in[213] ),    .DI86  (RAM3_data_in[214] ),    .DI87  (RAM3_data_in[215] ),
    .DI88  (RAM3_data_in[216] ),    .DI89  (RAM3_data_in[217] ),    .DI90  (RAM3_data_in[218] ),    .DI91  (RAM3_data_in[219] ),
    .DI92  (RAM3_data_in[220] ),    .DI93  (RAM3_data_in[221] ),    .DI94  (RAM3_data_in[222] ),    .DI95  (RAM3_data_in[223] ),
    .DI96  (RAM3_data_in[224] ),    .DI97  (RAM3_data_in[225] ),    .DI98  (RAM3_data_in[226] ),    .DI99  (RAM3_data_in[227] ),
    .DI100 (RAM3_data_in[228] ),    .DI101 (RAM3_data_in[229] ),    .DI102 (RAM3_data_in[230] ),    .DI103 (RAM3_data_in[231] ),
    .DI104 (RAM3_data_in[232] ),    .DI105 (RAM3_data_in[233] ),    .DI106 (RAM3_data_in[234] ),    .DI107 (RAM3_data_in[235] ),
    .DI108 (RAM3_data_in[236] ),    .DI109 (RAM3_data_in[237] ),    .DI110 (RAM3_data_in[238] ),    .DI111 (RAM3_data_in[239] ),
    .DI112 (RAM3_data_in[240] ),    .DI113 (RAM3_data_in[241] ),    .DI114 (RAM3_data_in[242] ),    .DI115 (RAM3_data_in[243] ),
    .DI116 (RAM3_data_in[244] ),    .DI117 (RAM3_data_in[245] ),    .DI118 (RAM3_data_in[246] ),    .DI119 (RAM3_data_in[247] ),
    .DI120 (RAM3_data_in[248] ),    .DI121 (RAM3_data_in[249] ),    .DI122 (RAM3_data_in[250] ),    .DI123 (RAM3_data_in[251] ),
    .DI124 (RAM3_data_in[252] ),    .DI125 (RAM3_data_in[253] ),    .DI126 (RAM3_data_in[254] ),    .DI127 (RAM3_data_in[255] ),

    .A0   (RAM_addr[0]   ),.A1   (RAM_addr[1]   ),.A2   (RAM_addr[2]   ),.A3   (RAM_addr[3]   ),.A4   (RAM_addr[4]   ),.A5   (RAM_addr[5]   ),.A6   (RAM_addr[6]   ),
    .DVSE (1'b0  ),.DVS0 (1'b0  ),.DVS1 (1'b0  ),.DVS2 (1'b0  ),.DVS3 (1'b0  ),
    .WEB0 (~w_WEB3_8[0] ),.WEB1 (~w_WEB3_8[1] ),.WEB2 (~w_WEB3_8[2] ),.WEB3 (~w_WEB3_8[3] ),
    .WEB4 (~w_WEB3_8[4] ),.WEB5 (~w_WEB3_8[5] ),.WEB6 (~w_WEB3_8[6] ),.WEB7 (~w_WEB3_8[7] ),

    .CK    (clka   ),
    .CSB   (1'b0   )
);

    
SYKB110_128X16X8CM2 u_L2data4_SYKB110_128X16X8CM2(
    .DO0   (RAM4_data_out[0  ] ),    .DO1   (RAM4_data_out[1  ] ),    .DO2   (RAM4_data_out[2  ] ),    .DO3   (RAM4_data_out[3  ] ),
    .DO4   (RAM4_data_out[4  ] ),    .DO5   (RAM4_data_out[5  ] ),    .DO6   (RAM4_data_out[6  ] ),    .DO7   (RAM4_data_out[7  ] ),
    .DO8   (RAM4_data_out[8  ] ),    .DO9   (RAM4_data_out[9  ] ),    .DO10  (RAM4_data_out[10 ] ),    .DO11  (RAM4_data_out[11 ] ),
    .DO12  (RAM4_data_out[12 ] ),    .DO13  (RAM4_data_out[13 ] ),    .DO14  (RAM4_data_out[14 ] ),    .DO15  (RAM4_data_out[15 ] ),
    .DO16  (RAM4_data_out[16 ] ),    .DO17  (RAM4_data_out[17 ] ),    .DO18  (RAM4_data_out[18 ] ),    .DO19  (RAM4_data_out[19 ] ),
    .DO20  (RAM4_data_out[20 ] ),    .DO21  (RAM4_data_out[21 ] ),    .DO22  (RAM4_data_out[22 ] ),    .DO23  (RAM4_data_out[23 ] ),
    .DO24  (RAM4_data_out[24 ] ),    .DO25  (RAM4_data_out[25 ] ),    .DO26  (RAM4_data_out[26 ] ),    .DO27  (RAM4_data_out[27 ] ),
    .DO28  (RAM4_data_out[28 ] ),    .DO29  (RAM4_data_out[29 ] ),    .DO30  (RAM4_data_out[30 ] ),    .DO31  (RAM4_data_out[31 ] ),
    .DO32  (RAM4_data_out[32 ] ),    .DO33  (RAM4_data_out[33 ] ),    .DO34  (RAM4_data_out[34 ] ),    .DO35  (RAM4_data_out[35 ] ),
    .DO36  (RAM4_data_out[36 ] ),    .DO37  (RAM4_data_out[37 ] ),    .DO38  (RAM4_data_out[38 ] ),    .DO39  (RAM4_data_out[39 ] ),
    .DO40  (RAM4_data_out[40 ] ),    .DO41  (RAM4_data_out[41 ] ),    .DO42  (RAM4_data_out[42 ] ),    .DO43  (RAM4_data_out[43 ] ),
    .DO44  (RAM4_data_out[44 ] ),    .DO45  (RAM4_data_out[45 ] ),    .DO46  (RAM4_data_out[46 ] ),    .DO47  (RAM4_data_out[47 ] ),
    .DO48  (RAM4_data_out[48 ] ),    .DO49  (RAM4_data_out[49 ] ),    .DO50  (RAM4_data_out[50 ] ),    .DO51  (RAM4_data_out[51 ] ),
    .DO52  (RAM4_data_out[52 ] ),    .DO53  (RAM4_data_out[53 ] ),    .DO54  (RAM4_data_out[54 ] ),    .DO55  (RAM4_data_out[55 ] ),
    .DO56  (RAM4_data_out[56 ] ),    .DO57  (RAM4_data_out[57 ] ),    .DO58  (RAM4_data_out[58 ] ),    .DO59  (RAM4_data_out[59 ] ),
    .DO60  (RAM4_data_out[60 ] ),    .DO61  (RAM4_data_out[61 ] ),    .DO62  (RAM4_data_out[62 ] ),    .DO63  (RAM4_data_out[63 ] ),
    .DO64  (RAM4_data_out[64 ] ),    .DO65  (RAM4_data_out[65 ] ),    .DO66  (RAM4_data_out[66 ] ),    .DO67  (RAM4_data_out[67 ] ),
    .DO68  (RAM4_data_out[68 ] ),    .DO69  (RAM4_data_out[69 ] ),    .DO70  (RAM4_data_out[70 ] ),    .DO71  (RAM4_data_out[71 ] ),
    .DO72  (RAM4_data_out[72 ] ),    .DO73  (RAM4_data_out[73 ] ),    .DO74  (RAM4_data_out[74 ] ),    .DO75  (RAM4_data_out[75 ] ),
    .DO76  (RAM4_data_out[76 ] ),    .DO77  (RAM4_data_out[77 ] ),    .DO78  (RAM4_data_out[78 ] ),    .DO79  (RAM4_data_out[79 ] ),
    .DO80  (RAM4_data_out[80 ] ),    .DO81  (RAM4_data_out[81 ] ),    .DO82  (RAM4_data_out[82 ] ),    .DO83  (RAM4_data_out[83 ] ),
    .DO84  (RAM4_data_out[84 ] ),    .DO85  (RAM4_data_out[85 ] ),    .DO86  (RAM4_data_out[86 ] ),    .DO87  (RAM4_data_out[87 ] ),
    .DO88  (RAM4_data_out[88 ] ),    .DO89  (RAM4_data_out[89 ] ),    .DO90  (RAM4_data_out[90 ] ),    .DO91  (RAM4_data_out[91 ] ),
    .DO92  (RAM4_data_out[92 ] ),    .DO93  (RAM4_data_out[93 ] ),    .DO94  (RAM4_data_out[94 ] ),    .DO95  (RAM4_data_out[95 ] ),
    .DO96  (RAM4_data_out[96 ] ),    .DO97  (RAM4_data_out[97 ] ),    .DO98  (RAM4_data_out[98 ] ),    .DO99  (RAM4_data_out[99 ] ),
    .DO100 (RAM4_data_out[100] ),    .DO101 (RAM4_data_out[101] ),    .DO102 (RAM4_data_out[102] ),    .DO103 (RAM4_data_out[103] ),
    .DO104 (RAM4_data_out[104] ),    .DO105 (RAM4_data_out[105] ),    .DO106 (RAM4_data_out[106] ),    .DO107 (RAM4_data_out[107] ),
    .DO108 (RAM4_data_out[108] ),    .DO109 (RAM4_data_out[109] ),    .DO110 (RAM4_data_out[110] ),    .DO111 (RAM4_data_out[111] ),
    .DO112 (RAM4_data_out[112] ),    .DO113 (RAM4_data_out[113] ),    .DO114 (RAM4_data_out[114] ),    .DO115 (RAM4_data_out[115] ),
    .DO116 (RAM4_data_out[116] ),    .DO117 (RAM4_data_out[117] ),    .DO118 (RAM4_data_out[118] ),    .DO119 (RAM4_data_out[119] ),
    .DO120 (RAM4_data_out[120] ),    .DO121 (RAM4_data_out[121] ),    .DO122 (RAM4_data_out[122] ),    .DO123 (RAM4_data_out[123] ),
    .DO124 (RAM4_data_out[124] ),    .DO125 (RAM4_data_out[125] ),    .DO126 (RAM4_data_out[126] ),    .DO127 (RAM4_data_out[127] ),

    .DI0   (RAM4_data_in[0  ] ),    .DI1   (RAM4_data_in[1  ] ),    .DI2   (RAM4_data_in[2  ] ),    .DI3   (RAM4_data_in[3  ] ),
    .DI4   (RAM4_data_in[4  ] ),    .DI5   (RAM4_data_in[5  ] ),    .DI6   (RAM4_data_in[6  ] ),    .DI7   (RAM4_data_in[7  ] ),
    .DI8   (RAM4_data_in[8  ] ),    .DI9   (RAM4_data_in[9  ] ),    .DI10  (RAM4_data_in[10 ] ),    .DI11  (RAM4_data_in[11 ] ),
    .DI12  (RAM4_data_in[12 ] ),    .DI13  (RAM4_data_in[13 ] ),    .DI14  (RAM4_data_in[14 ] ),    .DI15  (RAM4_data_in[15 ] ),
    .DI16  (RAM4_data_in[16 ] ),    .DI17  (RAM4_data_in[17 ] ),    .DI18  (RAM4_data_in[18 ] ),    .DI19  (RAM4_data_in[19 ] ),
    .DI20  (RAM4_data_in[20 ] ),    .DI21  (RAM4_data_in[21 ] ),    .DI22  (RAM4_data_in[22 ] ),    .DI23  (RAM4_data_in[23 ] ),
    .DI24  (RAM4_data_in[24 ] ),    .DI25  (RAM4_data_in[25 ] ),    .DI26  (RAM4_data_in[26 ] ),    .DI27  (RAM4_data_in[27 ] ),
    .DI28  (RAM4_data_in[28 ] ),    .DI29  (RAM4_data_in[29 ] ),    .DI30  (RAM4_data_in[30 ] ),    .DI31  (RAM4_data_in[31 ] ),
    .DI32  (RAM4_data_in[32 ] ),    .DI33  (RAM4_data_in[33 ] ),    .DI34  (RAM4_data_in[34 ] ),    .DI35  (RAM4_data_in[35 ] ),
    .DI36  (RAM4_data_in[36 ] ),    .DI37  (RAM4_data_in[37 ] ),    .DI38  (RAM4_data_in[38 ] ),    .DI39  (RAM4_data_in[39 ] ),
    .DI40  (RAM4_data_in[40 ] ),    .DI41  (RAM4_data_in[41 ] ),    .DI42  (RAM4_data_in[42 ] ),    .DI43  (RAM4_data_in[43 ] ),
    .DI44  (RAM4_data_in[44 ] ),    .DI45  (RAM4_data_in[45 ] ),    .DI46  (RAM4_data_in[46 ] ),    .DI47  (RAM4_data_in[47 ] ),
    .DI48  (RAM4_data_in[48 ] ),    .DI49  (RAM4_data_in[49 ] ),    .DI50  (RAM4_data_in[50 ] ),    .DI51  (RAM4_data_in[51 ] ),
    .DI52  (RAM4_data_in[52 ] ),    .DI53  (RAM4_data_in[53 ] ),    .DI54  (RAM4_data_in[54 ] ),    .DI55  (RAM4_data_in[55 ] ),
    .DI56  (RAM4_data_in[56 ] ),    .DI57  (RAM4_data_in[57 ] ),    .DI58  (RAM4_data_in[58 ] ),    .DI59  (RAM4_data_in[59 ] ),
    .DI60  (RAM4_data_in[60 ] ),    .DI61  (RAM4_data_in[61 ] ),    .DI62  (RAM4_data_in[62 ] ),    .DI63  (RAM4_data_in[63 ] ),
    .DI64  (RAM4_data_in[64 ] ),    .DI65  (RAM4_data_in[65 ] ),    .DI66  (RAM4_data_in[66 ] ),    .DI67  (RAM4_data_in[67 ] ),
    .DI68  (RAM4_data_in[68 ] ),    .DI69  (RAM4_data_in[69 ] ),    .DI70  (RAM4_data_in[70 ] ),    .DI71  (RAM4_data_in[71 ] ),
    .DI72  (RAM4_data_in[72 ] ),    .DI73  (RAM4_data_in[73 ] ),    .DI74  (RAM4_data_in[74 ] ),    .DI75  (RAM4_data_in[75 ] ),
    .DI76  (RAM4_data_in[76 ] ),    .DI77  (RAM4_data_in[77 ] ),    .DI78  (RAM4_data_in[78 ] ),    .DI79  (RAM4_data_in[79 ] ),
    .DI80  (RAM4_data_in[80 ] ),    .DI81  (RAM4_data_in[81 ] ),    .DI82  (RAM4_data_in[82 ] ),    .DI83  (RAM4_data_in[83 ] ),
    .DI84  (RAM4_data_in[84 ] ),    .DI85  (RAM4_data_in[85 ] ),    .DI86  (RAM4_data_in[86 ] ),    .DI87  (RAM4_data_in[87 ] ),
    .DI88  (RAM4_data_in[88 ] ),    .DI89  (RAM4_data_in[89 ] ),    .DI90  (RAM4_data_in[90 ] ),    .DI91  (RAM4_data_in[91 ] ),
    .DI92  (RAM4_data_in[92 ] ),    .DI93  (RAM4_data_in[93 ] ),    .DI94  (RAM4_data_in[94 ] ),    .DI95  (RAM4_data_in[95 ] ),
    .DI96  (RAM4_data_in[96 ] ),    .DI97  (RAM4_data_in[97 ] ),    .DI98  (RAM4_data_in[98 ] ),    .DI99  (RAM4_data_in[99 ] ),
    .DI100 (RAM4_data_in[100] ),    .DI101 (RAM4_data_in[101] ),    .DI102 (RAM4_data_in[102] ),    .DI103 (RAM4_data_in[103] ),
    .DI104 (RAM4_data_in[104] ),    .DI105 (RAM4_data_in[105] ),    .DI106 (RAM4_data_in[106] ),    .DI107 (RAM4_data_in[107] ),
    .DI108 (RAM4_data_in[108] ),    .DI109 (RAM4_data_in[109] ),    .DI110 (RAM4_data_in[110] ),    .DI111 (RAM4_data_in[111] ),
    .DI112 (RAM4_data_in[112] ),    .DI113 (RAM4_data_in[113] ),    .DI114 (RAM4_data_in[114] ),    .DI115 (RAM4_data_in[115] ),
    .DI116 (RAM4_data_in[116] ),    .DI117 (RAM4_data_in[117] ),    .DI118 (RAM4_data_in[118] ),    .DI119 (RAM4_data_in[119] ),
    .DI120 (RAM4_data_in[120] ),    .DI121 (RAM4_data_in[121] ),    .DI122 (RAM4_data_in[122] ),    .DI123 (RAM4_data_in[123] ),
    .DI124 (RAM4_data_in[124] ),    .DI125 (RAM4_data_in[125] ),    .DI126 (RAM4_data_in[126] ),    .DI127 (RAM4_data_in[127] ),

    .A0   (RAM_addr[0]   ),.A1   (RAM_addr[1]   ),.A2   (RAM_addr[2]   ),.A3   (RAM_addr[3]   ),.A4   (RAM_addr[4]   ),.A5   (RAM_addr[5]   ),.A6   (RAM_addr[6]   ),
    .DVSE (1'b0  ),.DVS0 (1'b0  ),.DVS1 (1'b0  ),.DVS2 (1'b0  ),.DVS3 (1'b0  ),
    .WEB0 (~w_WEB4_8[0] ),.WEB1 (~w_WEB4_8[1] ),.WEB2 (~w_WEB4_8[2] ),.WEB3 (~w_WEB4_8[3] ),
    .WEB4 (~w_WEB4_8[4] ),.WEB5 (~w_WEB4_8[5] ),.WEB6 (~w_WEB4_8[6] ),.WEB7 (~w_WEB4_8[7] ),

    .CK    (clka   ),
    .CSB   (1'b0   )
);


SYKB110_128X16X8CM2 u_L2data5_SYKB110_128X16X8CM2(
    .DO0   (RAM5_data_out[128] ),    .DO1   (RAM5_data_out[129] ),    .DO2   (RAM5_data_out[130] ),    .DO3   (RAM5_data_out[131] ),
    .DO4   (RAM5_data_out[132] ),    .DO5   (RAM5_data_out[133] ),    .DO6   (RAM5_data_out[134] ),    .DO7   (RAM5_data_out[135] ),
    .DO8   (RAM5_data_out[136] ),    .DO9   (RAM5_data_out[137] ),    .DO10  (RAM5_data_out[138] ),    .DO11  (RAM5_data_out[139] ),
    .DO12  (RAM5_data_out[140] ),    .DO13  (RAM5_data_out[141] ),    .DO14  (RAM5_data_out[142] ),    .DO15  (RAM5_data_out[143] ),
    .DO16  (RAM5_data_out[144] ),    .DO17  (RAM5_data_out[145] ),    .DO18  (RAM5_data_out[146] ),    .DO19  (RAM5_data_out[147] ),
    .DO20  (RAM5_data_out[148] ),    .DO21  (RAM5_data_out[149] ),    .DO22  (RAM5_data_out[150] ),    .DO23  (RAM5_data_out[151] ),
    .DO24  (RAM5_data_out[152] ),    .DO25  (RAM5_data_out[153] ),    .DO26  (RAM5_data_out[154] ),    .DO27  (RAM5_data_out[155] ),
    .DO28  (RAM5_data_out[156] ),    .DO29  (RAM5_data_out[157] ),    .DO30  (RAM5_data_out[158] ),    .DO31  (RAM5_data_out[159] ),
    .DO32  (RAM5_data_out[160] ),    .DO33  (RAM5_data_out[161] ),    .DO34  (RAM5_data_out[162] ),    .DO35  (RAM5_data_out[163] ),
    .DO36  (RAM5_data_out[164] ),    .DO37  (RAM5_data_out[165] ),    .DO38  (RAM5_data_out[166] ),    .DO39  (RAM5_data_out[167] ),
    .DO40  (RAM5_data_out[168] ),    .DO41  (RAM5_data_out[169] ),    .DO42  (RAM5_data_out[170] ),    .DO43  (RAM5_data_out[171] ),
    .DO44  (RAM5_data_out[172] ),    .DO45  (RAM5_data_out[173] ),    .DO46  (RAM5_data_out[174] ),    .DO47  (RAM5_data_out[175] ),
    .DO48  (RAM5_data_out[176] ),    .DO49  (RAM5_data_out[177] ),    .DO50  (RAM5_data_out[178] ),    .DO51  (RAM5_data_out[179] ),
    .DO52  (RAM5_data_out[180] ),    .DO53  (RAM5_data_out[181] ),    .DO54  (RAM5_data_out[182] ),    .DO55  (RAM5_data_out[183] ),
    .DO56  (RAM5_data_out[184] ),    .DO57  (RAM5_data_out[185] ),    .DO58  (RAM5_data_out[186] ),    .DO59  (RAM5_data_out[187] ),
    .DO60  (RAM5_data_out[188] ),    .DO61  (RAM5_data_out[189] ),    .DO62  (RAM5_data_out[190] ),    .DO63  (RAM5_data_out[191] ),
    .DO64  (RAM5_data_out[192] ),    .DO65  (RAM5_data_out[193] ),    .DO66  (RAM5_data_out[194] ),    .DO67  (RAM5_data_out[195] ),
    .DO68  (RAM5_data_out[196] ),    .DO69  (RAM5_data_out[197] ),    .DO70  (RAM5_data_out[198] ),    .DO71  (RAM5_data_out[199] ),
    .DO72  (RAM5_data_out[200] ),    .DO73  (RAM5_data_out[201] ),    .DO74  (RAM5_data_out[202] ),    .DO75  (RAM5_data_out[203] ),
    .DO76  (RAM5_data_out[204] ),    .DO77  (RAM5_data_out[205] ),    .DO78  (RAM5_data_out[206] ),    .DO79  (RAM5_data_out[207] ),
    .DO80  (RAM5_data_out[208] ),    .DO81  (RAM5_data_out[209] ),    .DO82  (RAM5_data_out[210] ),    .DO83  (RAM5_data_out[211] ),
    .DO84  (RAM5_data_out[212] ),    .DO85  (RAM5_data_out[213] ),    .DO86  (RAM5_data_out[214] ),    .DO87  (RAM5_data_out[215] ),
    .DO88  (RAM5_data_out[216] ),    .DO89  (RAM5_data_out[217] ),    .DO90  (RAM5_data_out[218] ),    .DO91  (RAM5_data_out[219] ),
    .DO92  (RAM5_data_out[220] ),    .DO93  (RAM5_data_out[221] ),    .DO94  (RAM5_data_out[222] ),    .DO95  (RAM5_data_out[223] ),
    .DO96  (RAM5_data_out[224] ),    .DO97  (RAM5_data_out[225] ),    .DO98  (RAM5_data_out[226] ),    .DO99  (RAM5_data_out[227] ),
    .DO100 (RAM5_data_out[228] ),    .DO101 (RAM5_data_out[229] ),    .DO102 (RAM5_data_out[230] ),    .DO103 (RAM5_data_out[231] ),
    .DO104 (RAM5_data_out[232] ),    .DO105 (RAM5_data_out[233] ),    .DO106 (RAM5_data_out[234] ),    .DO107 (RAM5_data_out[235] ),
    .DO108 (RAM5_data_out[236] ),    .DO109 (RAM5_data_out[237] ),    .DO110 (RAM5_data_out[238] ),    .DO111 (RAM5_data_out[239] ),
    .DO112 (RAM5_data_out[240] ),    .DO113 (RAM5_data_out[241] ),    .DO114 (RAM5_data_out[242] ),    .DO115 (RAM5_data_out[243] ),
    .DO116 (RAM5_data_out[244] ),    .DO117 (RAM5_data_out[245] ),    .DO118 (RAM5_data_out[246] ),    .DO119 (RAM5_data_out[247] ),
    .DO120 (RAM5_data_out[248] ),    .DO121 (RAM5_data_out[249] ),    .DO122 (RAM5_data_out[250] ),    .DO123 (RAM5_data_out[251] ),
    .DO124 (RAM5_data_out[252] ),    .DO125 (RAM5_data_out[253] ),    .DO126 (RAM5_data_out[254] ),    .DO127 (RAM5_data_out[255] ),

    .DI0   (RAM5_data_in[128] ),    .DI1   (RAM5_data_in[129] ),    .DI2   (RAM5_data_in[130] ),    .DI3   (RAM5_data_in[131] ),
    .DI4   (RAM5_data_in[132] ),    .DI5   (RAM5_data_in[133] ),    .DI6   (RAM5_data_in[134] ),    .DI7   (RAM5_data_in[135] ),
    .DI8   (RAM5_data_in[136] ),    .DI9   (RAM5_data_in[137] ),    .DI10  (RAM5_data_in[138] ),    .DI11  (RAM5_data_in[139] ),
    .DI12  (RAM5_data_in[140] ),    .DI13  (RAM5_data_in[141] ),    .DI14  (RAM5_data_in[142] ),    .DI15  (RAM5_data_in[143] ),
    .DI16  (RAM5_data_in[144] ),    .DI17  (RAM5_data_in[145] ),    .DI18  (RAM5_data_in[146] ),    .DI19  (RAM5_data_in[147] ),
    .DI20  (RAM5_data_in[148] ),    .DI21  (RAM5_data_in[149] ),    .DI22  (RAM5_data_in[150] ),    .DI23  (RAM5_data_in[151] ),
    .DI24  (RAM5_data_in[152] ),    .DI25  (RAM5_data_in[153] ),    .DI26  (RAM5_data_in[154] ),    .DI27  (RAM5_data_in[155] ),
    .DI28  (RAM5_data_in[156] ),    .DI29  (RAM5_data_in[157] ),    .DI30  (RAM5_data_in[158] ),    .DI31  (RAM5_data_in[159] ),
    .DI32  (RAM5_data_in[160] ),    .DI33  (RAM5_data_in[161] ),    .DI34  (RAM5_data_in[162] ),    .DI35  (RAM5_data_in[163] ),
    .DI36  (RAM5_data_in[164] ),    .DI37  (RAM5_data_in[165] ),    .DI38  (RAM5_data_in[166] ),    .DI39  (RAM5_data_in[167] ),
    .DI40  (RAM5_data_in[168] ),    .DI41  (RAM5_data_in[169] ),    .DI42  (RAM5_data_in[170] ),    .DI43  (RAM5_data_in[171] ),
    .DI44  (RAM5_data_in[172] ),    .DI45  (RAM5_data_in[173] ),    .DI46  (RAM5_data_in[174] ),    .DI47  (RAM5_data_in[175] ),
    .DI48  (RAM5_data_in[176] ),    .DI49  (RAM5_data_in[177] ),    .DI50  (RAM5_data_in[178] ),    .DI51  (RAM5_data_in[179] ),
    .DI52  (RAM5_data_in[180] ),    .DI53  (RAM5_data_in[181] ),    .DI54  (RAM5_data_in[182] ),    .DI55  (RAM5_data_in[183] ),
    .DI56  (RAM5_data_in[184] ),    .DI57  (RAM5_data_in[185] ),    .DI58  (RAM5_data_in[186] ),    .DI59  (RAM5_data_in[187] ),
    .DI60  (RAM5_data_in[188] ),    .DI61  (RAM5_data_in[189] ),    .DI62  (RAM5_data_in[190] ),    .DI63  (RAM5_data_in[191] ),
    .DI64  (RAM5_data_in[192] ),    .DI65  (RAM5_data_in[193] ),    .DI66  (RAM5_data_in[194] ),    .DI67  (RAM5_data_in[195] ),
    .DI68  (RAM5_data_in[196] ),    .DI69  (RAM5_data_in[197] ),    .DI70  (RAM5_data_in[198] ),    .DI71  (RAM5_data_in[199] ),
    .DI72  (RAM5_data_in[200] ),    .DI73  (RAM5_data_in[201] ),    .DI74  (RAM5_data_in[202] ),    .DI75  (RAM5_data_in[203] ),
    .DI76  (RAM5_data_in[204] ),    .DI77  (RAM5_data_in[205] ),    .DI78  (RAM5_data_in[206] ),    .DI79  (RAM5_data_in[207] ),
    .DI80  (RAM5_data_in[208] ),    .DI81  (RAM5_data_in[209] ),    .DI82  (RAM5_data_in[210] ),    .DI83  (RAM5_data_in[211] ),
    .DI84  (RAM5_data_in[212] ),    .DI85  (RAM5_data_in[213] ),    .DI86  (RAM5_data_in[214] ),    .DI87  (RAM5_data_in[215] ),
    .DI88  (RAM5_data_in[216] ),    .DI89  (RAM5_data_in[217] ),    .DI90  (RAM5_data_in[218] ),    .DI91  (RAM5_data_in[219] ),
    .DI92  (RAM5_data_in[220] ),    .DI93  (RAM5_data_in[221] ),    .DI94  (RAM5_data_in[222] ),    .DI95  (RAM5_data_in[223] ),
    .DI96  (RAM5_data_in[224] ),    .DI97  (RAM5_data_in[225] ),    .DI98  (RAM5_data_in[226] ),    .DI99  (RAM5_data_in[227] ),
    .DI100 (RAM5_data_in[228] ),    .DI101 (RAM5_data_in[229] ),    .DI102 (RAM5_data_in[230] ),    .DI103 (RAM5_data_in[231] ),
    .DI104 (RAM5_data_in[232] ),    .DI105 (RAM5_data_in[233] ),    .DI106 (RAM5_data_in[234] ),    .DI107 (RAM5_data_in[235] ),
    .DI108 (RAM5_data_in[236] ),    .DI109 (RAM5_data_in[237] ),    .DI110 (RAM5_data_in[238] ),    .DI111 (RAM5_data_in[239] ),
    .DI112 (RAM5_data_in[240] ),    .DI113 (RAM5_data_in[241] ),    .DI114 (RAM5_data_in[242] ),    .DI115 (RAM5_data_in[243] ),
    .DI116 (RAM5_data_in[244] ),    .DI117 (RAM5_data_in[245] ),    .DI118 (RAM5_data_in[246] ),    .DI119 (RAM5_data_in[247] ),
    .DI120 (RAM5_data_in[248] ),    .DI121 (RAM5_data_in[249] ),    .DI122 (RAM5_data_in[250] ),    .DI123 (RAM5_data_in[251] ),
    .DI124 (RAM5_data_in[252] ),    .DI125 (RAM5_data_in[253] ),    .DI126 (RAM5_data_in[254] ),    .DI127 (RAM5_data_in[255] ),

    .A0   (RAM_addr[0]   ),.A1   (RAM_addr[1]   ),.A2   (RAM_addr[2]   ),.A3   (RAM_addr[3]   ),.A4   (RAM_addr[4]   ),.A5   (RAM_addr[5]   ),.A6   (RAM_addr[6]   ),
    .DVSE (1'b0  ),.DVS0 (1'b0  ),.DVS1 (1'b0  ),.DVS2 (1'b0  ),.DVS3 (1'b0  ),
    .WEB0 (~w_WEB5_8[0] ),.WEB1 (~w_WEB5_8[1] ),.WEB2 (~w_WEB5_8[2] ),.WEB3 (~w_WEB5_8[3] ),
    .WEB4 (~w_WEB5_8[4] ),.WEB5 (~w_WEB5_8[5] ),.WEB6 (~w_WEB5_8[6] ),.WEB7 (~w_WEB5_8[7] ),

    .CK    (clka   ),
    .CSB   (1'b0   )
);


SYKB110_128X16X8CM2 u_L2data6_SYKB110_128X16X8CM2(
    .DO0   (RAM6_data_out[0  ] ),    .DO1   (RAM6_data_out[1  ] ),    .DO2   (RAM6_data_out[2  ] ),    .DO3   (RAM6_data_out[3  ] ),
    .DO4   (RAM6_data_out[4  ] ),    .DO5   (RAM6_data_out[5  ] ),    .DO6   (RAM6_data_out[6  ] ),    .DO7   (RAM6_data_out[7  ] ),
    .DO8   (RAM6_data_out[8  ] ),    .DO9   (RAM6_data_out[9  ] ),    .DO10  (RAM6_data_out[10 ] ),    .DO11  (RAM6_data_out[11 ] ),
    .DO12  (RAM6_data_out[12 ] ),    .DO13  (RAM6_data_out[13 ] ),    .DO14  (RAM6_data_out[14 ] ),    .DO15  (RAM6_data_out[15 ] ),
    .DO16  (RAM6_data_out[16 ] ),    .DO17  (RAM6_data_out[17 ] ),    .DO18  (RAM6_data_out[18 ] ),    .DO19  (RAM6_data_out[19 ] ),
    .DO20  (RAM6_data_out[20 ] ),    .DO21  (RAM6_data_out[21 ] ),    .DO22  (RAM6_data_out[22 ] ),    .DO23  (RAM6_data_out[23 ] ),
    .DO24  (RAM6_data_out[24 ] ),    .DO25  (RAM6_data_out[25 ] ),    .DO26  (RAM6_data_out[26 ] ),    .DO27  (RAM6_data_out[27 ] ),
    .DO28  (RAM6_data_out[28 ] ),    .DO29  (RAM6_data_out[29 ] ),    .DO30  (RAM6_data_out[30 ] ),    .DO31  (RAM6_data_out[31 ] ),
    .DO32  (RAM6_data_out[32 ] ),    .DO33  (RAM6_data_out[33 ] ),    .DO34  (RAM6_data_out[34 ] ),    .DO35  (RAM6_data_out[35 ] ),
    .DO36  (RAM6_data_out[36 ] ),    .DO37  (RAM6_data_out[37 ] ),    .DO38  (RAM6_data_out[38 ] ),    .DO39  (RAM6_data_out[39 ] ),
    .DO40  (RAM6_data_out[40 ] ),    .DO41  (RAM6_data_out[41 ] ),    .DO42  (RAM6_data_out[42 ] ),    .DO43  (RAM6_data_out[43 ] ),
    .DO44  (RAM6_data_out[44 ] ),    .DO45  (RAM6_data_out[45 ] ),    .DO46  (RAM6_data_out[46 ] ),    .DO47  (RAM6_data_out[47 ] ),
    .DO48  (RAM6_data_out[48 ] ),    .DO49  (RAM6_data_out[49 ] ),    .DO50  (RAM6_data_out[50 ] ),    .DO51  (RAM6_data_out[51 ] ),
    .DO52  (RAM6_data_out[52 ] ),    .DO53  (RAM6_data_out[53 ] ),    .DO54  (RAM6_data_out[54 ] ),    .DO55  (RAM6_data_out[55 ] ),
    .DO56  (RAM6_data_out[56 ] ),    .DO57  (RAM6_data_out[57 ] ),    .DO58  (RAM6_data_out[58 ] ),    .DO59  (RAM6_data_out[59 ] ),
    .DO60  (RAM6_data_out[60 ] ),    .DO61  (RAM6_data_out[61 ] ),    .DO62  (RAM6_data_out[62 ] ),    .DO63  (RAM6_data_out[63 ] ),
    .DO64  (RAM6_data_out[64 ] ),    .DO65  (RAM6_data_out[65 ] ),    .DO66  (RAM6_data_out[66 ] ),    .DO67  (RAM6_data_out[67 ] ),
    .DO68  (RAM6_data_out[68 ] ),    .DO69  (RAM6_data_out[69 ] ),    .DO70  (RAM6_data_out[70 ] ),    .DO71  (RAM6_data_out[71 ] ),
    .DO72  (RAM6_data_out[72 ] ),    .DO73  (RAM6_data_out[73 ] ),    .DO74  (RAM6_data_out[74 ] ),    .DO75  (RAM6_data_out[75 ] ),
    .DO76  (RAM6_data_out[76 ] ),    .DO77  (RAM6_data_out[77 ] ),    .DO78  (RAM6_data_out[78 ] ),    .DO79  (RAM6_data_out[79 ] ),
    .DO80  (RAM6_data_out[80 ] ),    .DO81  (RAM6_data_out[81 ] ),    .DO82  (RAM6_data_out[82 ] ),    .DO83  (RAM6_data_out[83 ] ),
    .DO84  (RAM6_data_out[84 ] ),    .DO85  (RAM6_data_out[85 ] ),    .DO86  (RAM6_data_out[86 ] ),    .DO87  (RAM6_data_out[87 ] ),
    .DO88  (RAM6_data_out[88 ] ),    .DO89  (RAM6_data_out[89 ] ),    .DO90  (RAM6_data_out[90 ] ),    .DO91  (RAM6_data_out[91 ] ),
    .DO92  (RAM6_data_out[92 ] ),    .DO93  (RAM6_data_out[93 ] ),    .DO94  (RAM6_data_out[94 ] ),    .DO95  (RAM6_data_out[95 ] ),
    .DO96  (RAM6_data_out[96 ] ),    .DO97  (RAM6_data_out[97 ] ),    .DO98  (RAM6_data_out[98 ] ),    .DO99  (RAM6_data_out[99 ] ),
    .DO100 (RAM6_data_out[100] ),    .DO101 (RAM6_data_out[101] ),    .DO102 (RAM6_data_out[102] ),    .DO103 (RAM6_data_out[103] ),
    .DO104 (RAM6_data_out[104] ),    .DO105 (RAM6_data_out[105] ),    .DO106 (RAM6_data_out[106] ),    .DO107 (RAM6_data_out[107] ),
    .DO108 (RAM6_data_out[108] ),    .DO109 (RAM6_data_out[109] ),    .DO110 (RAM6_data_out[110] ),    .DO111 (RAM6_data_out[111] ),
    .DO112 (RAM6_data_out[112] ),    .DO113 (RAM6_data_out[113] ),    .DO114 (RAM6_data_out[114] ),    .DO115 (RAM6_data_out[115] ),
    .DO116 (RAM6_data_out[116] ),    .DO117 (RAM6_data_out[117] ),    .DO118 (RAM6_data_out[118] ),    .DO119 (RAM6_data_out[119] ),
    .DO120 (RAM6_data_out[120] ),    .DO121 (RAM6_data_out[121] ),    .DO122 (RAM6_data_out[122] ),    .DO123 (RAM6_data_out[123] ),
    .DO124 (RAM6_data_out[124] ),    .DO125 (RAM6_data_out[125] ),    .DO126 (RAM6_data_out[126] ),    .DO127 (RAM6_data_out[127] ),

    .DI0   (RAM6_data_in[0  ] ),    .DI1   (RAM6_data_in[1  ] ),    .DI2   (RAM6_data_in[2  ] ),    .DI3   (RAM6_data_in[3  ] ),
    .DI4   (RAM6_data_in[4  ] ),    .DI5   (RAM6_data_in[5  ] ),    .DI6   (RAM6_data_in[6  ] ),    .DI7   (RAM6_data_in[7  ] ),
    .DI8   (RAM6_data_in[8  ] ),    .DI9   (RAM6_data_in[9  ] ),    .DI10  (RAM6_data_in[10 ] ),    .DI11  (RAM6_data_in[11 ] ),
    .DI12  (RAM6_data_in[12 ] ),    .DI13  (RAM6_data_in[13 ] ),    .DI14  (RAM6_data_in[14 ] ),    .DI15  (RAM6_data_in[15 ] ),
    .DI16  (RAM6_data_in[16 ] ),    .DI17  (RAM6_data_in[17 ] ),    .DI18  (RAM6_data_in[18 ] ),    .DI19  (RAM6_data_in[19 ] ),
    .DI20  (RAM6_data_in[20 ] ),    .DI21  (RAM6_data_in[21 ] ),    .DI22  (RAM6_data_in[22 ] ),    .DI23  (RAM6_data_in[23 ] ),
    .DI24  (RAM6_data_in[24 ] ),    .DI25  (RAM6_data_in[25 ] ),    .DI26  (RAM6_data_in[26 ] ),    .DI27  (RAM6_data_in[27 ] ),
    .DI28  (RAM6_data_in[28 ] ),    .DI29  (RAM6_data_in[29 ] ),    .DI30  (RAM6_data_in[30 ] ),    .DI31  (RAM6_data_in[31 ] ),
    .DI32  (RAM6_data_in[32 ] ),    .DI33  (RAM6_data_in[33 ] ),    .DI34  (RAM6_data_in[34 ] ),    .DI35  (RAM6_data_in[35 ] ),
    .DI36  (RAM6_data_in[36 ] ),    .DI37  (RAM6_data_in[37 ] ),    .DI38  (RAM6_data_in[38 ] ),    .DI39  (RAM6_data_in[39 ] ),
    .DI40  (RAM6_data_in[40 ] ),    .DI41  (RAM6_data_in[41 ] ),    .DI42  (RAM6_data_in[42 ] ),    .DI43  (RAM6_data_in[43 ] ),
    .DI44  (RAM6_data_in[44 ] ),    .DI45  (RAM6_data_in[45 ] ),    .DI46  (RAM6_data_in[46 ] ),    .DI47  (RAM6_data_in[47 ] ),
    .DI48  (RAM6_data_in[48 ] ),    .DI49  (RAM6_data_in[49 ] ),    .DI50  (RAM6_data_in[50 ] ),    .DI51  (RAM6_data_in[51 ] ),
    .DI52  (RAM6_data_in[52 ] ),    .DI53  (RAM6_data_in[53 ] ),    .DI54  (RAM6_data_in[54 ] ),    .DI55  (RAM6_data_in[55 ] ),
    .DI56  (RAM6_data_in[56 ] ),    .DI57  (RAM6_data_in[57 ] ),    .DI58  (RAM6_data_in[58 ] ),    .DI59  (RAM6_data_in[59 ] ),
    .DI60  (RAM6_data_in[60 ] ),    .DI61  (RAM6_data_in[61 ] ),    .DI62  (RAM6_data_in[62 ] ),    .DI63  (RAM6_data_in[63 ] ),
    .DI64  (RAM6_data_in[64 ] ),    .DI65  (RAM6_data_in[65 ] ),    .DI66  (RAM6_data_in[66 ] ),    .DI67  (RAM6_data_in[67 ] ),
    .DI68  (RAM6_data_in[68 ] ),    .DI69  (RAM6_data_in[69 ] ),    .DI70  (RAM6_data_in[70 ] ),    .DI71  (RAM6_data_in[71 ] ),
    .DI72  (RAM6_data_in[72 ] ),    .DI73  (RAM6_data_in[73 ] ),    .DI74  (RAM6_data_in[74 ] ),    .DI75  (RAM6_data_in[75 ] ),
    .DI76  (RAM6_data_in[76 ] ),    .DI77  (RAM6_data_in[77 ] ),    .DI78  (RAM6_data_in[78 ] ),    .DI79  (RAM6_data_in[79 ] ),
    .DI80  (RAM6_data_in[80 ] ),    .DI81  (RAM6_data_in[81 ] ),    .DI82  (RAM6_data_in[82 ] ),    .DI83  (RAM6_data_in[83 ] ),
    .DI84  (RAM6_data_in[84 ] ),    .DI85  (RAM6_data_in[85 ] ),    .DI86  (RAM6_data_in[86 ] ),    .DI87  (RAM6_data_in[87 ] ),
    .DI88  (RAM6_data_in[88 ] ),    .DI89  (RAM6_data_in[89 ] ),    .DI90  (RAM6_data_in[90 ] ),    .DI91  (RAM6_data_in[91 ] ),
    .DI92  (RAM6_data_in[92 ] ),    .DI93  (RAM6_data_in[93 ] ),    .DI94  (RAM6_data_in[94 ] ),    .DI95  (RAM6_data_in[95 ] ),
    .DI96  (RAM6_data_in[96 ] ),    .DI97  (RAM6_data_in[97 ] ),    .DI98  (RAM6_data_in[98 ] ),    .DI99  (RAM6_data_in[99 ] ),
    .DI100 (RAM6_data_in[100] ),    .DI101 (RAM6_data_in[101] ),    .DI102 (RAM6_data_in[102] ),    .DI103 (RAM6_data_in[103] ),
    .DI104 (RAM6_data_in[104] ),    .DI105 (RAM6_data_in[105] ),    .DI106 (RAM6_data_in[106] ),    .DI107 (RAM6_data_in[107] ),
    .DI108 (RAM6_data_in[108] ),    .DI109 (RAM6_data_in[109] ),    .DI110 (RAM6_data_in[110] ),    .DI111 (RAM6_data_in[111] ),
    .DI112 (RAM6_data_in[112] ),    .DI113 (RAM6_data_in[113] ),    .DI114 (RAM6_data_in[114] ),    .DI115 (RAM6_data_in[115] ),
    .DI116 (RAM6_data_in[116] ),    .DI117 (RAM6_data_in[117] ),    .DI118 (RAM6_data_in[118] ),    .DI119 (RAM6_data_in[119] ),
    .DI120 (RAM6_data_in[120] ),    .DI121 (RAM6_data_in[121] ),    .DI122 (RAM6_data_in[122] ),    .DI123 (RAM6_data_in[123] ),
    .DI124 (RAM6_data_in[124] ),    .DI125 (RAM6_data_in[125] ),    .DI126 (RAM6_data_in[126] ),    .DI127 (RAM6_data_in[127] ),

    .A0   (RAM_addr[0]   ),.A1   (RAM_addr[1]   ),.A2   (RAM_addr[2]   ),.A3   (RAM_addr[3]   ),.A4   (RAM_addr[4]   ),.A5   (RAM_addr[5]   ),.A6   (RAM_addr[6]   ),
    .DVSE (1'b0  ),.DVS0 (1'b0  ),.DVS1 (1'b0  ),.DVS2 (1'b0  ),.DVS3 (1'b0  ),
    .WEB0 (~w_WEB6_8[0] ),.WEB1 (~w_WEB6_8[1] ),.WEB2 (~w_WEB6_8[2] ),.WEB3 (~w_WEB6_8[3] ),
    .WEB4 (~w_WEB6_8[4] ),.WEB5 (~w_WEB6_8[5] ),.WEB6 (~w_WEB6_8[6] ),.WEB7 (~w_WEB6_8[7] ),

    .CK    (clka   ),
    .CSB   (1'b0   )
);


SYKB110_128X16X8CM2 u_L2data7_SYKB110_128X16X8CM2(
    .DO0   (RAM7_data_out[128] ),    .DO1   (RAM7_data_out[129] ),    .DO2   (RAM7_data_out[130] ),    .DO3   (RAM7_data_out[131] ),
    .DO4   (RAM7_data_out[132] ),    .DO5   (RAM7_data_out[133] ),    .DO6   (RAM7_data_out[134] ),    .DO7   (RAM7_data_out[135] ),
    .DO8   (RAM7_data_out[136] ),    .DO9   (RAM7_data_out[137] ),    .DO10  (RAM7_data_out[138] ),    .DO11  (RAM7_data_out[139] ),
    .DO12  (RAM7_data_out[140] ),    .DO13  (RAM7_data_out[141] ),    .DO14  (RAM7_data_out[142] ),    .DO15  (RAM7_data_out[143] ),
    .DO16  (RAM7_data_out[144] ),    .DO17  (RAM7_data_out[145] ),    .DO18  (RAM7_data_out[146] ),    .DO19  (RAM7_data_out[147] ),
    .DO20  (RAM7_data_out[148] ),    .DO21  (RAM7_data_out[149] ),    .DO22  (RAM7_data_out[150] ),    .DO23  (RAM7_data_out[151] ),
    .DO24  (RAM7_data_out[152] ),    .DO25  (RAM7_data_out[153] ),    .DO26  (RAM7_data_out[154] ),    .DO27  (RAM7_data_out[155] ),
    .DO28  (RAM7_data_out[156] ),    .DO29  (RAM7_data_out[157] ),    .DO30  (RAM7_data_out[158] ),    .DO31  (RAM7_data_out[159] ),
    .DO32  (RAM7_data_out[160] ),    .DO33  (RAM7_data_out[161] ),    .DO34  (RAM7_data_out[162] ),    .DO35  (RAM7_data_out[163] ),
    .DO36  (RAM7_data_out[164] ),    .DO37  (RAM7_data_out[165] ),    .DO38  (RAM7_data_out[166] ),    .DO39  (RAM7_data_out[167] ),
    .DO40  (RAM7_data_out[168] ),    .DO41  (RAM7_data_out[169] ),    .DO42  (RAM7_data_out[170] ),    .DO43  (RAM7_data_out[171] ),
    .DO44  (RAM7_data_out[172] ),    .DO45  (RAM7_data_out[173] ),    .DO46  (RAM7_data_out[174] ),    .DO47  (RAM7_data_out[175] ),
    .DO48  (RAM7_data_out[176] ),    .DO49  (RAM7_data_out[177] ),    .DO50  (RAM7_data_out[178] ),    .DO51  (RAM7_data_out[179] ),
    .DO52  (RAM7_data_out[180] ),    .DO53  (RAM7_data_out[181] ),    .DO54  (RAM7_data_out[182] ),    .DO55  (RAM7_data_out[183] ),
    .DO56  (RAM7_data_out[184] ),    .DO57  (RAM7_data_out[185] ),    .DO58  (RAM7_data_out[186] ),    .DO59  (RAM7_data_out[187] ),
    .DO60  (RAM7_data_out[188] ),    .DO61  (RAM7_data_out[189] ),    .DO62  (RAM7_data_out[190] ),    .DO63  (RAM7_data_out[191] ),
    .DO64  (RAM7_data_out[192] ),    .DO65  (RAM7_data_out[193] ),    .DO66  (RAM7_data_out[194] ),    .DO67  (RAM7_data_out[195] ),
    .DO68  (RAM7_data_out[196] ),    .DO69  (RAM7_data_out[197] ),    .DO70  (RAM7_data_out[198] ),    .DO71  (RAM7_data_out[199] ),
    .DO72  (RAM7_data_out[200] ),    .DO73  (RAM7_data_out[201] ),    .DO74  (RAM7_data_out[202] ),    .DO75  (RAM7_data_out[203] ),
    .DO76  (RAM7_data_out[204] ),    .DO77  (RAM7_data_out[205] ),    .DO78  (RAM7_data_out[206] ),    .DO79  (RAM7_data_out[207] ),
    .DO80  (RAM7_data_out[208] ),    .DO81  (RAM7_data_out[209] ),    .DO82  (RAM7_data_out[210] ),    .DO83  (RAM7_data_out[211] ),
    .DO84  (RAM7_data_out[212] ),    .DO85  (RAM7_data_out[213] ),    .DO86  (RAM7_data_out[214] ),    .DO87  (RAM7_data_out[215] ),
    .DO88  (RAM7_data_out[216] ),    .DO89  (RAM7_data_out[217] ),    .DO90  (RAM7_data_out[218] ),    .DO91  (RAM7_data_out[219] ),
    .DO92  (RAM7_data_out[220] ),    .DO93  (RAM7_data_out[221] ),    .DO94  (RAM7_data_out[222] ),    .DO95  (RAM7_data_out[223] ),
    .DO96  (RAM7_data_out[224] ),    .DO97  (RAM7_data_out[225] ),    .DO98  (RAM7_data_out[226] ),    .DO99  (RAM7_data_out[227] ),
    .DO100 (RAM7_data_out[228] ),    .DO101 (RAM7_data_out[229] ),    .DO102 (RAM7_data_out[230] ),    .DO103 (RAM7_data_out[231] ),
    .DO104 (RAM7_data_out[232] ),    .DO105 (RAM7_data_out[233] ),    .DO106 (RAM7_data_out[234] ),    .DO107 (RAM7_data_out[235] ),
    .DO108 (RAM7_data_out[236] ),    .DO109 (RAM7_data_out[237] ),    .DO110 (RAM7_data_out[238] ),    .DO111 (RAM7_data_out[239] ),
    .DO112 (RAM7_data_out[240] ),    .DO113 (RAM7_data_out[241] ),    .DO114 (RAM7_data_out[242] ),    .DO115 (RAM7_data_out[243] ),
    .DO116 (RAM7_data_out[244] ),    .DO117 (RAM7_data_out[245] ),    .DO118 (RAM7_data_out[246] ),    .DO119 (RAM7_data_out[247] ),
    .DO120 (RAM7_data_out[248] ),    .DO121 (RAM7_data_out[249] ),    .DO122 (RAM7_data_out[250] ),    .DO123 (RAM7_data_out[251] ),
    .DO124 (RAM7_data_out[252] ),    .DO125 (RAM7_data_out[253] ),    .DO126 (RAM7_data_out[254] ),    .DO127 (RAM7_data_out[255] ),

    .DI0   (RAM7_data_in[128] ),    .DI1   (RAM7_data_in[129] ),    .DI2   (RAM7_data_in[130] ),    .DI3   (RAM7_data_in[131] ),
    .DI4   (RAM7_data_in[132] ),    .DI5   (RAM7_data_in[133] ),    .DI6   (RAM7_data_in[134] ),    .DI7   (RAM7_data_in[135] ),
    .DI8   (RAM7_data_in[136] ),    .DI9   (RAM7_data_in[137] ),    .DI10  (RAM7_data_in[138] ),    .DI11  (RAM7_data_in[139] ),
    .DI12  (RAM7_data_in[140] ),    .DI13  (RAM7_data_in[141] ),    .DI14  (RAM7_data_in[142] ),    .DI15  (RAM7_data_in[143] ),
    .DI16  (RAM7_data_in[144] ),    .DI17  (RAM7_data_in[145] ),    .DI18  (RAM7_data_in[146] ),    .DI19  (RAM7_data_in[147] ),
    .DI20  (RAM7_data_in[148] ),    .DI21  (RAM7_data_in[149] ),    .DI22  (RAM7_data_in[150] ),    .DI23  (RAM7_data_in[151] ),
    .DI24  (RAM7_data_in[152] ),    .DI25  (RAM7_data_in[153] ),    .DI26  (RAM7_data_in[154] ),    .DI27  (RAM7_data_in[155] ),
    .DI28  (RAM7_data_in[156] ),    .DI29  (RAM7_data_in[157] ),    .DI30  (RAM7_data_in[158] ),    .DI31  (RAM7_data_in[159] ),
    .DI32  (RAM7_data_in[160] ),    .DI33  (RAM7_data_in[161] ),    .DI34  (RAM7_data_in[162] ),    .DI35  (RAM7_data_in[163] ),
    .DI36  (RAM7_data_in[164] ),    .DI37  (RAM7_data_in[165] ),    .DI38  (RAM7_data_in[166] ),    .DI39  (RAM7_data_in[167] ),
    .DI40  (RAM7_data_in[168] ),    .DI41  (RAM7_data_in[169] ),    .DI42  (RAM7_data_in[170] ),    .DI43  (RAM7_data_in[171] ),
    .DI44  (RAM7_data_in[172] ),    .DI45  (RAM7_data_in[173] ),    .DI46  (RAM7_data_in[174] ),    .DI47  (RAM7_data_in[175] ),
    .DI48  (RAM7_data_in[176] ),    .DI49  (RAM7_data_in[177] ),    .DI50  (RAM7_data_in[178] ),    .DI51  (RAM7_data_in[179] ),
    .DI52  (RAM7_data_in[180] ),    .DI53  (RAM7_data_in[181] ),    .DI54  (RAM7_data_in[182] ),    .DI55  (RAM7_data_in[183] ),
    .DI56  (RAM7_data_in[184] ),    .DI57  (RAM7_data_in[185] ),    .DI58  (RAM7_data_in[186] ),    .DI59  (RAM7_data_in[187] ),
    .DI60  (RAM7_data_in[188] ),    .DI61  (RAM7_data_in[189] ),    .DI62  (RAM7_data_in[190] ),    .DI63  (RAM7_data_in[191] ),
    .DI64  (RAM7_data_in[192] ),    .DI65  (RAM7_data_in[193] ),    .DI66  (RAM7_data_in[194] ),    .DI67  (RAM7_data_in[195] ),
    .DI68  (RAM7_data_in[196] ),    .DI69  (RAM7_data_in[197] ),    .DI70  (RAM7_data_in[198] ),    .DI71  (RAM7_data_in[199] ),
    .DI72  (RAM7_data_in[200] ),    .DI73  (RAM7_data_in[201] ),    .DI74  (RAM7_data_in[202] ),    .DI75  (RAM7_data_in[203] ),
    .DI76  (RAM7_data_in[204] ),    .DI77  (RAM7_data_in[205] ),    .DI78  (RAM7_data_in[206] ),    .DI79  (RAM7_data_in[207] ),
    .DI80  (RAM7_data_in[208] ),    .DI81  (RAM7_data_in[209] ),    .DI82  (RAM7_data_in[210] ),    .DI83  (RAM7_data_in[211] ),
    .DI84  (RAM7_data_in[212] ),    .DI85  (RAM7_data_in[213] ),    .DI86  (RAM7_data_in[214] ),    .DI87  (RAM7_data_in[215] ),
    .DI88  (RAM7_data_in[216] ),    .DI89  (RAM7_data_in[217] ),    .DI90  (RAM7_data_in[218] ),    .DI91  (RAM7_data_in[219] ),
    .DI92  (RAM7_data_in[220] ),    .DI93  (RAM7_data_in[221] ),    .DI94  (RAM7_data_in[222] ),    .DI95  (RAM7_data_in[223] ),
    .DI96  (RAM7_data_in[224] ),    .DI97  (RAM7_data_in[225] ),    .DI98  (RAM7_data_in[226] ),    .DI99  (RAM7_data_in[227] ),
    .DI100 (RAM7_data_in[228] ),    .DI101 (RAM7_data_in[229] ),    .DI102 (RAM7_data_in[230] ),    .DI103 (RAM7_data_in[231] ),
    .DI104 (RAM7_data_in[232] ),    .DI105 (RAM7_data_in[233] ),    .DI106 (RAM7_data_in[234] ),    .DI107 (RAM7_data_in[235] ),
    .DI108 (RAM7_data_in[236] ),    .DI109 (RAM7_data_in[237] ),    .DI110 (RAM7_data_in[238] ),    .DI111 (RAM7_data_in[239] ),
    .DI112 (RAM7_data_in[240] ),    .DI113 (RAM7_data_in[241] ),    .DI114 (RAM7_data_in[242] ),    .DI115 (RAM7_data_in[243] ),
    .DI116 (RAM7_data_in[244] ),    .DI117 (RAM7_data_in[245] ),    .DI118 (RAM7_data_in[246] ),    .DI119 (RAM7_data_in[247] ),
    .DI120 (RAM7_data_in[248] ),    .DI121 (RAM7_data_in[249] ),    .DI122 (RAM7_data_in[250] ),    .DI123 (RAM7_data_in[251] ),
    .DI124 (RAM7_data_in[252] ),    .DI125 (RAM7_data_in[253] ),    .DI126 (RAM7_data_in[254] ),    .DI127 (RAM7_data_in[255] ),

    .A0   (RAM_addr[0]   ),.A1   (RAM_addr[1]   ),.A2   (RAM_addr[2]   ),.A3   (RAM_addr[3]   ),.A4   (RAM_addr[4]   ),.A5   (RAM_addr[5]   ),.A6   (RAM_addr[6]   ),
    .DVSE (1'b0  ),.DVS0 (1'b0  ),.DVS1 (1'b0  ),.DVS2 (1'b0  ),.DVS3 (1'b0  ),
    .WEB0 (~w_WEB7_8[0] ),.WEB1 (~w_WEB7_8[1] ),.WEB2 (~w_WEB7_8[2] ),.WEB3 (~w_WEB7_8[3] ),
    .WEB4 (~w_WEB7_8[4] ),.WEB5 (~w_WEB7_8[5] ),.WEB6 (~w_WEB7_8[6] ),.WEB7 (~w_WEB7_8[7] ),

    .CK    (clka   ),
    .CSB   (1'b0   )
);


SYKB110_128X16X8CM2 u_L2data8_SYKB110_128X16X8CM2(
    .DO0   (RAM8_data_out[0  ] ),    .DO1   (RAM8_data_out[1  ] ),    .DO2   (RAM8_data_out[2  ] ),    .DO3   (RAM8_data_out[3  ] ),
    .DO4   (RAM8_data_out[4  ] ),    .DO5   (RAM8_data_out[5  ] ),    .DO6   (RAM8_data_out[6  ] ),    .DO7   (RAM8_data_out[7  ] ),
    .DO8   (RAM8_data_out[8  ] ),    .DO9   (RAM8_data_out[9  ] ),    .DO10  (RAM8_data_out[10 ] ),    .DO11  (RAM8_data_out[11 ] ),
    .DO12  (RAM8_data_out[12 ] ),    .DO13  (RAM8_data_out[13 ] ),    .DO14  (RAM8_data_out[14 ] ),    .DO15  (RAM8_data_out[15 ] ),
    .DO16  (RAM8_data_out[16 ] ),    .DO17  (RAM8_data_out[17 ] ),    .DO18  (RAM8_data_out[18 ] ),    .DO19  (RAM8_data_out[19 ] ),
    .DO20  (RAM8_data_out[20 ] ),    .DO21  (RAM8_data_out[21 ] ),    .DO22  (RAM8_data_out[22 ] ),    .DO23  (RAM8_data_out[23 ] ),
    .DO24  (RAM8_data_out[24 ] ),    .DO25  (RAM8_data_out[25 ] ),    .DO26  (RAM8_data_out[26 ] ),    .DO27  (RAM8_data_out[27 ] ),
    .DO28  (RAM8_data_out[28 ] ),    .DO29  (RAM8_data_out[29 ] ),    .DO30  (RAM8_data_out[30 ] ),    .DO31  (RAM8_data_out[31 ] ),
    .DO32  (RAM8_data_out[32 ] ),    .DO33  (RAM8_data_out[33 ] ),    .DO34  (RAM8_data_out[34 ] ),    .DO35  (RAM8_data_out[35 ] ),
    .DO36  (RAM8_data_out[36 ] ),    .DO37  (RAM8_data_out[37 ] ),    .DO38  (RAM8_data_out[38 ] ),    .DO39  (RAM8_data_out[39 ] ),
    .DO40  (RAM8_data_out[40 ] ),    .DO41  (RAM8_data_out[41 ] ),    .DO42  (RAM8_data_out[42 ] ),    .DO43  (RAM8_data_out[43 ] ),
    .DO44  (RAM8_data_out[44 ] ),    .DO45  (RAM8_data_out[45 ] ),    .DO46  (RAM8_data_out[46 ] ),    .DO47  (RAM8_data_out[47 ] ),
    .DO48  (RAM8_data_out[48 ] ),    .DO49  (RAM8_data_out[49 ] ),    .DO50  (RAM8_data_out[50 ] ),    .DO51  (RAM8_data_out[51 ] ),
    .DO52  (RAM8_data_out[52 ] ),    .DO53  (RAM8_data_out[53 ] ),    .DO54  (RAM8_data_out[54 ] ),    .DO55  (RAM8_data_out[55 ] ),
    .DO56  (RAM8_data_out[56 ] ),    .DO57  (RAM8_data_out[57 ] ),    .DO58  (RAM8_data_out[58 ] ),    .DO59  (RAM8_data_out[59 ] ),
    .DO60  (RAM8_data_out[60 ] ),    .DO61  (RAM8_data_out[61 ] ),    .DO62  (RAM8_data_out[62 ] ),    .DO63  (RAM8_data_out[63 ] ),
    .DO64  (RAM8_data_out[64 ] ),    .DO65  (RAM8_data_out[65 ] ),    .DO66  (RAM8_data_out[66 ] ),    .DO67  (RAM8_data_out[67 ] ),
    .DO68  (RAM8_data_out[68 ] ),    .DO69  (RAM8_data_out[69 ] ),    .DO70  (RAM8_data_out[70 ] ),    .DO71  (RAM8_data_out[71 ] ),
    .DO72  (RAM8_data_out[72 ] ),    .DO73  (RAM8_data_out[73 ] ),    .DO74  (RAM8_data_out[74 ] ),    .DO75  (RAM8_data_out[75 ] ),
    .DO76  (RAM8_data_out[76 ] ),    .DO77  (RAM8_data_out[77 ] ),    .DO78  (RAM8_data_out[78 ] ),    .DO79  (RAM8_data_out[79 ] ),
    .DO80  (RAM8_data_out[80 ] ),    .DO81  (RAM8_data_out[81 ] ),    .DO82  (RAM8_data_out[82 ] ),    .DO83  (RAM8_data_out[83 ] ),
    .DO84  (RAM8_data_out[84 ] ),    .DO85  (RAM8_data_out[85 ] ),    .DO86  (RAM8_data_out[86 ] ),    .DO87  (RAM8_data_out[87 ] ),
    .DO88  (RAM8_data_out[88 ] ),    .DO89  (RAM8_data_out[89 ] ),    .DO90  (RAM8_data_out[90 ] ),    .DO91  (RAM8_data_out[91 ] ),
    .DO92  (RAM8_data_out[92 ] ),    .DO93  (RAM8_data_out[93 ] ),    .DO94  (RAM8_data_out[94 ] ),    .DO95  (RAM8_data_out[95 ] ),
    .DO96  (RAM8_data_out[96 ] ),    .DO97  (RAM8_data_out[97 ] ),    .DO98  (RAM8_data_out[98 ] ),    .DO99  (RAM8_data_out[99 ] ),
    .DO100 (RAM8_data_out[100] ),    .DO101 (RAM8_data_out[101] ),    .DO102 (RAM8_data_out[102] ),    .DO103 (RAM8_data_out[103] ),
    .DO104 (RAM8_data_out[104] ),    .DO105 (RAM8_data_out[105] ),    .DO106 (RAM8_data_out[106] ),    .DO107 (RAM8_data_out[107] ),
    .DO108 (RAM8_data_out[108] ),    .DO109 (RAM8_data_out[109] ),    .DO110 (RAM8_data_out[110] ),    .DO111 (RAM8_data_out[111] ),
    .DO112 (RAM8_data_out[112] ),    .DO113 (RAM8_data_out[113] ),    .DO114 (RAM8_data_out[114] ),    .DO115 (RAM8_data_out[115] ),
    .DO116 (RAM8_data_out[116] ),    .DO117 (RAM8_data_out[117] ),    .DO118 (RAM8_data_out[118] ),    .DO119 (RAM8_data_out[119] ),
    .DO120 (RAM8_data_out[120] ),    .DO121 (RAM8_data_out[121] ),    .DO122 (RAM8_data_out[122] ),    .DO123 (RAM8_data_out[123] ),
    .DO124 (RAM8_data_out[124] ),    .DO125 (RAM8_data_out[125] ),    .DO126 (RAM8_data_out[126] ),    .DO127 (RAM8_data_out[127] ),

    .DI0   (RAM8_data_in[0  ] ),    .DI1   (RAM8_data_in[1  ] ),    .DI2   (RAM8_data_in[2  ] ),    .DI3   (RAM8_data_in[3  ] ),
    .DI4   (RAM8_data_in[4  ] ),    .DI5   (RAM8_data_in[5  ] ),    .DI6   (RAM8_data_in[6  ] ),    .DI7   (RAM8_data_in[7  ] ),
    .DI8   (RAM8_data_in[8  ] ),    .DI9   (RAM8_data_in[9  ] ),    .DI10  (RAM8_data_in[10 ] ),    .DI11  (RAM8_data_in[11 ] ),
    .DI12  (RAM8_data_in[12 ] ),    .DI13  (RAM8_data_in[13 ] ),    .DI14  (RAM8_data_in[14 ] ),    .DI15  (RAM8_data_in[15 ] ),
    .DI16  (RAM8_data_in[16 ] ),    .DI17  (RAM8_data_in[17 ] ),    .DI18  (RAM8_data_in[18 ] ),    .DI19  (RAM8_data_in[19 ] ),
    .DI20  (RAM8_data_in[20 ] ),    .DI21  (RAM8_data_in[21 ] ),    .DI22  (RAM8_data_in[22 ] ),    .DI23  (RAM8_data_in[23 ] ),
    .DI24  (RAM8_data_in[24 ] ),    .DI25  (RAM8_data_in[25 ] ),    .DI26  (RAM8_data_in[26 ] ),    .DI27  (RAM8_data_in[27 ] ),
    .DI28  (RAM8_data_in[28 ] ),    .DI29  (RAM8_data_in[29 ] ),    .DI30  (RAM8_data_in[30 ] ),    .DI31  (RAM8_data_in[31 ] ),
    .DI32  (RAM8_data_in[32 ] ),    .DI33  (RAM8_data_in[33 ] ),    .DI34  (RAM8_data_in[34 ] ),    .DI35  (RAM8_data_in[35 ] ),
    .DI36  (RAM8_data_in[36 ] ),    .DI37  (RAM8_data_in[37 ] ),    .DI38  (RAM8_data_in[38 ] ),    .DI39  (RAM8_data_in[39 ] ),
    .DI40  (RAM8_data_in[40 ] ),    .DI41  (RAM8_data_in[41 ] ),    .DI42  (RAM8_data_in[42 ] ),    .DI43  (RAM8_data_in[43 ] ),
    .DI44  (RAM8_data_in[44 ] ),    .DI45  (RAM8_data_in[45 ] ),    .DI46  (RAM8_data_in[46 ] ),    .DI47  (RAM8_data_in[47 ] ),
    .DI48  (RAM8_data_in[48 ] ),    .DI49  (RAM8_data_in[49 ] ),    .DI50  (RAM8_data_in[50 ] ),    .DI51  (RAM8_data_in[51 ] ),
    .DI52  (RAM8_data_in[52 ] ),    .DI53  (RAM8_data_in[53 ] ),    .DI54  (RAM8_data_in[54 ] ),    .DI55  (RAM8_data_in[55 ] ),
    .DI56  (RAM8_data_in[56 ] ),    .DI57  (RAM8_data_in[57 ] ),    .DI58  (RAM8_data_in[58 ] ),    .DI59  (RAM8_data_in[59 ] ),
    .DI60  (RAM8_data_in[60 ] ),    .DI61  (RAM8_data_in[61 ] ),    .DI62  (RAM8_data_in[62 ] ),    .DI63  (RAM8_data_in[63 ] ),
    .DI64  (RAM8_data_in[64 ] ),    .DI65  (RAM8_data_in[65 ] ),    .DI66  (RAM8_data_in[66 ] ),    .DI67  (RAM8_data_in[67 ] ),
    .DI68  (RAM8_data_in[68 ] ),    .DI69  (RAM8_data_in[69 ] ),    .DI70  (RAM8_data_in[70 ] ),    .DI71  (RAM8_data_in[71 ] ),
    .DI72  (RAM8_data_in[72 ] ),    .DI73  (RAM8_data_in[73 ] ),    .DI74  (RAM8_data_in[74 ] ),    .DI75  (RAM8_data_in[75 ] ),
    .DI76  (RAM8_data_in[76 ] ),    .DI77  (RAM8_data_in[77 ] ),    .DI78  (RAM8_data_in[78 ] ),    .DI79  (RAM8_data_in[79 ] ),
    .DI80  (RAM8_data_in[80 ] ),    .DI81  (RAM8_data_in[81 ] ),    .DI82  (RAM8_data_in[82 ] ),    .DI83  (RAM8_data_in[83 ] ),
    .DI84  (RAM8_data_in[84 ] ),    .DI85  (RAM8_data_in[85 ] ),    .DI86  (RAM8_data_in[86 ] ),    .DI87  (RAM8_data_in[87 ] ),
    .DI88  (RAM8_data_in[88 ] ),    .DI89  (RAM8_data_in[89 ] ),    .DI90  (RAM8_data_in[90 ] ),    .DI91  (RAM8_data_in[91 ] ),
    .DI92  (RAM8_data_in[92 ] ),    .DI93  (RAM8_data_in[93 ] ),    .DI94  (RAM8_data_in[94 ] ),    .DI95  (RAM8_data_in[95 ] ),
    .DI96  (RAM8_data_in[96 ] ),    .DI97  (RAM8_data_in[97 ] ),    .DI98  (RAM8_data_in[98 ] ),    .DI99  (RAM8_data_in[99 ] ),
    .DI100 (RAM8_data_in[100] ),    .DI101 (RAM8_data_in[101] ),    .DI102 (RAM8_data_in[102] ),    .DI103 (RAM8_data_in[103] ),
    .DI104 (RAM8_data_in[104] ),    .DI105 (RAM8_data_in[105] ),    .DI106 (RAM8_data_in[106] ),    .DI107 (RAM8_data_in[107] ),
    .DI108 (RAM8_data_in[108] ),    .DI109 (RAM8_data_in[109] ),    .DI110 (RAM8_data_in[110] ),    .DI111 (RAM8_data_in[111] ),
    .DI112 (RAM8_data_in[112] ),    .DI113 (RAM8_data_in[113] ),    .DI114 (RAM8_data_in[114] ),    .DI115 (RAM8_data_in[115] ),
    .DI116 (RAM8_data_in[116] ),    .DI117 (RAM8_data_in[117] ),    .DI118 (RAM8_data_in[118] ),    .DI119 (RAM8_data_in[119] ),
    .DI120 (RAM8_data_in[120] ),    .DI121 (RAM8_data_in[121] ),    .DI122 (RAM8_data_in[122] ),    .DI123 (RAM8_data_in[123] ),
    .DI124 (RAM8_data_in[124] ),    .DI125 (RAM8_data_in[125] ),    .DI126 (RAM8_data_in[126] ),    .DI127 (RAM8_data_in[127] ),

    .A0   (RAM_addr[0]   ),.A1   (RAM_addr[1]   ),.A2   (RAM_addr[2]   ),.A3   (RAM_addr[3]   ),.A4   (RAM_addr[4]   ),.A5   (RAM_addr[5]   ),.A6   (RAM_addr[6]   ),
    .DVSE (1'b0  ),.DVS0 (1'b0  ),.DVS1 (1'b0  ),.DVS2 (1'b0  ),.DVS3 (1'b0  ),
    .WEB0 (~w_WEB8_8[0] ),.WEB1 (~w_WEB8_8[1] ),.WEB2 (~w_WEB8_8[2] ),.WEB3 (~w_WEB8_8[3] ),
    .WEB4 (~w_WEB8_8[4] ),.WEB5 (~w_WEB8_8[5] ),.WEB6 (~w_WEB8_8[6] ),.WEB7 (~w_WEB8_8[7] ),

    .CK    (clka   ),
    .CSB   (1'b0   )
);


SYKB110_128X16X8CM2 u_L2data9_SYKB110_128X16X8CM2(
    .DO0   (RAM9_data_out[128] ),    .DO1   (RAM9_data_out[129] ),    .DO2   (RAM9_data_out[130] ),    .DO3   (RAM9_data_out[131] ),
    .DO4   (RAM9_data_out[132] ),    .DO5   (RAM9_data_out[133] ),    .DO6   (RAM9_data_out[134] ),    .DO7   (RAM9_data_out[135] ),
    .DO8   (RAM9_data_out[136] ),    .DO9   (RAM9_data_out[137] ),    .DO10  (RAM9_data_out[138] ),    .DO11  (RAM9_data_out[139] ),
    .DO12  (RAM9_data_out[140] ),    .DO13  (RAM9_data_out[141] ),    .DO14  (RAM9_data_out[142] ),    .DO15  (RAM9_data_out[143] ),
    .DO16  (RAM9_data_out[144] ),    .DO17  (RAM9_data_out[145] ),    .DO18  (RAM9_data_out[146] ),    .DO19  (RAM9_data_out[147] ),
    .DO20  (RAM9_data_out[148] ),    .DO21  (RAM9_data_out[149] ),    .DO22  (RAM9_data_out[150] ),    .DO23  (RAM9_data_out[151] ),
    .DO24  (RAM9_data_out[152] ),    .DO25  (RAM9_data_out[153] ),    .DO26  (RAM9_data_out[154] ),    .DO27  (RAM9_data_out[155] ),
    .DO28  (RAM9_data_out[156] ),    .DO29  (RAM9_data_out[157] ),    .DO30  (RAM9_data_out[158] ),    .DO31  (RAM9_data_out[159] ),
    .DO32  (RAM9_data_out[160] ),    .DO33  (RAM9_data_out[161] ),    .DO34  (RAM9_data_out[162] ),    .DO35  (RAM9_data_out[163] ),
    .DO36  (RAM9_data_out[164] ),    .DO37  (RAM9_data_out[165] ),    .DO38  (RAM9_data_out[166] ),    .DO39  (RAM9_data_out[167] ),
    .DO40  (RAM9_data_out[168] ),    .DO41  (RAM9_data_out[169] ),    .DO42  (RAM9_data_out[170] ),    .DO43  (RAM9_data_out[171] ),
    .DO44  (RAM9_data_out[172] ),    .DO45  (RAM9_data_out[173] ),    .DO46  (RAM9_data_out[174] ),    .DO47  (RAM9_data_out[175] ),
    .DO48  (RAM9_data_out[176] ),    .DO49  (RAM9_data_out[177] ),    .DO50  (RAM9_data_out[178] ),    .DO51  (RAM9_data_out[179] ),
    .DO52  (RAM9_data_out[180] ),    .DO53  (RAM9_data_out[181] ),    .DO54  (RAM9_data_out[182] ),    .DO55  (RAM9_data_out[183] ),
    .DO56  (RAM9_data_out[184] ),    .DO57  (RAM9_data_out[185] ),    .DO58  (RAM9_data_out[186] ),    .DO59  (RAM9_data_out[187] ),
    .DO60  (RAM9_data_out[188] ),    .DO61  (RAM9_data_out[189] ),    .DO62  (RAM9_data_out[190] ),    .DO63  (RAM9_data_out[191] ),
    .DO64  (RAM9_data_out[192] ),    .DO65  (RAM9_data_out[193] ),    .DO66  (RAM9_data_out[194] ),    .DO67  (RAM9_data_out[195] ),
    .DO68  (RAM9_data_out[196] ),    .DO69  (RAM9_data_out[197] ),    .DO70  (RAM9_data_out[198] ),    .DO71  (RAM9_data_out[199] ),
    .DO72  (RAM9_data_out[200] ),    .DO73  (RAM9_data_out[201] ),    .DO74  (RAM9_data_out[202] ),    .DO75  (RAM9_data_out[203] ),
    .DO76  (RAM9_data_out[204] ),    .DO77  (RAM9_data_out[205] ),    .DO78  (RAM9_data_out[206] ),    .DO79  (RAM9_data_out[207] ),
    .DO80  (RAM9_data_out[208] ),    .DO81  (RAM9_data_out[209] ),    .DO82  (RAM9_data_out[210] ),    .DO83  (RAM9_data_out[211] ),
    .DO84  (RAM9_data_out[212] ),    .DO85  (RAM9_data_out[213] ),    .DO86  (RAM9_data_out[214] ),    .DO87  (RAM9_data_out[215] ),
    .DO88  (RAM9_data_out[216] ),    .DO89  (RAM9_data_out[217] ),    .DO90  (RAM9_data_out[218] ),    .DO91  (RAM9_data_out[219] ),
    .DO92  (RAM9_data_out[220] ),    .DO93  (RAM9_data_out[221] ),    .DO94  (RAM9_data_out[222] ),    .DO95  (RAM9_data_out[223] ),
    .DO96  (RAM9_data_out[224] ),    .DO97  (RAM9_data_out[225] ),    .DO98  (RAM9_data_out[226] ),    .DO99  (RAM9_data_out[227] ),
    .DO100 (RAM9_data_out[228] ),    .DO101 (RAM9_data_out[229] ),    .DO102 (RAM9_data_out[230] ),    .DO103 (RAM9_data_out[231] ),
    .DO104 (RAM9_data_out[232] ),    .DO105 (RAM9_data_out[233] ),    .DO106 (RAM9_data_out[234] ),    .DO107 (RAM9_data_out[235] ),
    .DO108 (RAM9_data_out[236] ),    .DO109 (RAM9_data_out[237] ),    .DO110 (RAM9_data_out[238] ),    .DO111 (RAM9_data_out[239] ),
    .DO112 (RAM9_data_out[240] ),    .DO113 (RAM9_data_out[241] ),    .DO114 (RAM9_data_out[242] ),    .DO115 (RAM9_data_out[243] ),
    .DO116 (RAM9_data_out[244] ),    .DO117 (RAM9_data_out[245] ),    .DO118 (RAM9_data_out[246] ),    .DO119 (RAM9_data_out[247] ),
    .DO120 (RAM9_data_out[248] ),    .DO121 (RAM9_data_out[249] ),    .DO122 (RAM9_data_out[250] ),    .DO123 (RAM9_data_out[251] ),
    .DO124 (RAM9_data_out[252] ),    .DO125 (RAM9_data_out[253] ),    .DO126 (RAM9_data_out[254] ),    .DO127 (RAM9_data_out[255] ),

    .DI0   (RAM9_data_in[128] ),    .DI1   (RAM9_data_in[129] ),    .DI2   (RAM9_data_in[130] ),    .DI3   (RAM9_data_in[131] ),
    .DI4   (RAM9_data_in[132] ),    .DI5   (RAM9_data_in[133] ),    .DI6   (RAM9_data_in[134] ),    .DI7   (RAM9_data_in[135] ),
    .DI8   (RAM9_data_in[136] ),    .DI9   (RAM9_data_in[137] ),    .DI10  (RAM9_data_in[138] ),    .DI11  (RAM9_data_in[139] ),
    .DI12  (RAM9_data_in[140] ),    .DI13  (RAM9_data_in[141] ),    .DI14  (RAM9_data_in[142] ),    .DI15  (RAM9_data_in[143] ),
    .DI16  (RAM9_data_in[144] ),    .DI17  (RAM9_data_in[145] ),    .DI18  (RAM9_data_in[146] ),    .DI19  (RAM9_data_in[147] ),
    .DI20  (RAM9_data_in[148] ),    .DI21  (RAM9_data_in[149] ),    .DI22  (RAM9_data_in[150] ),    .DI23  (RAM9_data_in[151] ),
    .DI24  (RAM9_data_in[152] ),    .DI25  (RAM9_data_in[153] ),    .DI26  (RAM9_data_in[154] ),    .DI27  (RAM9_data_in[155] ),
    .DI28  (RAM9_data_in[156] ),    .DI29  (RAM9_data_in[157] ),    .DI30  (RAM9_data_in[158] ),    .DI31  (RAM9_data_in[159] ),
    .DI32  (RAM9_data_in[160] ),    .DI33  (RAM9_data_in[161] ),    .DI34  (RAM9_data_in[162] ),    .DI35  (RAM9_data_in[163] ),
    .DI36  (RAM9_data_in[164] ),    .DI37  (RAM9_data_in[165] ),    .DI38  (RAM9_data_in[166] ),    .DI39  (RAM9_data_in[167] ),
    .DI40  (RAM9_data_in[168] ),    .DI41  (RAM9_data_in[169] ),    .DI42  (RAM9_data_in[170] ),    .DI43  (RAM9_data_in[171] ),
    .DI44  (RAM9_data_in[172] ),    .DI45  (RAM9_data_in[173] ),    .DI46  (RAM9_data_in[174] ),    .DI47  (RAM9_data_in[175] ),
    .DI48  (RAM9_data_in[176] ),    .DI49  (RAM9_data_in[177] ),    .DI50  (RAM9_data_in[178] ),    .DI51  (RAM9_data_in[179] ),
    .DI52  (RAM9_data_in[180] ),    .DI53  (RAM9_data_in[181] ),    .DI54  (RAM9_data_in[182] ),    .DI55  (RAM9_data_in[183] ),
    .DI56  (RAM9_data_in[184] ),    .DI57  (RAM9_data_in[185] ),    .DI58  (RAM9_data_in[186] ),    .DI59  (RAM9_data_in[187] ),
    .DI60  (RAM9_data_in[188] ),    .DI61  (RAM9_data_in[189] ),    .DI62  (RAM9_data_in[190] ),    .DI63  (RAM9_data_in[191] ),
    .DI64  (RAM9_data_in[192] ),    .DI65  (RAM9_data_in[193] ),    .DI66  (RAM9_data_in[194] ),    .DI67  (RAM9_data_in[195] ),
    .DI68  (RAM9_data_in[196] ),    .DI69  (RAM9_data_in[197] ),    .DI70  (RAM9_data_in[198] ),    .DI71  (RAM9_data_in[199] ),
    .DI72  (RAM9_data_in[200] ),    .DI73  (RAM9_data_in[201] ),    .DI74  (RAM9_data_in[202] ),    .DI75  (RAM9_data_in[203] ),
    .DI76  (RAM9_data_in[204] ),    .DI77  (RAM9_data_in[205] ),    .DI78  (RAM9_data_in[206] ),    .DI79  (RAM9_data_in[207] ),
    .DI80  (RAM9_data_in[208] ),    .DI81  (RAM9_data_in[209] ),    .DI82  (RAM9_data_in[210] ),    .DI83  (RAM9_data_in[211] ),
    .DI84  (RAM9_data_in[212] ),    .DI85  (RAM9_data_in[213] ),    .DI86  (RAM9_data_in[214] ),    .DI87  (RAM9_data_in[215] ),
    .DI88  (RAM9_data_in[216] ),    .DI89  (RAM9_data_in[217] ),    .DI90  (RAM9_data_in[218] ),    .DI91  (RAM9_data_in[219] ),
    .DI92  (RAM9_data_in[220] ),    .DI93  (RAM9_data_in[221] ),    .DI94  (RAM9_data_in[222] ),    .DI95  (RAM9_data_in[223] ),
    .DI96  (RAM9_data_in[224] ),    .DI97  (RAM9_data_in[225] ),    .DI98  (RAM9_data_in[226] ),    .DI99  (RAM9_data_in[227] ),
    .DI100 (RAM9_data_in[228] ),    .DI101 (RAM9_data_in[229] ),    .DI102 (RAM9_data_in[230] ),    .DI103 (RAM9_data_in[231] ),
    .DI104 (RAM9_data_in[232] ),    .DI105 (RAM9_data_in[233] ),    .DI106 (RAM9_data_in[234] ),    .DI107 (RAM9_data_in[235] ),
    .DI108 (RAM9_data_in[236] ),    .DI109 (RAM9_data_in[237] ),    .DI110 (RAM9_data_in[238] ),    .DI111 (RAM9_data_in[239] ),
    .DI112 (RAM9_data_in[240] ),    .DI113 (RAM9_data_in[241] ),    .DI114 (RAM9_data_in[242] ),    .DI115 (RAM9_data_in[243] ),
    .DI116 (RAM9_data_in[244] ),    .DI117 (RAM9_data_in[245] ),    .DI118 (RAM9_data_in[246] ),    .DI119 (RAM9_data_in[247] ),
    .DI120 (RAM9_data_in[248] ),    .DI121 (RAM9_data_in[249] ),    .DI122 (RAM9_data_in[250] ),    .DI123 (RAM9_data_in[251] ),
    .DI124 (RAM9_data_in[252] ),    .DI125 (RAM9_data_in[253] ),    .DI126 (RAM9_data_in[254] ),    .DI127 (RAM9_data_in[255] ),

    .A0   (RAM_addr[0]   ),.A1   (RAM_addr[1]   ),.A2   (RAM_addr[2]   ),.A3   (RAM_addr[3]   ),.A4   (RAM_addr[4]   ),.A5   (RAM_addr[5]   ),.A6   (RAM_addr[6]   ),
    .DVSE (1'b0  ),.DVS0 (1'b0  ),.DVS1 (1'b0  ),.DVS2 (1'b0  ),.DVS3 (1'b0  ),
    .WEB0 (~w_WEB9_8[0] ),.WEB1 (~w_WEB9_8[1] ),.WEB2 (~w_WEB9_8[2] ),.WEB3 (~w_WEB9_8[3] ),
    .WEB4 (~w_WEB9_8[4] ),.WEB5 (~w_WEB9_8[5] ),.WEB6 (~w_WEB9_8[6] ),.WEB7 (~w_WEB9_8[7] ),

    .CK    (clka   ),
    .CSB   (1'b0   )
);


SYKB110_128X16X8CM2 u_L2data10_SYKB110_128X16X8CM2(
    .DO0   (RAM10_data_out[0  ] ),    .DO1   (RAM10_data_out[1  ] ),    .DO2   (RAM10_data_out[2  ] ),    .DO3   (RAM10_data_out[3  ] ),
    .DO4   (RAM10_data_out[4  ] ),    .DO5   (RAM10_data_out[5  ] ),    .DO6   (RAM10_data_out[6  ] ),    .DO7   (RAM10_data_out[7  ] ),
    .DO8   (RAM10_data_out[8  ] ),    .DO9   (RAM10_data_out[9  ] ),    .DO10  (RAM10_data_out[10 ] ),    .DO11  (RAM10_data_out[11 ] ),
    .DO12  (RAM10_data_out[12 ] ),    .DO13  (RAM10_data_out[13 ] ),    .DO14  (RAM10_data_out[14 ] ),    .DO15  (RAM10_data_out[15 ] ),
    .DO16  (RAM10_data_out[16 ] ),    .DO17  (RAM10_data_out[17 ] ),    .DO18  (RAM10_data_out[18 ] ),    .DO19  (RAM10_data_out[19 ] ),
    .DO20  (RAM10_data_out[20 ] ),    .DO21  (RAM10_data_out[21 ] ),    .DO22  (RAM10_data_out[22 ] ),    .DO23  (RAM10_data_out[23 ] ),
    .DO24  (RAM10_data_out[24 ] ),    .DO25  (RAM10_data_out[25 ] ),    .DO26  (RAM10_data_out[26 ] ),    .DO27  (RAM10_data_out[27 ] ),
    .DO28  (RAM10_data_out[28 ] ),    .DO29  (RAM10_data_out[29 ] ),    .DO30  (RAM10_data_out[30 ] ),    .DO31  (RAM10_data_out[31 ] ),
    .DO32  (RAM10_data_out[32 ] ),    .DO33  (RAM10_data_out[33 ] ),    .DO34  (RAM10_data_out[34 ] ),    .DO35  (RAM10_data_out[35 ] ),
    .DO36  (RAM10_data_out[36 ] ),    .DO37  (RAM10_data_out[37 ] ),    .DO38  (RAM10_data_out[38 ] ),    .DO39  (RAM10_data_out[39 ] ),
    .DO40  (RAM10_data_out[40 ] ),    .DO41  (RAM10_data_out[41 ] ),    .DO42  (RAM10_data_out[42 ] ),    .DO43  (RAM10_data_out[43 ] ),
    .DO44  (RAM10_data_out[44 ] ),    .DO45  (RAM10_data_out[45 ] ),    .DO46  (RAM10_data_out[46 ] ),    .DO47  (RAM10_data_out[47 ] ),
    .DO48  (RAM10_data_out[48 ] ),    .DO49  (RAM10_data_out[49 ] ),    .DO50  (RAM10_data_out[50 ] ),    .DO51  (RAM10_data_out[51 ] ),
    .DO52  (RAM10_data_out[52 ] ),    .DO53  (RAM10_data_out[53 ] ),    .DO54  (RAM10_data_out[54 ] ),    .DO55  (RAM10_data_out[55 ] ),
    .DO56  (RAM10_data_out[56 ] ),    .DO57  (RAM10_data_out[57 ] ),    .DO58  (RAM10_data_out[58 ] ),    .DO59  (RAM10_data_out[59 ] ),
    .DO60  (RAM10_data_out[60 ] ),    .DO61  (RAM10_data_out[61 ] ),    .DO62  (RAM10_data_out[62 ] ),    .DO63  (RAM10_data_out[63 ] ),
    .DO64  (RAM10_data_out[64 ] ),    .DO65  (RAM10_data_out[65 ] ),    .DO66  (RAM10_data_out[66 ] ),    .DO67  (RAM10_data_out[67 ] ),
    .DO68  (RAM10_data_out[68 ] ),    .DO69  (RAM10_data_out[69 ] ),    .DO70  (RAM10_data_out[70 ] ),    .DO71  (RAM10_data_out[71 ] ),
    .DO72  (RAM10_data_out[72 ] ),    .DO73  (RAM10_data_out[73 ] ),    .DO74  (RAM10_data_out[74 ] ),    .DO75  (RAM10_data_out[75 ] ),
    .DO76  (RAM10_data_out[76 ] ),    .DO77  (RAM10_data_out[77 ] ),    .DO78  (RAM10_data_out[78 ] ),    .DO79  (RAM10_data_out[79 ] ),
    .DO80  (RAM10_data_out[80 ] ),    .DO81  (RAM10_data_out[81 ] ),    .DO82  (RAM10_data_out[82 ] ),    .DO83  (RAM10_data_out[83 ] ),
    .DO84  (RAM10_data_out[84 ] ),    .DO85  (RAM10_data_out[85 ] ),    .DO86  (RAM10_data_out[86 ] ),    .DO87  (RAM10_data_out[87 ] ),
    .DO88  (RAM10_data_out[88 ] ),    .DO89  (RAM10_data_out[89 ] ),    .DO90  (RAM10_data_out[90 ] ),    .DO91  (RAM10_data_out[91 ] ),
    .DO92  (RAM10_data_out[92 ] ),    .DO93  (RAM10_data_out[93 ] ),    .DO94  (RAM10_data_out[94 ] ),    .DO95  (RAM10_data_out[95 ] ),
    .DO96  (RAM10_data_out[96 ] ),    .DO97  (RAM10_data_out[97 ] ),    .DO98  (RAM10_data_out[98 ] ),    .DO99  (RAM10_data_out[99 ] ),
    .DO100 (RAM10_data_out[100] ),    .DO101 (RAM10_data_out[101] ),    .DO102 (RAM10_data_out[102] ),    .DO103 (RAM10_data_out[103] ),
    .DO104 (RAM10_data_out[104] ),    .DO105 (RAM10_data_out[105] ),    .DO106 (RAM10_data_out[106] ),    .DO107 (RAM10_data_out[107] ),
    .DO108 (RAM10_data_out[108] ),    .DO109 (RAM10_data_out[109] ),    .DO110 (RAM10_data_out[110] ),    .DO111 (RAM10_data_out[111] ),
    .DO112 (RAM10_data_out[112] ),    .DO113 (RAM10_data_out[113] ),    .DO114 (RAM10_data_out[114] ),    .DO115 (RAM10_data_out[115] ),
    .DO116 (RAM10_data_out[116] ),    .DO117 (RAM10_data_out[117] ),    .DO118 (RAM10_data_out[118] ),    .DO119 (RAM10_data_out[119] ),
    .DO120 (RAM10_data_out[120] ),    .DO121 (RAM10_data_out[121] ),    .DO122 (RAM10_data_out[122] ),    .DO123 (RAM10_data_out[123] ),
    .DO124 (RAM10_data_out[124] ),    .DO125 (RAM10_data_out[125] ),    .DO126 (RAM10_data_out[126] ),    .DO127 (RAM10_data_out[127] ),

    .DI0   (RAM10_data_in[0  ] ),    .DI1   (RAM10_data_in[1  ] ),    .DI2   (RAM10_data_in[2  ] ),    .DI3   (RAM10_data_in[3  ] ),
    .DI4   (RAM10_data_in[4  ] ),    .DI5   (RAM10_data_in[5  ] ),    .DI6   (RAM10_data_in[6  ] ),    .DI7   (RAM10_data_in[7  ] ),
    .DI8   (RAM10_data_in[8  ] ),    .DI9   (RAM10_data_in[9  ] ),    .DI10  (RAM10_data_in[10 ] ),    .DI11  (RAM10_data_in[11 ] ),
    .DI12  (RAM10_data_in[12 ] ),    .DI13  (RAM10_data_in[13 ] ),    .DI14  (RAM10_data_in[14 ] ),    .DI15  (RAM10_data_in[15 ] ),
    .DI16  (RAM10_data_in[16 ] ),    .DI17  (RAM10_data_in[17 ] ),    .DI18  (RAM10_data_in[18 ] ),    .DI19  (RAM10_data_in[19 ] ),
    .DI20  (RAM10_data_in[20 ] ),    .DI21  (RAM10_data_in[21 ] ),    .DI22  (RAM10_data_in[22 ] ),    .DI23  (RAM10_data_in[23 ] ),
    .DI24  (RAM10_data_in[24 ] ),    .DI25  (RAM10_data_in[25 ] ),    .DI26  (RAM10_data_in[26 ] ),    .DI27  (RAM10_data_in[27 ] ),
    .DI28  (RAM10_data_in[28 ] ),    .DI29  (RAM10_data_in[29 ] ),    .DI30  (RAM10_data_in[30 ] ),    .DI31  (RAM10_data_in[31 ] ),
    .DI32  (RAM10_data_in[32 ] ),    .DI33  (RAM10_data_in[33 ] ),    .DI34  (RAM10_data_in[34 ] ),    .DI35  (RAM10_data_in[35 ] ),
    .DI36  (RAM10_data_in[36 ] ),    .DI37  (RAM10_data_in[37 ] ),    .DI38  (RAM10_data_in[38 ] ),    .DI39  (RAM10_data_in[39 ] ),
    .DI40  (RAM10_data_in[40 ] ),    .DI41  (RAM10_data_in[41 ] ),    .DI42  (RAM10_data_in[42 ] ),    .DI43  (RAM10_data_in[43 ] ),
    .DI44  (RAM10_data_in[44 ] ),    .DI45  (RAM10_data_in[45 ] ),    .DI46  (RAM10_data_in[46 ] ),    .DI47  (RAM10_data_in[47 ] ),
    .DI48  (RAM10_data_in[48 ] ),    .DI49  (RAM10_data_in[49 ] ),    .DI50  (RAM10_data_in[50 ] ),    .DI51  (RAM10_data_in[51 ] ),
    .DI52  (RAM10_data_in[52 ] ),    .DI53  (RAM10_data_in[53 ] ),    .DI54  (RAM10_data_in[54 ] ),    .DI55  (RAM10_data_in[55 ] ),
    .DI56  (RAM10_data_in[56 ] ),    .DI57  (RAM10_data_in[57 ] ),    .DI58  (RAM10_data_in[58 ] ),    .DI59  (RAM10_data_in[59 ] ),
    .DI60  (RAM10_data_in[60 ] ),    .DI61  (RAM10_data_in[61 ] ),    .DI62  (RAM10_data_in[62 ] ),    .DI63  (RAM10_data_in[63 ] ),
    .DI64  (RAM10_data_in[64 ] ),    .DI65  (RAM10_data_in[65 ] ),    .DI66  (RAM10_data_in[66 ] ),    .DI67  (RAM10_data_in[67 ] ),
    .DI68  (RAM10_data_in[68 ] ),    .DI69  (RAM10_data_in[69 ] ),    .DI70  (RAM10_data_in[70 ] ),    .DI71  (RAM10_data_in[71 ] ),
    .DI72  (RAM10_data_in[72 ] ),    .DI73  (RAM10_data_in[73 ] ),    .DI74  (RAM10_data_in[74 ] ),    .DI75  (RAM10_data_in[75 ] ),
    .DI76  (RAM10_data_in[76 ] ),    .DI77  (RAM10_data_in[77 ] ),    .DI78  (RAM10_data_in[78 ] ),    .DI79  (RAM10_data_in[79 ] ),
    .DI80  (RAM10_data_in[80 ] ),    .DI81  (RAM10_data_in[81 ] ),    .DI82  (RAM10_data_in[82 ] ),    .DI83  (RAM10_data_in[83 ] ),
    .DI84  (RAM10_data_in[84 ] ),    .DI85  (RAM10_data_in[85 ] ),    .DI86  (RAM10_data_in[86 ] ),    .DI87  (RAM10_data_in[87 ] ),
    .DI88  (RAM10_data_in[88 ] ),    .DI89  (RAM10_data_in[89 ] ),    .DI90  (RAM10_data_in[90 ] ),    .DI91  (RAM10_data_in[91 ] ),
    .DI92  (RAM10_data_in[92 ] ),    .DI93  (RAM10_data_in[93 ] ),    .DI94  (RAM10_data_in[94 ] ),    .DI95  (RAM10_data_in[95 ] ),
    .DI96  (RAM10_data_in[96 ] ),    .DI97  (RAM10_data_in[97 ] ),    .DI98  (RAM10_data_in[98 ] ),    .DI99  (RAM10_data_in[99 ] ),
    .DI100 (RAM10_data_in[100] ),    .DI101 (RAM10_data_in[101] ),    .DI102 (RAM10_data_in[102] ),    .DI103 (RAM10_data_in[103] ),
    .DI104 (RAM10_data_in[104] ),    .DI105 (RAM10_data_in[105] ),    .DI106 (RAM10_data_in[106] ),    .DI107 (RAM10_data_in[107] ),
    .DI108 (RAM10_data_in[108] ),    .DI109 (RAM10_data_in[109] ),    .DI110 (RAM10_data_in[110] ),    .DI111 (RAM10_data_in[111] ),
    .DI112 (RAM10_data_in[112] ),    .DI113 (RAM10_data_in[113] ),    .DI114 (RAM10_data_in[114] ),    .DI115 (RAM10_data_in[115] ),
    .DI116 (RAM10_data_in[116] ),    .DI117 (RAM10_data_in[117] ),    .DI118 (RAM10_data_in[118] ),    .DI119 (RAM10_data_in[119] ),
    .DI120 (RAM10_data_in[120] ),    .DI121 (RAM10_data_in[121] ),    .DI122 (RAM10_data_in[122] ),    .DI123 (RAM10_data_in[123] ),
    .DI124 (RAM10_data_in[124] ),    .DI125 (RAM10_data_in[125] ),    .DI126 (RAM10_data_in[126] ),    .DI127 (RAM10_data_in[127] ),

    .A0   (RAM_addr[0]   ),.A1   (RAM_addr[1]   ),.A2   (RAM_addr[2]   ),.A3   (RAM_addr[3]   ),.A4   (RAM_addr[4]   ),.A5   (RAM_addr[5]   ),.A6   (RAM_addr[6]   ),
    .DVSE (1'b0  ),.DVS0 (1'b0  ),.DVS1 (1'b0  ),.DVS2 (1'b0  ),.DVS3 (1'b0  ),
    .WEB0 (~w_WEB10_8[0] ),.WEB1 (~w_WEB10_8[1] ),.WEB2 (~w_WEB10_8[2] ),.WEB3 (~w_WEB10_8[3] ),
    .WEB4 (~w_WEB10_8[4] ),.WEB5 (~w_WEB10_8[5] ),.WEB6 (~w_WEB10_8[6] ),.WEB7 (~w_WEB10_8[7] ),

    .CK    (clka   ),
    .CSB   (1'b0   )
);


SYKB110_128X16X8CM2 u_L2data11_SYKB110_128X16X8CM2(
    .DO0   (RAM11_data_out[128] ),    .DO1   (RAM11_data_out[129] ),    .DO2   (RAM11_data_out[130] ),    .DO3   (RAM11_data_out[131] ),
    .DO4   (RAM11_data_out[132] ),    .DO5   (RAM11_data_out[133] ),    .DO6   (RAM11_data_out[134] ),    .DO7   (RAM11_data_out[135] ),
    .DO8   (RAM11_data_out[136] ),    .DO9   (RAM11_data_out[137] ),    .DO10  (RAM11_data_out[138] ),    .DO11  (RAM11_data_out[139] ),
    .DO12  (RAM11_data_out[140] ),    .DO13  (RAM11_data_out[141] ),    .DO14  (RAM11_data_out[142] ),    .DO15  (RAM11_data_out[143] ),
    .DO16  (RAM11_data_out[144] ),    .DO17  (RAM11_data_out[145] ),    .DO18  (RAM11_data_out[146] ),    .DO19  (RAM11_data_out[147] ),
    .DO20  (RAM11_data_out[148] ),    .DO21  (RAM11_data_out[149] ),    .DO22  (RAM11_data_out[150] ),    .DO23  (RAM11_data_out[151] ),
    .DO24  (RAM11_data_out[152] ),    .DO25  (RAM11_data_out[153] ),    .DO26  (RAM11_data_out[154] ),    .DO27  (RAM11_data_out[155] ),
    .DO28  (RAM11_data_out[156] ),    .DO29  (RAM11_data_out[157] ),    .DO30  (RAM11_data_out[158] ),    .DO31  (RAM11_data_out[159] ),
    .DO32  (RAM11_data_out[160] ),    .DO33  (RAM11_data_out[161] ),    .DO34  (RAM11_data_out[162] ),    .DO35  (RAM11_data_out[163] ),
    .DO36  (RAM11_data_out[164] ),    .DO37  (RAM11_data_out[165] ),    .DO38  (RAM11_data_out[166] ),    .DO39  (RAM11_data_out[167] ),
    .DO40  (RAM11_data_out[168] ),    .DO41  (RAM11_data_out[169] ),    .DO42  (RAM11_data_out[170] ),    .DO43  (RAM11_data_out[171] ),
    .DO44  (RAM11_data_out[172] ),    .DO45  (RAM11_data_out[173] ),    .DO46  (RAM11_data_out[174] ),    .DO47  (RAM11_data_out[175] ),
    .DO48  (RAM11_data_out[176] ),    .DO49  (RAM11_data_out[177] ),    .DO50  (RAM11_data_out[178] ),    .DO51  (RAM11_data_out[179] ),
    .DO52  (RAM11_data_out[180] ),    .DO53  (RAM11_data_out[181] ),    .DO54  (RAM11_data_out[182] ),    .DO55  (RAM11_data_out[183] ),
    .DO56  (RAM11_data_out[184] ),    .DO57  (RAM11_data_out[185] ),    .DO58  (RAM11_data_out[186] ),    .DO59  (RAM11_data_out[187] ),
    .DO60  (RAM11_data_out[188] ),    .DO61  (RAM11_data_out[189] ),    .DO62  (RAM11_data_out[190] ),    .DO63  (RAM11_data_out[191] ),
    .DO64  (RAM11_data_out[192] ),    .DO65  (RAM11_data_out[193] ),    .DO66  (RAM11_data_out[194] ),    .DO67  (RAM11_data_out[195] ),
    .DO68  (RAM11_data_out[196] ),    .DO69  (RAM11_data_out[197] ),    .DO70  (RAM11_data_out[198] ),    .DO71  (RAM11_data_out[199] ),
    .DO72  (RAM11_data_out[200] ),    .DO73  (RAM11_data_out[201] ),    .DO74  (RAM11_data_out[202] ),    .DO75  (RAM11_data_out[203] ),
    .DO76  (RAM11_data_out[204] ),    .DO77  (RAM11_data_out[205] ),    .DO78  (RAM11_data_out[206] ),    .DO79  (RAM11_data_out[207] ),
    .DO80  (RAM11_data_out[208] ),    .DO81  (RAM11_data_out[209] ),    .DO82  (RAM11_data_out[210] ),    .DO83  (RAM11_data_out[211] ),
    .DO84  (RAM11_data_out[212] ),    .DO85  (RAM11_data_out[213] ),    .DO86  (RAM11_data_out[214] ),    .DO87  (RAM11_data_out[215] ),
    .DO88  (RAM11_data_out[216] ),    .DO89  (RAM11_data_out[217] ),    .DO90  (RAM11_data_out[218] ),    .DO91  (RAM11_data_out[219] ),
    .DO92  (RAM11_data_out[220] ),    .DO93  (RAM11_data_out[221] ),    .DO94  (RAM11_data_out[222] ),    .DO95  (RAM11_data_out[223] ),
    .DO96  (RAM11_data_out[224] ),    .DO97  (RAM11_data_out[225] ),    .DO98  (RAM11_data_out[226] ),    .DO99  (RAM11_data_out[227] ),
    .DO100 (RAM11_data_out[228] ),    .DO101 (RAM11_data_out[229] ),    .DO102 (RAM11_data_out[230] ),    .DO103 (RAM11_data_out[231] ),
    .DO104 (RAM11_data_out[232] ),    .DO105 (RAM11_data_out[233] ),    .DO106 (RAM11_data_out[234] ),    .DO107 (RAM11_data_out[235] ),
    .DO108 (RAM11_data_out[236] ),    .DO109 (RAM11_data_out[237] ),    .DO110 (RAM11_data_out[238] ),    .DO111 (RAM11_data_out[239] ),
    .DO112 (RAM11_data_out[240] ),    .DO113 (RAM11_data_out[241] ),    .DO114 (RAM11_data_out[242] ),    .DO115 (RAM11_data_out[243] ),
    .DO116 (RAM11_data_out[244] ),    .DO117 (RAM11_data_out[245] ),    .DO118 (RAM11_data_out[246] ),    .DO119 (RAM11_data_out[247] ),
    .DO120 (RAM11_data_out[248] ),    .DO121 (RAM11_data_out[249] ),    .DO122 (RAM11_data_out[250] ),    .DO123 (RAM11_data_out[251] ),
    .DO124 (RAM11_data_out[252] ),    .DO125 (RAM11_data_out[253] ),    .DO126 (RAM11_data_out[254] ),    .DO127 (RAM11_data_out[255] ),

    .DI0   (RAM11_data_in[128] ),    .DI1   (RAM11_data_in[129] ),    .DI2   (RAM11_data_in[130] ),    .DI3   (RAM11_data_in[131] ),
    .DI4   (RAM11_data_in[132] ),    .DI5   (RAM11_data_in[133] ),    .DI6   (RAM11_data_in[134] ),    .DI7   (RAM11_data_in[135] ),
    .DI8   (RAM11_data_in[136] ),    .DI9   (RAM11_data_in[137] ),    .DI10  (RAM11_data_in[138] ),    .DI11  (RAM11_data_in[139] ),
    .DI12  (RAM11_data_in[140] ),    .DI13  (RAM11_data_in[141] ),    .DI14  (RAM11_data_in[142] ),    .DI15  (RAM11_data_in[143] ),
    .DI16  (RAM11_data_in[144] ),    .DI17  (RAM11_data_in[145] ),    .DI18  (RAM11_data_in[146] ),    .DI19  (RAM11_data_in[147] ),
    .DI20  (RAM11_data_in[148] ),    .DI21  (RAM11_data_in[149] ),    .DI22  (RAM11_data_in[150] ),    .DI23  (RAM11_data_in[151] ),
    .DI24  (RAM11_data_in[152] ),    .DI25  (RAM11_data_in[153] ),    .DI26  (RAM11_data_in[154] ),    .DI27  (RAM11_data_in[155] ),
    .DI28  (RAM11_data_in[156] ),    .DI29  (RAM11_data_in[157] ),    .DI30  (RAM11_data_in[158] ),    .DI31  (RAM11_data_in[159] ),
    .DI32  (RAM11_data_in[160] ),    .DI33  (RAM11_data_in[161] ),    .DI34  (RAM11_data_in[162] ),    .DI35  (RAM11_data_in[163] ),
    .DI36  (RAM11_data_in[164] ),    .DI37  (RAM11_data_in[165] ),    .DI38  (RAM11_data_in[166] ),    .DI39  (RAM11_data_in[167] ),
    .DI40  (RAM11_data_in[168] ),    .DI41  (RAM11_data_in[169] ),    .DI42  (RAM11_data_in[170] ),    .DI43  (RAM11_data_in[171] ),
    .DI44  (RAM11_data_in[172] ),    .DI45  (RAM11_data_in[173] ),    .DI46  (RAM11_data_in[174] ),    .DI47  (RAM11_data_in[175] ),
    .DI48  (RAM11_data_in[176] ),    .DI49  (RAM11_data_in[177] ),    .DI50  (RAM11_data_in[178] ),    .DI51  (RAM11_data_in[179] ),
    .DI52  (RAM11_data_in[180] ),    .DI53  (RAM11_data_in[181] ),    .DI54  (RAM11_data_in[182] ),    .DI55  (RAM11_data_in[183] ),
    .DI56  (RAM11_data_in[184] ),    .DI57  (RAM11_data_in[185] ),    .DI58  (RAM11_data_in[186] ),    .DI59  (RAM11_data_in[187] ),
    .DI60  (RAM11_data_in[188] ),    .DI61  (RAM11_data_in[189] ),    .DI62  (RAM11_data_in[190] ),    .DI63  (RAM11_data_in[191] ),
    .DI64  (RAM11_data_in[192] ),    .DI65  (RAM11_data_in[193] ),    .DI66  (RAM11_data_in[194] ),    .DI67  (RAM11_data_in[195] ),
    .DI68  (RAM11_data_in[196] ),    .DI69  (RAM11_data_in[197] ),    .DI70  (RAM11_data_in[198] ),    .DI71  (RAM11_data_in[199] ),
    .DI72  (RAM11_data_in[200] ),    .DI73  (RAM11_data_in[201] ),    .DI74  (RAM11_data_in[202] ),    .DI75  (RAM11_data_in[203] ),
    .DI76  (RAM11_data_in[204] ),    .DI77  (RAM11_data_in[205] ),    .DI78  (RAM11_data_in[206] ),    .DI79  (RAM11_data_in[207] ),
    .DI80  (RAM11_data_in[208] ),    .DI81  (RAM11_data_in[209] ),    .DI82  (RAM11_data_in[210] ),    .DI83  (RAM11_data_in[211] ),
    .DI84  (RAM11_data_in[212] ),    .DI85  (RAM11_data_in[213] ),    .DI86  (RAM11_data_in[214] ),    .DI87  (RAM11_data_in[215] ),
    .DI88  (RAM11_data_in[216] ),    .DI89  (RAM11_data_in[217] ),    .DI90  (RAM11_data_in[218] ),    .DI91  (RAM11_data_in[219] ),
    .DI92  (RAM11_data_in[220] ),    .DI93  (RAM11_data_in[221] ),    .DI94  (RAM11_data_in[222] ),    .DI95  (RAM11_data_in[223] ),
    .DI96  (RAM11_data_in[224] ),    .DI97  (RAM11_data_in[225] ),    .DI98  (RAM11_data_in[226] ),    .DI99  (RAM11_data_in[227] ),
    .DI100 (RAM11_data_in[228] ),    .DI101 (RAM11_data_in[229] ),    .DI102 (RAM11_data_in[230] ),    .DI103 (RAM11_data_in[231] ),
    .DI104 (RAM11_data_in[232] ),    .DI105 (RAM11_data_in[233] ),    .DI106 (RAM11_data_in[234] ),    .DI107 (RAM11_data_in[235] ),
    .DI108 (RAM11_data_in[236] ),    .DI109 (RAM11_data_in[237] ),    .DI110 (RAM11_data_in[238] ),    .DI111 (RAM11_data_in[239] ),
    .DI112 (RAM11_data_in[240] ),    .DI113 (RAM11_data_in[241] ),    .DI114 (RAM11_data_in[242] ),    .DI115 (RAM11_data_in[243] ),
    .DI116 (RAM11_data_in[244] ),    .DI117 (RAM11_data_in[245] ),    .DI118 (RAM11_data_in[246] ),    .DI119 (RAM11_data_in[247] ),
    .DI120 (RAM11_data_in[248] ),    .DI121 (RAM11_data_in[249] ),    .DI122 (RAM11_data_in[250] ),    .DI123 (RAM11_data_in[251] ),
    .DI124 (RAM11_data_in[252] ),    .DI125 (RAM11_data_in[253] ),    .DI126 (RAM11_data_in[254] ),    .DI127 (RAM11_data_in[255] ),

    .A0   (RAM_addr[0]   ),.A1   (RAM_addr[1]   ),.A2   (RAM_addr[2]   ),.A3   (RAM_addr[3]   ),.A4   (RAM_addr[4]   ),.A5   (RAM_addr[5]   ),.A6   (RAM_addr[6]   ),
    .DVSE (1'b0  ),.DVS0 (1'b0  ),.DVS1 (1'b0  ),.DVS2 (1'b0  ),.DVS3 (1'b0  ),
    .WEB0 (~w_WEB11_8[0] ),.WEB1 (~w_WEB11_8[1] ),.WEB2 (~w_WEB11_8[2] ),.WEB3 (~w_WEB11_8[3] ),
    .WEB4 (~w_WEB11_8[4] ),.WEB5 (~w_WEB11_8[5] ),.WEB6 (~w_WEB11_8[6] ),.WEB7 (~w_WEB11_8[7] ),

    .CK    (clka   ),
    .CSB   (1'b0   )
);


SYKB110_128X16X8CM2 u_L2data12_SYKB110_128X16X8CM2(
    .DO0   (RAM12_data_out[0  ] ),    .DO1   (RAM12_data_out[1  ] ),    .DO2   (RAM12_data_out[2  ] ),    .DO3   (RAM12_data_out[3  ] ),
    .DO4   (RAM12_data_out[4  ] ),    .DO5   (RAM12_data_out[5  ] ),    .DO6   (RAM12_data_out[6  ] ),    .DO7   (RAM12_data_out[7  ] ),
    .DO8   (RAM12_data_out[8  ] ),    .DO9   (RAM12_data_out[9  ] ),    .DO10  (RAM12_data_out[10 ] ),    .DO11  (RAM12_data_out[11 ] ),
    .DO12  (RAM12_data_out[12 ] ),    .DO13  (RAM12_data_out[13 ] ),    .DO14  (RAM12_data_out[14 ] ),    .DO15  (RAM12_data_out[15 ] ),
    .DO16  (RAM12_data_out[16 ] ),    .DO17  (RAM12_data_out[17 ] ),    .DO18  (RAM12_data_out[18 ] ),    .DO19  (RAM12_data_out[19 ] ),
    .DO20  (RAM12_data_out[20 ] ),    .DO21  (RAM12_data_out[21 ] ),    .DO22  (RAM12_data_out[22 ] ),    .DO23  (RAM12_data_out[23 ] ),
    .DO24  (RAM12_data_out[24 ] ),    .DO25  (RAM12_data_out[25 ] ),    .DO26  (RAM12_data_out[26 ] ),    .DO27  (RAM12_data_out[27 ] ),
    .DO28  (RAM12_data_out[28 ] ),    .DO29  (RAM12_data_out[29 ] ),    .DO30  (RAM12_data_out[30 ] ),    .DO31  (RAM12_data_out[31 ] ),
    .DO32  (RAM12_data_out[32 ] ),    .DO33  (RAM12_data_out[33 ] ),    .DO34  (RAM12_data_out[34 ] ),    .DO35  (RAM12_data_out[35 ] ),
    .DO36  (RAM12_data_out[36 ] ),    .DO37  (RAM12_data_out[37 ] ),    .DO38  (RAM12_data_out[38 ] ),    .DO39  (RAM12_data_out[39 ] ),
    .DO40  (RAM12_data_out[40 ] ),    .DO41  (RAM12_data_out[41 ] ),    .DO42  (RAM12_data_out[42 ] ),    .DO43  (RAM12_data_out[43 ] ),
    .DO44  (RAM12_data_out[44 ] ),    .DO45  (RAM12_data_out[45 ] ),    .DO46  (RAM12_data_out[46 ] ),    .DO47  (RAM12_data_out[47 ] ),
    .DO48  (RAM12_data_out[48 ] ),    .DO49  (RAM12_data_out[49 ] ),    .DO50  (RAM12_data_out[50 ] ),    .DO51  (RAM12_data_out[51 ] ),
    .DO52  (RAM12_data_out[52 ] ),    .DO53  (RAM12_data_out[53 ] ),    .DO54  (RAM12_data_out[54 ] ),    .DO55  (RAM12_data_out[55 ] ),
    .DO56  (RAM12_data_out[56 ] ),    .DO57  (RAM12_data_out[57 ] ),    .DO58  (RAM12_data_out[58 ] ),    .DO59  (RAM12_data_out[59 ] ),
    .DO60  (RAM12_data_out[60 ] ),    .DO61  (RAM12_data_out[61 ] ),    .DO62  (RAM12_data_out[62 ] ),    .DO63  (RAM12_data_out[63 ] ),
    .DO64  (RAM12_data_out[64 ] ),    .DO65  (RAM12_data_out[65 ] ),    .DO66  (RAM12_data_out[66 ] ),    .DO67  (RAM12_data_out[67 ] ),
    .DO68  (RAM12_data_out[68 ] ),    .DO69  (RAM12_data_out[69 ] ),    .DO70  (RAM12_data_out[70 ] ),    .DO71  (RAM12_data_out[71 ] ),
    .DO72  (RAM12_data_out[72 ] ),    .DO73  (RAM12_data_out[73 ] ),    .DO74  (RAM12_data_out[74 ] ),    .DO75  (RAM12_data_out[75 ] ),
    .DO76  (RAM12_data_out[76 ] ),    .DO77  (RAM12_data_out[77 ] ),    .DO78  (RAM12_data_out[78 ] ),    .DO79  (RAM12_data_out[79 ] ),
    .DO80  (RAM12_data_out[80 ] ),    .DO81  (RAM12_data_out[81 ] ),    .DO82  (RAM12_data_out[82 ] ),    .DO83  (RAM12_data_out[83 ] ),
    .DO84  (RAM12_data_out[84 ] ),    .DO85  (RAM12_data_out[85 ] ),    .DO86  (RAM12_data_out[86 ] ),    .DO87  (RAM12_data_out[87 ] ),
    .DO88  (RAM12_data_out[88 ] ),    .DO89  (RAM12_data_out[89 ] ),    .DO90  (RAM12_data_out[90 ] ),    .DO91  (RAM12_data_out[91 ] ),
    .DO92  (RAM12_data_out[92 ] ),    .DO93  (RAM12_data_out[93 ] ),    .DO94  (RAM12_data_out[94 ] ),    .DO95  (RAM12_data_out[95 ] ),
    .DO96  (RAM12_data_out[96 ] ),    .DO97  (RAM12_data_out[97 ] ),    .DO98  (RAM12_data_out[98 ] ),    .DO99  (RAM12_data_out[99 ] ),
    .DO100 (RAM12_data_out[100] ),    .DO101 (RAM12_data_out[101] ),    .DO102 (RAM12_data_out[102] ),    .DO103 (RAM12_data_out[103] ),
    .DO104 (RAM12_data_out[104] ),    .DO105 (RAM12_data_out[105] ),    .DO106 (RAM12_data_out[106] ),    .DO107 (RAM12_data_out[107] ),
    .DO108 (RAM12_data_out[108] ),    .DO109 (RAM12_data_out[109] ),    .DO110 (RAM12_data_out[110] ),    .DO111 (RAM12_data_out[111] ),
    .DO112 (RAM12_data_out[112] ),    .DO113 (RAM12_data_out[113] ),    .DO114 (RAM12_data_out[114] ),    .DO115 (RAM12_data_out[115] ),
    .DO116 (RAM12_data_out[116] ),    .DO117 (RAM12_data_out[117] ),    .DO118 (RAM12_data_out[118] ),    .DO119 (RAM12_data_out[119] ),
    .DO120 (RAM12_data_out[120] ),    .DO121 (RAM12_data_out[121] ),    .DO122 (RAM12_data_out[122] ),    .DO123 (RAM12_data_out[123] ),
    .DO124 (RAM12_data_out[124] ),    .DO125 (RAM12_data_out[125] ),    .DO126 (RAM12_data_out[126] ),    .DO127 (RAM12_data_out[127] ),

    .DI0   (RAM12_data_in[0  ] ),    .DI1   (RAM12_data_in[1  ] ),    .DI2   (RAM12_data_in[2  ] ),    .DI3   (RAM12_data_in[3  ] ),
    .DI4   (RAM12_data_in[4  ] ),    .DI5   (RAM12_data_in[5  ] ),    .DI6   (RAM12_data_in[6  ] ),    .DI7   (RAM12_data_in[7  ] ),
    .DI8   (RAM12_data_in[8  ] ),    .DI9   (RAM12_data_in[9  ] ),    .DI10  (RAM12_data_in[10 ] ),    .DI11  (RAM12_data_in[11 ] ),
    .DI12  (RAM12_data_in[12 ] ),    .DI13  (RAM12_data_in[13 ] ),    .DI14  (RAM12_data_in[14 ] ),    .DI15  (RAM12_data_in[15 ] ),
    .DI16  (RAM12_data_in[16 ] ),    .DI17  (RAM12_data_in[17 ] ),    .DI18  (RAM12_data_in[18 ] ),    .DI19  (RAM12_data_in[19 ] ),
    .DI20  (RAM12_data_in[20 ] ),    .DI21  (RAM12_data_in[21 ] ),    .DI22  (RAM12_data_in[22 ] ),    .DI23  (RAM12_data_in[23 ] ),
    .DI24  (RAM12_data_in[24 ] ),    .DI25  (RAM12_data_in[25 ] ),    .DI26  (RAM12_data_in[26 ] ),    .DI27  (RAM12_data_in[27 ] ),
    .DI28  (RAM12_data_in[28 ] ),    .DI29  (RAM12_data_in[29 ] ),    .DI30  (RAM12_data_in[30 ] ),    .DI31  (RAM12_data_in[31 ] ),
    .DI32  (RAM12_data_in[32 ] ),    .DI33  (RAM12_data_in[33 ] ),    .DI34  (RAM12_data_in[34 ] ),    .DI35  (RAM12_data_in[35 ] ),
    .DI36  (RAM12_data_in[36 ] ),    .DI37  (RAM12_data_in[37 ] ),    .DI38  (RAM12_data_in[38 ] ),    .DI39  (RAM12_data_in[39 ] ),
    .DI40  (RAM12_data_in[40 ] ),    .DI41  (RAM12_data_in[41 ] ),    .DI42  (RAM12_data_in[42 ] ),    .DI43  (RAM12_data_in[43 ] ),
    .DI44  (RAM12_data_in[44 ] ),    .DI45  (RAM12_data_in[45 ] ),    .DI46  (RAM12_data_in[46 ] ),    .DI47  (RAM12_data_in[47 ] ),
    .DI48  (RAM12_data_in[48 ] ),    .DI49  (RAM12_data_in[49 ] ),    .DI50  (RAM12_data_in[50 ] ),    .DI51  (RAM12_data_in[51 ] ),
    .DI52  (RAM12_data_in[52 ] ),    .DI53  (RAM12_data_in[53 ] ),    .DI54  (RAM12_data_in[54 ] ),    .DI55  (RAM12_data_in[55 ] ),
    .DI56  (RAM12_data_in[56 ] ),    .DI57  (RAM12_data_in[57 ] ),    .DI58  (RAM12_data_in[58 ] ),    .DI59  (RAM12_data_in[59 ] ),
    .DI60  (RAM12_data_in[60 ] ),    .DI61  (RAM12_data_in[61 ] ),    .DI62  (RAM12_data_in[62 ] ),    .DI63  (RAM12_data_in[63 ] ),
    .DI64  (RAM12_data_in[64 ] ),    .DI65  (RAM12_data_in[65 ] ),    .DI66  (RAM12_data_in[66 ] ),    .DI67  (RAM12_data_in[67 ] ),
    .DI68  (RAM12_data_in[68 ] ),    .DI69  (RAM12_data_in[69 ] ),    .DI70  (RAM12_data_in[70 ] ),    .DI71  (RAM12_data_in[71 ] ),
    .DI72  (RAM12_data_in[72 ] ),    .DI73  (RAM12_data_in[73 ] ),    .DI74  (RAM12_data_in[74 ] ),    .DI75  (RAM12_data_in[75 ] ),
    .DI76  (RAM12_data_in[76 ] ),    .DI77  (RAM12_data_in[77 ] ),    .DI78  (RAM12_data_in[78 ] ),    .DI79  (RAM12_data_in[79 ] ),
    .DI80  (RAM12_data_in[80 ] ),    .DI81  (RAM12_data_in[81 ] ),    .DI82  (RAM12_data_in[82 ] ),    .DI83  (RAM12_data_in[83 ] ),
    .DI84  (RAM12_data_in[84 ] ),    .DI85  (RAM12_data_in[85 ] ),    .DI86  (RAM12_data_in[86 ] ),    .DI87  (RAM12_data_in[87 ] ),
    .DI88  (RAM12_data_in[88 ] ),    .DI89  (RAM12_data_in[89 ] ),    .DI90  (RAM12_data_in[90 ] ),    .DI91  (RAM12_data_in[91 ] ),
    .DI92  (RAM12_data_in[92 ] ),    .DI93  (RAM12_data_in[93 ] ),    .DI94  (RAM12_data_in[94 ] ),    .DI95  (RAM12_data_in[95 ] ),
    .DI96  (RAM12_data_in[96 ] ),    .DI97  (RAM12_data_in[97 ] ),    .DI98  (RAM12_data_in[98 ] ),    .DI99  (RAM12_data_in[99 ] ),
    .DI100 (RAM12_data_in[100] ),    .DI101 (RAM12_data_in[101] ),    .DI102 (RAM12_data_in[102] ),    .DI103 (RAM12_data_in[103] ),
    .DI104 (RAM12_data_in[104] ),    .DI105 (RAM12_data_in[105] ),    .DI106 (RAM12_data_in[106] ),    .DI107 (RAM12_data_in[107] ),
    .DI108 (RAM12_data_in[108] ),    .DI109 (RAM12_data_in[109] ),    .DI110 (RAM12_data_in[110] ),    .DI111 (RAM12_data_in[111] ),
    .DI112 (RAM12_data_in[112] ),    .DI113 (RAM12_data_in[113] ),    .DI114 (RAM12_data_in[114] ),    .DI115 (RAM12_data_in[115] ),
    .DI116 (RAM12_data_in[116] ),    .DI117 (RAM12_data_in[117] ),    .DI118 (RAM12_data_in[118] ),    .DI119 (RAM12_data_in[119] ),
    .DI120 (RAM12_data_in[120] ),    .DI121 (RAM12_data_in[121] ),    .DI122 (RAM12_data_in[122] ),    .DI123 (RAM12_data_in[123] ),
    .DI124 (RAM12_data_in[124] ),    .DI125 (RAM12_data_in[125] ),    .DI126 (RAM12_data_in[126] ),    .DI127 (RAM12_data_in[127] ),

    .A0   (RAM_addr[0]   ),.A1   (RAM_addr[1]   ),.A2   (RAM_addr[2]   ),.A3   (RAM_addr[3]   ),.A4   (RAM_addr[4]   ),.A5   (RAM_addr[5]   ),.A6   (RAM_addr[6]   ),
    .DVSE (1'b0  ),.DVS0 (1'b0  ),.DVS1 (1'b0  ),.DVS2 (1'b0  ),.DVS3 (1'b0  ),
    .WEB0 (~w_WEB12_8[0] ),.WEB1 (~w_WEB12_8[1] ),.WEB2 (~w_WEB12_8[2] ),.WEB3 (~w_WEB12_8[3] ),
    .WEB4 (~w_WEB12_8[4] ),.WEB5 (~w_WEB12_8[5] ),.WEB6 (~w_WEB12_8[6] ),.WEB7 (~w_WEB12_8[7] ),

    .CK    (clka   ),
    .CSB   (1'b0   )
);


SYKB110_128X16X8CM2 u_L2data13_SYKB110_128X16X8CM2(
    .DO0   (RAM13_data_out[128] ),    .DO1   (RAM13_data_out[129] ),    .DO2   (RAM13_data_out[130] ),    .DO3   (RAM13_data_out[131] ),
    .DO4   (RAM13_data_out[132] ),    .DO5   (RAM13_data_out[133] ),    .DO6   (RAM13_data_out[134] ),    .DO7   (RAM13_data_out[135] ),
    .DO8   (RAM13_data_out[136] ),    .DO9   (RAM13_data_out[137] ),    .DO10  (RAM13_data_out[138] ),    .DO11  (RAM13_data_out[139] ),
    .DO12  (RAM13_data_out[140] ),    .DO13  (RAM13_data_out[141] ),    .DO14  (RAM13_data_out[142] ),    .DO15  (RAM13_data_out[143] ),
    .DO16  (RAM13_data_out[144] ),    .DO17  (RAM13_data_out[145] ),    .DO18  (RAM13_data_out[146] ),    .DO19  (RAM13_data_out[147] ),
    .DO20  (RAM13_data_out[148] ),    .DO21  (RAM13_data_out[149] ),    .DO22  (RAM13_data_out[150] ),    .DO23  (RAM13_data_out[151] ),
    .DO24  (RAM13_data_out[152] ),    .DO25  (RAM13_data_out[153] ),    .DO26  (RAM13_data_out[154] ),    .DO27  (RAM13_data_out[155] ),
    .DO28  (RAM13_data_out[156] ),    .DO29  (RAM13_data_out[157] ),    .DO30  (RAM13_data_out[158] ),    .DO31  (RAM13_data_out[159] ),
    .DO32  (RAM13_data_out[160] ),    .DO33  (RAM13_data_out[161] ),    .DO34  (RAM13_data_out[162] ),    .DO35  (RAM13_data_out[163] ),
    .DO36  (RAM13_data_out[164] ),    .DO37  (RAM13_data_out[165] ),    .DO38  (RAM13_data_out[166] ),    .DO39  (RAM13_data_out[167] ),
    .DO40  (RAM13_data_out[168] ),    .DO41  (RAM13_data_out[169] ),    .DO42  (RAM13_data_out[170] ),    .DO43  (RAM13_data_out[171] ),
    .DO44  (RAM13_data_out[172] ),    .DO45  (RAM13_data_out[173] ),    .DO46  (RAM13_data_out[174] ),    .DO47  (RAM13_data_out[175] ),
    .DO48  (RAM13_data_out[176] ),    .DO49  (RAM13_data_out[177] ),    .DO50  (RAM13_data_out[178] ),    .DO51  (RAM13_data_out[179] ),
    .DO52  (RAM13_data_out[180] ),    .DO53  (RAM13_data_out[181] ),    .DO54  (RAM13_data_out[182] ),    .DO55  (RAM13_data_out[183] ),
    .DO56  (RAM13_data_out[184] ),    .DO57  (RAM13_data_out[185] ),    .DO58  (RAM13_data_out[186] ),    .DO59  (RAM13_data_out[187] ),
    .DO60  (RAM13_data_out[188] ),    .DO61  (RAM13_data_out[189] ),    .DO62  (RAM13_data_out[190] ),    .DO63  (RAM13_data_out[191] ),
    .DO64  (RAM13_data_out[192] ),    .DO65  (RAM13_data_out[193] ),    .DO66  (RAM13_data_out[194] ),    .DO67  (RAM13_data_out[195] ),
    .DO68  (RAM13_data_out[196] ),    .DO69  (RAM13_data_out[197] ),    .DO70  (RAM13_data_out[198] ),    .DO71  (RAM13_data_out[199] ),
    .DO72  (RAM13_data_out[200] ),    .DO73  (RAM13_data_out[201] ),    .DO74  (RAM13_data_out[202] ),    .DO75  (RAM13_data_out[203] ),
    .DO76  (RAM13_data_out[204] ),    .DO77  (RAM13_data_out[205] ),    .DO78  (RAM13_data_out[206] ),    .DO79  (RAM13_data_out[207] ),
    .DO80  (RAM13_data_out[208] ),    .DO81  (RAM13_data_out[209] ),    .DO82  (RAM13_data_out[210] ),    .DO83  (RAM13_data_out[211] ),
    .DO84  (RAM13_data_out[212] ),    .DO85  (RAM13_data_out[213] ),    .DO86  (RAM13_data_out[214] ),    .DO87  (RAM13_data_out[215] ),
    .DO88  (RAM13_data_out[216] ),    .DO89  (RAM13_data_out[217] ),    .DO90  (RAM13_data_out[218] ),    .DO91  (RAM13_data_out[219] ),
    .DO92  (RAM13_data_out[220] ),    .DO93  (RAM13_data_out[221] ),    .DO94  (RAM13_data_out[222] ),    .DO95  (RAM13_data_out[223] ),
    .DO96  (RAM13_data_out[224] ),    .DO97  (RAM13_data_out[225] ),    .DO98  (RAM13_data_out[226] ),    .DO99  (RAM13_data_out[227] ),
    .DO100 (RAM13_data_out[228] ),    .DO101 (RAM13_data_out[229] ),    .DO102 (RAM13_data_out[230] ),    .DO103 (RAM13_data_out[231] ),
    .DO104 (RAM13_data_out[232] ),    .DO105 (RAM13_data_out[233] ),    .DO106 (RAM13_data_out[234] ),    .DO107 (RAM13_data_out[235] ),
    .DO108 (RAM13_data_out[236] ),    .DO109 (RAM13_data_out[237] ),    .DO110 (RAM13_data_out[238] ),    .DO111 (RAM13_data_out[239] ),
    .DO112 (RAM13_data_out[240] ),    .DO113 (RAM13_data_out[241] ),    .DO114 (RAM13_data_out[242] ),    .DO115 (RAM13_data_out[243] ),
    .DO116 (RAM13_data_out[244] ),    .DO117 (RAM13_data_out[245] ),    .DO118 (RAM13_data_out[246] ),    .DO119 (RAM13_data_out[247] ),
    .DO120 (RAM13_data_out[248] ),    .DO121 (RAM13_data_out[249] ),    .DO122 (RAM13_data_out[250] ),    .DO123 (RAM13_data_out[251] ),
    .DO124 (RAM13_data_out[252] ),    .DO125 (RAM13_data_out[253] ),    .DO126 (RAM13_data_out[254] ),    .DO127 (RAM13_data_out[255] ),

    .DI0   (RAM13_data_in[128] ),    .DI1   (RAM13_data_in[129] ),    .DI2   (RAM13_data_in[130] ),    .DI3   (RAM13_data_in[131] ),
    .DI4   (RAM13_data_in[132] ),    .DI5   (RAM13_data_in[133] ),    .DI6   (RAM13_data_in[134] ),    .DI7   (RAM13_data_in[135] ),
    .DI8   (RAM13_data_in[136] ),    .DI9   (RAM13_data_in[137] ),    .DI10  (RAM13_data_in[138] ),    .DI11  (RAM13_data_in[139] ),
    .DI12  (RAM13_data_in[140] ),    .DI13  (RAM13_data_in[141] ),    .DI14  (RAM13_data_in[142] ),    .DI15  (RAM13_data_in[143] ),
    .DI16  (RAM13_data_in[144] ),    .DI17  (RAM13_data_in[145] ),    .DI18  (RAM13_data_in[146] ),    .DI19  (RAM13_data_in[147] ),
    .DI20  (RAM13_data_in[148] ),    .DI21  (RAM13_data_in[149] ),    .DI22  (RAM13_data_in[150] ),    .DI23  (RAM13_data_in[151] ),
    .DI24  (RAM13_data_in[152] ),    .DI25  (RAM13_data_in[153] ),    .DI26  (RAM13_data_in[154] ),    .DI27  (RAM13_data_in[155] ),
    .DI28  (RAM13_data_in[156] ),    .DI29  (RAM13_data_in[157] ),    .DI30  (RAM13_data_in[158] ),    .DI31  (RAM13_data_in[159] ),
    .DI32  (RAM13_data_in[160] ),    .DI33  (RAM13_data_in[161] ),    .DI34  (RAM13_data_in[162] ),    .DI35  (RAM13_data_in[163] ),
    .DI36  (RAM13_data_in[164] ),    .DI37  (RAM13_data_in[165] ),    .DI38  (RAM13_data_in[166] ),    .DI39  (RAM13_data_in[167] ),
    .DI40  (RAM13_data_in[168] ),    .DI41  (RAM13_data_in[169] ),    .DI42  (RAM13_data_in[170] ),    .DI43  (RAM13_data_in[171] ),
    .DI44  (RAM13_data_in[172] ),    .DI45  (RAM13_data_in[173] ),    .DI46  (RAM13_data_in[174] ),    .DI47  (RAM13_data_in[175] ),
    .DI48  (RAM13_data_in[176] ),    .DI49  (RAM13_data_in[177] ),    .DI50  (RAM13_data_in[178] ),    .DI51  (RAM13_data_in[179] ),
    .DI52  (RAM13_data_in[180] ),    .DI53  (RAM13_data_in[181] ),    .DI54  (RAM13_data_in[182] ),    .DI55  (RAM13_data_in[183] ),
    .DI56  (RAM13_data_in[184] ),    .DI57  (RAM13_data_in[185] ),    .DI58  (RAM13_data_in[186] ),    .DI59  (RAM13_data_in[187] ),
    .DI60  (RAM13_data_in[188] ),    .DI61  (RAM13_data_in[189] ),    .DI62  (RAM13_data_in[190] ),    .DI63  (RAM13_data_in[191] ),
    .DI64  (RAM13_data_in[192] ),    .DI65  (RAM13_data_in[193] ),    .DI66  (RAM13_data_in[194] ),    .DI67  (RAM13_data_in[195] ),
    .DI68  (RAM13_data_in[196] ),    .DI69  (RAM13_data_in[197] ),    .DI70  (RAM13_data_in[198] ),    .DI71  (RAM13_data_in[199] ),
    .DI72  (RAM13_data_in[200] ),    .DI73  (RAM13_data_in[201] ),    .DI74  (RAM13_data_in[202] ),    .DI75  (RAM13_data_in[203] ),
    .DI76  (RAM13_data_in[204] ),    .DI77  (RAM13_data_in[205] ),    .DI78  (RAM13_data_in[206] ),    .DI79  (RAM13_data_in[207] ),
    .DI80  (RAM13_data_in[208] ),    .DI81  (RAM13_data_in[209] ),    .DI82  (RAM13_data_in[210] ),    .DI83  (RAM13_data_in[211] ),
    .DI84  (RAM13_data_in[212] ),    .DI85  (RAM13_data_in[213] ),    .DI86  (RAM13_data_in[214] ),    .DI87  (RAM13_data_in[215] ),
    .DI88  (RAM13_data_in[216] ),    .DI89  (RAM13_data_in[217] ),    .DI90  (RAM13_data_in[218] ),    .DI91  (RAM13_data_in[219] ),
    .DI92  (RAM13_data_in[220] ),    .DI93  (RAM13_data_in[221] ),    .DI94  (RAM13_data_in[222] ),    .DI95  (RAM13_data_in[223] ),
    .DI96  (RAM13_data_in[224] ),    .DI97  (RAM13_data_in[225] ),    .DI98  (RAM13_data_in[226] ),    .DI99  (RAM13_data_in[227] ),
    .DI100 (RAM13_data_in[228] ),    .DI101 (RAM13_data_in[229] ),    .DI102 (RAM13_data_in[230] ),    .DI103 (RAM13_data_in[231] ),
    .DI104 (RAM13_data_in[232] ),    .DI105 (RAM13_data_in[233] ),    .DI106 (RAM13_data_in[234] ),    .DI107 (RAM13_data_in[235] ),
    .DI108 (RAM13_data_in[236] ),    .DI109 (RAM13_data_in[237] ),    .DI110 (RAM13_data_in[238] ),    .DI111 (RAM13_data_in[239] ),
    .DI112 (RAM13_data_in[240] ),    .DI113 (RAM13_data_in[241] ),    .DI114 (RAM13_data_in[242] ),    .DI115 (RAM13_data_in[243] ),
    .DI116 (RAM13_data_in[244] ),    .DI117 (RAM13_data_in[245] ),    .DI118 (RAM13_data_in[246] ),    .DI119 (RAM13_data_in[247] ),
    .DI120 (RAM13_data_in[248] ),    .DI121 (RAM13_data_in[249] ),    .DI122 (RAM13_data_in[250] ),    .DI123 (RAM13_data_in[251] ),
    .DI124 (RAM13_data_in[252] ),    .DI125 (RAM13_data_in[253] ),    .DI126 (RAM13_data_in[254] ),    .DI127 (RAM13_data_in[255] ),

    .A0   (RAM_addr[0]   ),.A1   (RAM_addr[1]   ),.A2   (RAM_addr[2]   ),.A3   (RAM_addr[3]   ),.A4   (RAM_addr[4]   ),.A5   (RAM_addr[5]   ),.A6   (RAM_addr[6]   ),
    .DVSE (1'b0  ),.DVS0 (1'b0  ),.DVS1 (1'b0  ),.DVS2 (1'b0  ),.DVS3 (1'b0  ),
    .WEB0 (~w_WEB13_8[0] ),.WEB1 (~w_WEB13_8[1] ),.WEB2 (~w_WEB13_8[2] ),.WEB3 (~w_WEB13_8[3] ),
    .WEB4 (~w_WEB13_8[4] ),.WEB5 (~w_WEB13_8[5] ),.WEB6 (~w_WEB13_8[6] ),.WEB7 (~w_WEB13_8[7] ),

    .CK    (clka   ),
    .CSB   (1'b0   )
);


SYKB110_128X16X8CM2 u_L2data14_SYKB110_128X16X8CM2(
    .DO0   (RAM14_data_out[0  ] ),    .DO1   (RAM14_data_out[1  ] ),    .DO2   (RAM14_data_out[2  ] ),    .DO3   (RAM14_data_out[3  ] ),
    .DO4   (RAM14_data_out[4  ] ),    .DO5   (RAM14_data_out[5  ] ),    .DO6   (RAM14_data_out[6  ] ),    .DO7   (RAM14_data_out[7  ] ),
    .DO8   (RAM14_data_out[8  ] ),    .DO9   (RAM14_data_out[9  ] ),    .DO10  (RAM14_data_out[10 ] ),    .DO11  (RAM14_data_out[11 ] ),
    .DO12  (RAM14_data_out[12 ] ),    .DO13  (RAM14_data_out[13 ] ),    .DO14  (RAM14_data_out[14 ] ),    .DO15  (RAM14_data_out[15 ] ),
    .DO16  (RAM14_data_out[16 ] ),    .DO17  (RAM14_data_out[17 ] ),    .DO18  (RAM14_data_out[18 ] ),    .DO19  (RAM14_data_out[19 ] ),
    .DO20  (RAM14_data_out[20 ] ),    .DO21  (RAM14_data_out[21 ] ),    .DO22  (RAM14_data_out[22 ] ),    .DO23  (RAM14_data_out[23 ] ),
    .DO24  (RAM14_data_out[24 ] ),    .DO25  (RAM14_data_out[25 ] ),    .DO26  (RAM14_data_out[26 ] ),    .DO27  (RAM14_data_out[27 ] ),
    .DO28  (RAM14_data_out[28 ] ),    .DO29  (RAM14_data_out[29 ] ),    .DO30  (RAM14_data_out[30 ] ),    .DO31  (RAM14_data_out[31 ] ),
    .DO32  (RAM14_data_out[32 ] ),    .DO33  (RAM14_data_out[33 ] ),    .DO34  (RAM14_data_out[34 ] ),    .DO35  (RAM14_data_out[35 ] ),
    .DO36  (RAM14_data_out[36 ] ),    .DO37  (RAM14_data_out[37 ] ),    .DO38  (RAM14_data_out[38 ] ),    .DO39  (RAM14_data_out[39 ] ),
    .DO40  (RAM14_data_out[40 ] ),    .DO41  (RAM14_data_out[41 ] ),    .DO42  (RAM14_data_out[42 ] ),    .DO43  (RAM14_data_out[43 ] ),
    .DO44  (RAM14_data_out[44 ] ),    .DO45  (RAM14_data_out[45 ] ),    .DO46  (RAM14_data_out[46 ] ),    .DO47  (RAM14_data_out[47 ] ),
    .DO48  (RAM14_data_out[48 ] ),    .DO49  (RAM14_data_out[49 ] ),    .DO50  (RAM14_data_out[50 ] ),    .DO51  (RAM14_data_out[51 ] ),
    .DO52  (RAM14_data_out[52 ] ),    .DO53  (RAM14_data_out[53 ] ),    .DO54  (RAM14_data_out[54 ] ),    .DO55  (RAM14_data_out[55 ] ),
    .DO56  (RAM14_data_out[56 ] ),    .DO57  (RAM14_data_out[57 ] ),    .DO58  (RAM14_data_out[58 ] ),    .DO59  (RAM14_data_out[59 ] ),
    .DO60  (RAM14_data_out[60 ] ),    .DO61  (RAM14_data_out[61 ] ),    .DO62  (RAM14_data_out[62 ] ),    .DO63  (RAM14_data_out[63 ] ),
    .DO64  (RAM14_data_out[64 ] ),    .DO65  (RAM14_data_out[65 ] ),    .DO66  (RAM14_data_out[66 ] ),    .DO67  (RAM14_data_out[67 ] ),
    .DO68  (RAM14_data_out[68 ] ),    .DO69  (RAM14_data_out[69 ] ),    .DO70  (RAM14_data_out[70 ] ),    .DO71  (RAM14_data_out[71 ] ),
    .DO72  (RAM14_data_out[72 ] ),    .DO73  (RAM14_data_out[73 ] ),    .DO74  (RAM14_data_out[74 ] ),    .DO75  (RAM14_data_out[75 ] ),
    .DO76  (RAM14_data_out[76 ] ),    .DO77  (RAM14_data_out[77 ] ),    .DO78  (RAM14_data_out[78 ] ),    .DO79  (RAM14_data_out[79 ] ),
    .DO80  (RAM14_data_out[80 ] ),    .DO81  (RAM14_data_out[81 ] ),    .DO82  (RAM14_data_out[82 ] ),    .DO83  (RAM14_data_out[83 ] ),
    .DO84  (RAM14_data_out[84 ] ),    .DO85  (RAM14_data_out[85 ] ),    .DO86  (RAM14_data_out[86 ] ),    .DO87  (RAM14_data_out[87 ] ),
    .DO88  (RAM14_data_out[88 ] ),    .DO89  (RAM14_data_out[89 ] ),    .DO90  (RAM14_data_out[90 ] ),    .DO91  (RAM14_data_out[91 ] ),
    .DO92  (RAM14_data_out[92 ] ),    .DO93  (RAM14_data_out[93 ] ),    .DO94  (RAM14_data_out[94 ] ),    .DO95  (RAM14_data_out[95 ] ),
    .DO96  (RAM14_data_out[96 ] ),    .DO97  (RAM14_data_out[97 ] ),    .DO98  (RAM14_data_out[98 ] ),    .DO99  (RAM14_data_out[99 ] ),
    .DO100 (RAM14_data_out[100] ),    .DO101 (RAM14_data_out[101] ),    .DO102 (RAM14_data_out[102] ),    .DO103 (RAM14_data_out[103] ),
    .DO104 (RAM14_data_out[104] ),    .DO105 (RAM14_data_out[105] ),    .DO106 (RAM14_data_out[106] ),    .DO107 (RAM14_data_out[107] ),
    .DO108 (RAM14_data_out[108] ),    .DO109 (RAM14_data_out[109] ),    .DO110 (RAM14_data_out[110] ),    .DO111 (RAM14_data_out[111] ),
    .DO112 (RAM14_data_out[112] ),    .DO113 (RAM14_data_out[113] ),    .DO114 (RAM14_data_out[114] ),    .DO115 (RAM14_data_out[115] ),
    .DO116 (RAM14_data_out[116] ),    .DO117 (RAM14_data_out[117] ),    .DO118 (RAM14_data_out[118] ),    .DO119 (RAM14_data_out[119] ),
    .DO120 (RAM14_data_out[120] ),    .DO121 (RAM14_data_out[121] ),    .DO122 (RAM14_data_out[122] ),    .DO123 (RAM14_data_out[123] ),
    .DO124 (RAM14_data_out[124] ),    .DO125 (RAM14_data_out[125] ),    .DO126 (RAM14_data_out[126] ),    .DO127 (RAM14_data_out[127] ),

    .DI0   (RAM14_data_in[0  ] ),    .DI1   (RAM14_data_in[1  ] ),    .DI2   (RAM14_data_in[2  ] ),    .DI3   (RAM14_data_in[3  ] ),
    .DI4   (RAM14_data_in[4  ] ),    .DI5   (RAM14_data_in[5  ] ),    .DI6   (RAM14_data_in[6  ] ),    .DI7   (RAM14_data_in[7  ] ),
    .DI8   (RAM14_data_in[8  ] ),    .DI9   (RAM14_data_in[9  ] ),    .DI10  (RAM14_data_in[10 ] ),    .DI11  (RAM14_data_in[11 ] ),
    .DI12  (RAM14_data_in[12 ] ),    .DI13  (RAM14_data_in[13 ] ),    .DI14  (RAM14_data_in[14 ] ),    .DI15  (RAM14_data_in[15 ] ),
    .DI16  (RAM14_data_in[16 ] ),    .DI17  (RAM14_data_in[17 ] ),    .DI18  (RAM14_data_in[18 ] ),    .DI19  (RAM14_data_in[19 ] ),
    .DI20  (RAM14_data_in[20 ] ),    .DI21  (RAM14_data_in[21 ] ),    .DI22  (RAM14_data_in[22 ] ),    .DI23  (RAM14_data_in[23 ] ),
    .DI24  (RAM14_data_in[24 ] ),    .DI25  (RAM14_data_in[25 ] ),    .DI26  (RAM14_data_in[26 ] ),    .DI27  (RAM14_data_in[27 ] ),
    .DI28  (RAM14_data_in[28 ] ),    .DI29  (RAM14_data_in[29 ] ),    .DI30  (RAM14_data_in[30 ] ),    .DI31  (RAM14_data_in[31 ] ),
    .DI32  (RAM14_data_in[32 ] ),    .DI33  (RAM14_data_in[33 ] ),    .DI34  (RAM14_data_in[34 ] ),    .DI35  (RAM14_data_in[35 ] ),
    .DI36  (RAM14_data_in[36 ] ),    .DI37  (RAM14_data_in[37 ] ),    .DI38  (RAM14_data_in[38 ] ),    .DI39  (RAM14_data_in[39 ] ),
    .DI40  (RAM14_data_in[40 ] ),    .DI41  (RAM14_data_in[41 ] ),    .DI42  (RAM14_data_in[42 ] ),    .DI43  (RAM14_data_in[43 ] ),
    .DI44  (RAM14_data_in[44 ] ),    .DI45  (RAM14_data_in[45 ] ),    .DI46  (RAM14_data_in[46 ] ),    .DI47  (RAM14_data_in[47 ] ),
    .DI48  (RAM14_data_in[48 ] ),    .DI49  (RAM14_data_in[49 ] ),    .DI50  (RAM14_data_in[50 ] ),    .DI51  (RAM14_data_in[51 ] ),
    .DI52  (RAM14_data_in[52 ] ),    .DI53  (RAM14_data_in[53 ] ),    .DI54  (RAM14_data_in[54 ] ),    .DI55  (RAM14_data_in[55 ] ),
    .DI56  (RAM14_data_in[56 ] ),    .DI57  (RAM14_data_in[57 ] ),    .DI58  (RAM14_data_in[58 ] ),    .DI59  (RAM14_data_in[59 ] ),
    .DI60  (RAM14_data_in[60 ] ),    .DI61  (RAM14_data_in[61 ] ),    .DI62  (RAM14_data_in[62 ] ),    .DI63  (RAM14_data_in[63 ] ),
    .DI64  (RAM14_data_in[64 ] ),    .DI65  (RAM14_data_in[65 ] ),    .DI66  (RAM14_data_in[66 ] ),    .DI67  (RAM14_data_in[67 ] ),
    .DI68  (RAM14_data_in[68 ] ),    .DI69  (RAM14_data_in[69 ] ),    .DI70  (RAM14_data_in[70 ] ),    .DI71  (RAM14_data_in[71 ] ),
    .DI72  (RAM14_data_in[72 ] ),    .DI73  (RAM14_data_in[73 ] ),    .DI74  (RAM14_data_in[74 ] ),    .DI75  (RAM14_data_in[75 ] ),
    .DI76  (RAM14_data_in[76 ] ),    .DI77  (RAM14_data_in[77 ] ),    .DI78  (RAM14_data_in[78 ] ),    .DI79  (RAM14_data_in[79 ] ),
    .DI80  (RAM14_data_in[80 ] ),    .DI81  (RAM14_data_in[81 ] ),    .DI82  (RAM14_data_in[82 ] ),    .DI83  (RAM14_data_in[83 ] ),
    .DI84  (RAM14_data_in[84 ] ),    .DI85  (RAM14_data_in[85 ] ),    .DI86  (RAM14_data_in[86 ] ),    .DI87  (RAM14_data_in[87 ] ),
    .DI88  (RAM14_data_in[88 ] ),    .DI89  (RAM14_data_in[89 ] ),    .DI90  (RAM14_data_in[90 ] ),    .DI91  (RAM14_data_in[91 ] ),
    .DI92  (RAM14_data_in[92 ] ),    .DI93  (RAM14_data_in[93 ] ),    .DI94  (RAM14_data_in[94 ] ),    .DI95  (RAM14_data_in[95 ] ),
    .DI96  (RAM14_data_in[96 ] ),    .DI97  (RAM14_data_in[97 ] ),    .DI98  (RAM14_data_in[98 ] ),    .DI99  (RAM14_data_in[99 ] ),
    .DI100 (RAM14_data_in[100] ),    .DI101 (RAM14_data_in[101] ),    .DI102 (RAM14_data_in[102] ),    .DI103 (RAM14_data_in[103] ),
    .DI104 (RAM14_data_in[104] ),    .DI105 (RAM14_data_in[105] ),    .DI106 (RAM14_data_in[106] ),    .DI107 (RAM14_data_in[107] ),
    .DI108 (RAM14_data_in[108] ),    .DI109 (RAM14_data_in[109] ),    .DI110 (RAM14_data_in[110] ),    .DI111 (RAM14_data_in[111] ),
    .DI112 (RAM14_data_in[112] ),    .DI113 (RAM14_data_in[113] ),    .DI114 (RAM14_data_in[114] ),    .DI115 (RAM14_data_in[115] ),
    .DI116 (RAM14_data_in[116] ),    .DI117 (RAM14_data_in[117] ),    .DI118 (RAM14_data_in[118] ),    .DI119 (RAM14_data_in[119] ),
    .DI120 (RAM14_data_in[120] ),    .DI121 (RAM14_data_in[121] ),    .DI122 (RAM14_data_in[122] ),    .DI123 (RAM14_data_in[123] ),
    .DI124 (RAM14_data_in[124] ),    .DI125 (RAM14_data_in[125] ),    .DI126 (RAM14_data_in[126] ),    .DI127 (RAM14_data_in[127] ),

    .A0   (RAM_addr[0]   ),.A1   (RAM_addr[1]   ),.A2   (RAM_addr[2]   ),.A3   (RAM_addr[3]   ),.A4   (RAM_addr[4]   ),.A5   (RAM_addr[5]   ),.A6   (RAM_addr[6]   ),
    .DVSE (1'b0  ),.DVS0 (1'b0  ),.DVS1 (1'b0  ),.DVS2 (1'b0  ),.DVS3 (1'b0  ),
    .WEB0 (~w_WEB14_8[0] ),.WEB1 (~w_WEB14_8[1] ),.WEB2 (~w_WEB14_8[2] ),.WEB3 (~w_WEB14_8[3] ),
    .WEB4 (~w_WEB14_8[4] ),.WEB5 (~w_WEB14_8[5] ),.WEB6 (~w_WEB14_8[6] ),.WEB7 (~w_WEB14_8[7] ),

    .CK    (clka   ),
    .CSB   (1'b0   )
);


SYKB110_128X16X8CM2 u_L2data15_SYKB110_128X16X8CM2(
    .DO0   (RAM15_data_out[128] ),    .DO1   (RAM15_data_out[129] ),    .DO2   (RAM15_data_out[130] ),    .DO3   (RAM15_data_out[131] ),
    .DO4   (RAM15_data_out[132] ),    .DO5   (RAM15_data_out[133] ),    .DO6   (RAM15_data_out[134] ),    .DO7   (RAM15_data_out[135] ),
    .DO8   (RAM15_data_out[136] ),    .DO9   (RAM15_data_out[137] ),    .DO10  (RAM15_data_out[138] ),    .DO11  (RAM15_data_out[139] ),
    .DO12  (RAM15_data_out[140] ),    .DO13  (RAM15_data_out[141] ),    .DO14  (RAM15_data_out[142] ),    .DO15  (RAM15_data_out[143] ),
    .DO16  (RAM15_data_out[144] ),    .DO17  (RAM15_data_out[145] ),    .DO18  (RAM15_data_out[146] ),    .DO19  (RAM15_data_out[147] ),
    .DO20  (RAM15_data_out[148] ),    .DO21  (RAM15_data_out[149] ),    .DO22  (RAM15_data_out[150] ),    .DO23  (RAM15_data_out[151] ),
    .DO24  (RAM15_data_out[152] ),    .DO25  (RAM15_data_out[153] ),    .DO26  (RAM15_data_out[154] ),    .DO27  (RAM15_data_out[155] ),
    .DO28  (RAM15_data_out[156] ),    .DO29  (RAM15_data_out[157] ),    .DO30  (RAM15_data_out[158] ),    .DO31  (RAM15_data_out[159] ),
    .DO32  (RAM15_data_out[160] ),    .DO33  (RAM15_data_out[161] ),    .DO34  (RAM15_data_out[162] ),    .DO35  (RAM15_data_out[163] ),
    .DO36  (RAM15_data_out[164] ),    .DO37  (RAM15_data_out[165] ),    .DO38  (RAM15_data_out[166] ),    .DO39  (RAM15_data_out[167] ),
    .DO40  (RAM15_data_out[168] ),    .DO41  (RAM15_data_out[169] ),    .DO42  (RAM15_data_out[170] ),    .DO43  (RAM15_data_out[171] ),
    .DO44  (RAM15_data_out[172] ),    .DO45  (RAM15_data_out[173] ),    .DO46  (RAM15_data_out[174] ),    .DO47  (RAM15_data_out[175] ),
    .DO48  (RAM15_data_out[176] ),    .DO49  (RAM15_data_out[177] ),    .DO50  (RAM15_data_out[178] ),    .DO51  (RAM15_data_out[179] ),
    .DO52  (RAM15_data_out[180] ),    .DO53  (RAM15_data_out[181] ),    .DO54  (RAM15_data_out[182] ),    .DO55  (RAM15_data_out[183] ),
    .DO56  (RAM15_data_out[184] ),    .DO57  (RAM15_data_out[185] ),    .DO58  (RAM15_data_out[186] ),    .DO59  (RAM15_data_out[187] ),
    .DO60  (RAM15_data_out[188] ),    .DO61  (RAM15_data_out[189] ),    .DO62  (RAM15_data_out[190] ),    .DO63  (RAM15_data_out[191] ),
    .DO64  (RAM15_data_out[192] ),    .DO65  (RAM15_data_out[193] ),    .DO66  (RAM15_data_out[194] ),    .DO67  (RAM15_data_out[195] ),
    .DO68  (RAM15_data_out[196] ),    .DO69  (RAM15_data_out[197] ),    .DO70  (RAM15_data_out[198] ),    .DO71  (RAM15_data_out[199] ),
    .DO72  (RAM15_data_out[200] ),    .DO73  (RAM15_data_out[201] ),    .DO74  (RAM15_data_out[202] ),    .DO75  (RAM15_data_out[203] ),
    .DO76  (RAM15_data_out[204] ),    .DO77  (RAM15_data_out[205] ),    .DO78  (RAM15_data_out[206] ),    .DO79  (RAM15_data_out[207] ),
    .DO80  (RAM15_data_out[208] ),    .DO81  (RAM15_data_out[209] ),    .DO82  (RAM15_data_out[210] ),    .DO83  (RAM15_data_out[211] ),
    .DO84  (RAM15_data_out[212] ),    .DO85  (RAM15_data_out[213] ),    .DO86  (RAM15_data_out[214] ),    .DO87  (RAM15_data_out[215] ),
    .DO88  (RAM15_data_out[216] ),    .DO89  (RAM15_data_out[217] ),    .DO90  (RAM15_data_out[218] ),    .DO91  (RAM15_data_out[219] ),
    .DO92  (RAM15_data_out[220] ),    .DO93  (RAM15_data_out[221] ),    .DO94  (RAM15_data_out[222] ),    .DO95  (RAM15_data_out[223] ),
    .DO96  (RAM15_data_out[224] ),    .DO97  (RAM15_data_out[225] ),    .DO98  (RAM15_data_out[226] ),    .DO99  (RAM15_data_out[227] ),
    .DO100 (RAM15_data_out[228] ),    .DO101 (RAM15_data_out[229] ),    .DO102 (RAM15_data_out[230] ),    .DO103 (RAM15_data_out[231] ),
    .DO104 (RAM15_data_out[232] ),    .DO105 (RAM15_data_out[233] ),    .DO106 (RAM15_data_out[234] ),    .DO107 (RAM15_data_out[235] ),
    .DO108 (RAM15_data_out[236] ),    .DO109 (RAM15_data_out[237] ),    .DO110 (RAM15_data_out[238] ),    .DO111 (RAM15_data_out[239] ),
    .DO112 (RAM15_data_out[240] ),    .DO113 (RAM15_data_out[241] ),    .DO114 (RAM15_data_out[242] ),    .DO115 (RAM15_data_out[243] ),
    .DO116 (RAM15_data_out[244] ),    .DO117 (RAM15_data_out[245] ),    .DO118 (RAM15_data_out[246] ),    .DO119 (RAM15_data_out[247] ),
    .DO120 (RAM15_data_out[248] ),    .DO121 (RAM15_data_out[249] ),    .DO122 (RAM15_data_out[250] ),    .DO123 (RAM15_data_out[251] ),
    .DO124 (RAM15_data_out[252] ),    .DO125 (RAM15_data_out[253] ),    .DO126 (RAM15_data_out[254] ),    .DO127 (RAM15_data_out[255] ),

    .DI0   (RAM15_data_in[128] ),    .DI1   (RAM15_data_in[129] ),    .DI2   (RAM15_data_in[130] ),    .DI3   (RAM15_data_in[131] ),
    .DI4   (RAM15_data_in[132] ),    .DI5   (RAM15_data_in[133] ),    .DI6   (RAM15_data_in[134] ),    .DI7   (RAM15_data_in[135] ),
    .DI8   (RAM15_data_in[136] ),    .DI9   (RAM15_data_in[137] ),    .DI10  (RAM15_data_in[138] ),    .DI11  (RAM15_data_in[139] ),
    .DI12  (RAM15_data_in[140] ),    .DI13  (RAM15_data_in[141] ),    .DI14  (RAM15_data_in[142] ),    .DI15  (RAM15_data_in[143] ),
    .DI16  (RAM15_data_in[144] ),    .DI17  (RAM15_data_in[145] ),    .DI18  (RAM15_data_in[146] ),    .DI19  (RAM15_data_in[147] ),
    .DI20  (RAM15_data_in[148] ),    .DI21  (RAM15_data_in[149] ),    .DI22  (RAM15_data_in[150] ),    .DI23  (RAM15_data_in[151] ),
    .DI24  (RAM15_data_in[152] ),    .DI25  (RAM15_data_in[153] ),    .DI26  (RAM15_data_in[154] ),    .DI27  (RAM15_data_in[155] ),
    .DI28  (RAM15_data_in[156] ),    .DI29  (RAM15_data_in[157] ),    .DI30  (RAM15_data_in[158] ),    .DI31  (RAM15_data_in[159] ),
    .DI32  (RAM15_data_in[160] ),    .DI33  (RAM15_data_in[161] ),    .DI34  (RAM15_data_in[162] ),    .DI35  (RAM15_data_in[163] ),
    .DI36  (RAM15_data_in[164] ),    .DI37  (RAM15_data_in[165] ),    .DI38  (RAM15_data_in[166] ),    .DI39  (RAM15_data_in[167] ),
    .DI40  (RAM15_data_in[168] ),    .DI41  (RAM15_data_in[169] ),    .DI42  (RAM15_data_in[170] ),    .DI43  (RAM15_data_in[171] ),
    .DI44  (RAM15_data_in[172] ),    .DI45  (RAM15_data_in[173] ),    .DI46  (RAM15_data_in[174] ),    .DI47  (RAM15_data_in[175] ),
    .DI48  (RAM15_data_in[176] ),    .DI49  (RAM15_data_in[177] ),    .DI50  (RAM15_data_in[178] ),    .DI51  (RAM15_data_in[179] ),
    .DI52  (RAM15_data_in[180] ),    .DI53  (RAM15_data_in[181] ),    .DI54  (RAM15_data_in[182] ),    .DI55  (RAM15_data_in[183] ),
    .DI56  (RAM15_data_in[184] ),    .DI57  (RAM15_data_in[185] ),    .DI58  (RAM15_data_in[186] ),    .DI59  (RAM15_data_in[187] ),
    .DI60  (RAM15_data_in[188] ),    .DI61  (RAM15_data_in[189] ),    .DI62  (RAM15_data_in[190] ),    .DI63  (RAM15_data_in[191] ),
    .DI64  (RAM15_data_in[192] ),    .DI65  (RAM15_data_in[193] ),    .DI66  (RAM15_data_in[194] ),    .DI67  (RAM15_data_in[195] ),
    .DI68  (RAM15_data_in[196] ),    .DI69  (RAM15_data_in[197] ),    .DI70  (RAM15_data_in[198] ),    .DI71  (RAM15_data_in[199] ),
    .DI72  (RAM15_data_in[200] ),    .DI73  (RAM15_data_in[201] ),    .DI74  (RAM15_data_in[202] ),    .DI75  (RAM15_data_in[203] ),
    .DI76  (RAM15_data_in[204] ),    .DI77  (RAM15_data_in[205] ),    .DI78  (RAM15_data_in[206] ),    .DI79  (RAM15_data_in[207] ),
    .DI80  (RAM15_data_in[208] ),    .DI81  (RAM15_data_in[209] ),    .DI82  (RAM15_data_in[210] ),    .DI83  (RAM15_data_in[211] ),
    .DI84  (RAM15_data_in[212] ),    .DI85  (RAM15_data_in[213] ),    .DI86  (RAM15_data_in[214] ),    .DI87  (RAM15_data_in[215] ),
    .DI88  (RAM15_data_in[216] ),    .DI89  (RAM15_data_in[217] ),    .DI90  (RAM15_data_in[218] ),    .DI91  (RAM15_data_in[219] ),
    .DI92  (RAM15_data_in[220] ),    .DI93  (RAM15_data_in[221] ),    .DI94  (RAM15_data_in[222] ),    .DI95  (RAM15_data_in[223] ),
    .DI96  (RAM15_data_in[224] ),    .DI97  (RAM15_data_in[225] ),    .DI98  (RAM15_data_in[226] ),    .DI99  (RAM15_data_in[227] ),
    .DI100 (RAM15_data_in[228] ),    .DI101 (RAM15_data_in[229] ),    .DI102 (RAM15_data_in[230] ),    .DI103 (RAM15_data_in[231] ),
    .DI104 (RAM15_data_in[232] ),    .DI105 (RAM15_data_in[233] ),    .DI106 (RAM15_data_in[234] ),    .DI107 (RAM15_data_in[235] ),
    .DI108 (RAM15_data_in[236] ),    .DI109 (RAM15_data_in[237] ),    .DI110 (RAM15_data_in[238] ),    .DI111 (RAM15_data_in[239] ),
    .DI112 (RAM15_data_in[240] ),    .DI113 (RAM15_data_in[241] ),    .DI114 (RAM15_data_in[242] ),    .DI115 (RAM15_data_in[243] ),
    .DI116 (RAM15_data_in[244] ),    .DI117 (RAM15_data_in[245] ),    .DI118 (RAM15_data_in[246] ),    .DI119 (RAM15_data_in[247] ),
    .DI120 (RAM15_data_in[248] ),    .DI121 (RAM15_data_in[249] ),    .DI122 (RAM15_data_in[250] ),    .DI123 (RAM15_data_in[251] ),
    .DI124 (RAM15_data_in[252] ),    .DI125 (RAM15_data_in[253] ),    .DI126 (RAM15_data_in[254] ),    .DI127 (RAM15_data_in[255] ),

    .A0   (RAM_addr[0]   ),.A1   (RAM_addr[1]   ),.A2   (RAM_addr[2]   ),.A3   (RAM_addr[3]   ),.A4   (RAM_addr[4]   ),.A5   (RAM_addr[5]   ),.A6   (RAM_addr[6]   ),
    .DVSE (1'b0  ),.DVS0 (1'b0  ),.DVS1 (1'b0  ),.DVS2 (1'b0  ),.DVS3 (1'b0  ),
    .WEB0 (~w_WEB15_8[0] ),.WEB1 (~w_WEB15_8[1] ),.WEB2 (~w_WEB15_8[2] ),.WEB3 (~w_WEB15_8[3] ),
    .WEB4 (~w_WEB15_8[4] ),.WEB5 (~w_WEB15_8[5] ),.WEB6 (~w_WEB15_8[6] ),.WEB7 (~w_WEB15_8[7] ),

    .CK    (clka   ),
    .CSB   (1'b0   )
);

endmodule